`timescale 1ns / 1ps
`include "Definition.h"
module vga_display_back(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input [2:0] choise,
    output [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;
reg [3:0] red, green, blue;

assign pixel_data = {red, green, blue};

reg [0:639] data [479:0];
//(*ram_style = "block"*) reg [0:639] data [199:0];
always @(posedge vga_clk) begin
if(choise == 0) begin
data[0]<=640'd0;
data[1]<=640'd0;
data[2]<=640'd0;
data[3]<=640'd0;
data[4]<=640'd0;
data[5]<=640'd0;
data[6]<=640'd0;
data[7]<=640'd0;
data[8]<=640'd0;
data[9]<=640'd0;
data[10]<=640'd0;
data[11]<=640'd0;
data[12]<=640'd0;
data[13]<=640'd0;
data[14]<=640'd0;
data[15]<=640'd0;
data[16]<=640'd0;
data[17]<=640'd0;
data[18]<=640'd0;
data[19]<=640'd0;
data[20]<=640'd0;
data[21]<=640'd0;
data[22]<=640'd0;
data[23]<=640'd0;
data[24]<=640'd0;
data[25]<=640'd0;
data[26]<=640'd0;
data[27]<=640'd0;
data[28]<=640'd0;
data[29]<=640'd0;
data[30]<=640'd0;
data[31]<=640'd85070591732710495944414412407740301312;
data[32]<=640'd730750818665451459101842416358132502628711530496;
data[33]<=640'd27021597764222976;
data[34]<=640'd9007199254740992;
data[35]<=640'd9007199254740992;
data[36]<=640'd9007199254740992;
data[37]<=640'd9007199254740992;
data[38]<=640'd9007199254740992;
data[39]<=640'd9007199254740992;
data[40]<=640'd13510798882111488;
data[41]<=640'd9007199254740992;
data[42]<=640'd9007199254740992;
data[43]<=640'd9007199254740992;
data[44]<=640'd9007199254740992;
data[45]<=640'd13510798882111488;
data[46]<=640'd9007199254740992;
data[47]<=640'd9007199254740992;
data[48]<=640'd9007199254740992;
data[49]<=640'd13510798882111488;
data[50]<=640'd31525197391593472;
data[51]<=640'd309787241346054520360140800;
data[52]<=640'd599375721660670508425266668362373856774380817170532873411752110287376594018075499955962254745047801101257078721539110295345450208080468874490806272;
data[53]<=640'd5027929472167778066878457916438579271401010308215785621888644634346722099039006813346457612736872842782101791232293722601083851606530876499670384477470720;
data[54]<=640'd26396628205467732864788082285642163171681467387598851022504789516166031859271295734080499794632056350026575515206137239670386077067062433013666803051659264;
data[55]<=640'd107052979177370224261959331447169757995624348293019147030047829383530188356005728063506518606159218349527795023329677542352008354006734679382389176714395648;
data[56]<=640'd214315455403593848371243628535063509913572769065503325629120859826805569962864356697324533626196254014778770029289013968377661500181271326886728884677509120;
data[57]<=640'd428840407856041074259963789741753073154462173194139026648524031365156604373179187965892171529647976321944478726877311152888398901532830347995215140384407552;
data[58]<=640'd857890312710984452973429432205287855794666022103459363145609269421919230326598971951740951076827667545097005016360117896252295914307608837212705991216332800;
data[59]<=640'd1715990122520767163402835295025441171969567992656791332698788381890886667082526282063613182540215233834685701369746996036155842454675129901135972923267350528;
data[60]<=640'd3381910457608045116620999402357853392069290396874125430328045293723256668427299865470942285888501138062814744645993448611444427055806175678689141383990607872;
data[61]<=640'd6760678458734064500004395559042319423859994262652645444346415197021551412634851879054371547607344496682524987027586199293328324311640523138232093438226989056;
data[62]<=640'd13518213642638457425626434681613824247268059382700472661371176154298941598148001792901619029354125148973649014067957618735459638875554094018914426032008200192;
data[63]<=640'd13303689508433767673001792403097267332445570694662408114543717372905665493958789517438273337383157632243321737455198609118372135649314003991232408626193760256;
data[64]<=640'd26604027063486494151856852108440019966858802187707887285518607084327113815165657061281383825521489522527025728247401310676293068991128914079610415427673391104;
data[65]<=640'd54066572828686917512538848091696728615772215835780101081038941672982135750213955630549554187526714626306345586352280791600468548118337364405108883342695071744;
data[66]<=640'd108126854402215468636948495822802328610646555176645496568601164575687211790167285726112387578570729443792281568925608496419361685686955605409517285680324018176;
data[67]<=640'd106410661329377119006977893772893853047864231581297737945232268808300772200366709756376036593409518210486072502430351275254099497567078879082869518791243464704;
data[68]<=640'd216247436575855479282092410736678649095590945920787579121648876487916844005673158738319991589732162304852207301197122119583818767818967446770323958965500641280;
data[69]<=640'd212814617933244944225846956985053715385389454010758270613221946629202400863949106570233714202028220831395569769179299962980594675440578057599903261196493520896;
data[70]<=640'd425630075491580350373514556489764094002022545108418790299028410609512909024529356069086987000409094756423964141442302784669197120254938147435314767835038744576;
data[71]<=640'd864977176477493792998426720553126075865707973051461377546367259004900087853513061839282910684749462706454618560081417516813094727567860441403240096422265094144;
data[72]<=640'd851247682632341467128970141392075156053575187939118035919251798845312188512943540402250903746277609282808142921882505770245391633396799966707883547220447854592;
data[73]<=640'd1729955184390208237472303383221228712183658530661859015675224928698743183157140205290275958981656649640543026924220237830657450719240773284034815281766284132352;
data[74]<=640'd1702495365258689079671238639778692186686648698691038037051379820481306262388471864585215024917390711291478313796939795069715334066961525319969474466567994474496;
data[75]<=640'd3459883972158554305902524366150836688105814640052773469618604938651459850491363095953710892695995849384108774563596257108611723471560113782663469689111389929472;
data[76]<=640'd3404966402678380287026472699061892275557714108338375202607199483365135647893772515601448216130947937129818071330403331790953794098718246683046836199909150949376;
data[77]<=640'd6919769620281112346282473663417035300574804215453964264447298784452164613972549122915290026490312135640287871664655176173607558561847291296195597047089902649344;
data[78]<=640'd6809932805344772864421133650764320560533861927265129952552077886232105511571101450500741662581779928543593774435373931650172041152181291712486836710752275922944;
data[79]<=640'd13839485504582804636771634314557442765540704517288645763211024595086836483792384167084161877332950073509926851413873715336011710023323021165928452172413373775872;
data[80]<=640'd13619811979458625123224703741313646734349949348047649061338701020815318781929897902843165232488609907086914327981229207162956470717094728387741441325879816880128;
data[81]<=640'd27678971009140035495573996324079679547060880019621936630943123616759766761141886885221954464300421961469106309459060756254840548257620172840974207485516475006976;
data[82]<=640'd27239623539897679053327564100571767080268538237049088531596804344288460452819900738111875815959250704898749886308357836242488687851363195978447168975123953745920;
data[83]<=640'd55357834755792656445893429784966008765323002970073268929816810071248050828911928509004133547621889284623934433607299484814503444967508689819300071169627483275264;
data[84]<=640'd54479247079796955661475752410167943692920068694349925510592349617495011916437736470975248442430863494517913342821690832962759812414814875610540376595600097935360;
data[85]<=640'd110715669511586911227044760910989549664951290921252942767736421845620006903796688988886746286888562537833446547416159306317038729986015682962372443556378803437568;
data[86]<=640'd108958279634617483897186059353955721834531173292492643743446586046970229497852579626815538309591923960744126037655557682374053725383735175296355788649654040657920;
data[87]<=640'd108958276282663903076283488369549075760180252722079693234698334086877633526618490491310064159152584231270217074212862956664341061242741187353202903905637178015744;
data[88]<=640'd221431335671170693240215314621644771431426395490521791277898172646833623334842425363648422135228700058062154206682413788871748700324389950795583538713360416636928;
data[89]<=640'd217916552565331002823165766959398391001306435154144838499707258298812106106143536212746440113533544594240287378617390005937186876393157600823930063484681833152512;
data[90]<=640'd442862242292490821964359011659308181960156777221913368692767379022222992390025038628709715690211444402007032171733189041754440386983041800259773752932296824979456;
data[91]<=640'd442862228884679695448036652215884974418818052233948439596294440625308896041677152899905542243931370874668803798369585865243004234553139213729170333811226439581696;
data[92]<=640'd435833105130508562534745063552623256078125856084596639737079105219936424717994818075581101639306710098286409836474796876868486384501888739015930737911622812041216;
data[93]<=640'd435833078314886309308436457572871538053355971474607200970256890968555190777274628892512546854519477174740741143016318386965325376872929856817777546809377032241152;
data[94]<=640'd421773972706900460565300364381239083639546980409929178366340363577876513135139219757465394741596352353179657050576974825036112800830974047350341605563815455358976;
data[95]<=640'd421773490025814980266866852072168080722746520326731594415381246511774577959324591550086354122775601042723754080244766925928918731942453508047105353713736589770752;
data[96]<=640'd168709267295369864355395194106365450110326787925898158555921256322683905591083810756201579645300549095178113289751200261547810419468161304768314266015640158470144;
data[97]<=640'd9007199271518208;
data[98]<=640'd9007199271518208;
data[99]<=640'd9007199305072640;
data[100]<=640'd13510798898888704;
data[101]<=640'd9007199271518208;
data[102]<=640'd9007199271518208;
data[103]<=640'd9007199271518208;
data[104]<=640'd9007199305072640;
data[105]<=640'd13510798898888704;
data[106]<=640'd9007199271518208;
data[107]<=640'd9007199271518208;
data[108]<=640'd9007199271518208;
data[109]<=640'd9007199271518208;
data[110]<=640'd13510798898888704;
data[111]<=640'd9007199271518208;
data[112]<=640'd9007199271518208;
data[113]<=640'd9007199271518208;
data[114]<=640'd9007199305072640;
data[115]<=640'd13510798898888704;
data[116]<=640'd9007199271518208;
data[117]<=640'd9007199271518208;
data[118]<=640'd9007199271518208;
data[119]<=640'd9007199305072640;
data[120]<=640'd9007199271518208;
data[121]<=640'd9007199271518208;
data[122]<=640'd9007199271518208;
data[123]<=640'd9007199271518208;
data[124]<=640'd9007199271518208;
data[125]<=640'd13510798898888704;
data[126]<=640'd9007199271518208;
data[127]<=640'd9007199271518208;
data[128]<=640'd9007199271518208;
data[129]<=640'd533996758980227548388856843498274930307712532674261077271556721709290300914980308412090940391424;
data[130]<=640'd1868988656430796558311506037023396764362175874785403194374430124751192900551531866420075563057152;
data[131]<=640'd70608395103938906748405908848113786735498346477469127413701232021435384158860502965062554256599959879843061883878768640;
data[132]<=640'd320259506364294327037405639924244233692028483547307954462621785835688912818792645285933467907937828686853293558248505344;
data[133]<=640'd1636695303852802729735721062057007209171471377742890289643062904937418624395482718595003351178232432600793374821907689755208590573672079544628279246848;
data[134]<=640'd1636695303852802729735721062058147030406720677237543099851066895318485373478903061535747386712734283593220464541437540325981490295668695865160609300480;
data[135]<=640'd1636695303852802729735721062065404564732046969152611200271195788852249740197418431205925877357108034363812204308885191990930668944454828233263325118464;
data[136]<=640'd1432108391621439505026886996886717169273864967559035645802998680124266543704676409646449470163531041179254364961423359278795446832131342830488728371200;
data[137]<=640'd1432108391621439505026886996904792918420473327686627080007019763244601044180741872875958218823407205924272963993675377937932973822672338671949406273536;
data[138]<=640'd1432108391621439505026886996940944416713690047941809952687036001327029501520034157640508399872311787975085208710858581108289465131830540530627962208256;
data[139]<=640'd1432108391621439505026886997013247413300123488452175689503120333808321972122134470033220033847614419284429732306322481390539143083906703564612258758656;
data[140]<=640'd1432108391621439505026886996992589414275428219734928335071630492107686374016258216053810355123933847131021312988412579121760328376010588614750415880192;
data[141]<=640'd1438501708263826107773067200574440595710413292009303674706163034184736318488786445288231027768489408390551455490014148558540112382132240449363983204352;
data[142]<=640'd1438501708263826107773067200905112324530611555697776182677881604841364878485544834097304301566202876957463908960600784381609845588812803537031045054464;
data[143]<=640'd1438501708263826107773067200823611324858682238667124598499346632091097017956705033809947116106813684914271999279295423637327699940550686502619315175424;
data[144]<=640'd1438501708263826107773067201323246436537238515940420174492130866768986460830840368098883116633055999418160435102198599573719690396074069642355528433664;
data[145]<=640'd1438501708263826107773067201322962740813441439457109761583034352706409608873262240980858385615278939318779762280298122657646878248325483011038393663488;
data[146]<=640'd1438501708263826107773067202312297309787738345839875981067882261633881989358028662215501224530230193504744836927753656721722281519100185974841261686784;
data[147]<=640'd1438501708263826107773067202309715054984254465367451376283259637096398556801914921456373845917349145277493652774308822503213564773201498818347301601280;
data[148]<=640'd1438501708263826107773067202309732707084522954598918008415798489359989066652640762027133268951647952458608815625633188054076831696503447797863775469568;
data[149]<=640'd1438501708263826107773067202309768050686478991570927280503415492089160941891970074339170593665702809496375178098731523621550020287451338742925027704832;
data[150]<=640'd1438501708263826107773067202309848736144526745273229086695513425302448813404944478720520681834899876522488497296199062363961010652565782525297207279616;
data[151]<=640'd1438501708263826107773067202640528024242994277653415346277159249999999682165383556445927478766297169811298765766314058727337797412710454030339030384640;
data[152]<=640'd1438501708263826107773067202640830631649982238765905294379567146994319168831492556122191299623390740742054492039624243994098153348564249012274095718400;
data[153]<=640'd1438501708263826107773067201485798409517193899444102656796441397993625284904625016300391696264886638598651896272353560065744139537532355271058561957888;
data[154]<=640'd1438501708263826107773067200987262772728632956610153777650158933238602953326497741304358027431757108917308735210185175675280377471521256380509953458176;
data[155]<=640'd1438501708263826107773067200655766444626819975358548998235631410281896786752360085236610547710231679244496890731981817430355582768606249983016532180992;
data[156]<=640'd1438501708263826107773067200398832502951340050453914034473356873165588656285070363517185675721137460733609444265944369714287184776974375807963321335808;
data[157]<=640'd1438501708263826107773067200326529466962317972766699079742782072606113783650612821291620594761390321761360491071143119989379591963352437851729424285696;
data[158]<=640'd1438501708263826107773067200326529466962317972766699079743694664723511633417261084960027996177541379601722830511428110910690354785646412696099586310144;
data[159]<=640'd1432108391621439505026886996868641420127256607431444208398647411592158318702671441836255319300660893909043208523209351375611244346730489970972357033984;
data[160]<=640'd1432108391621439505026886996868641420127256607431444208402297780061749717769264496509884924965265125270492566284349315060854295635906389348453005131776;
data[161]<=640'd1432108391621439505026886996868641420127256607431444208426285915719064625921161712936593762189807217074302631571840504992451489821919442400468675854336;
data[162]<=640'd1432108391621439505026886996868641420127256607431444208657823572933147652430778323663957321487561320571947609564146773027867885878219345772098355200000;
data[163]<=640'd1432108391621439505026886996868641420127256607431444208645308023894548569916744993354370102066061098761264097240238326107034567172473405049307561721856;
data[164]<=640'd1636695303852802729735721062055718605960824492694731914513886315868436735039865809623431264300745114147225121181134921005965207090773500786651179253760;
data[165]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[166]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[167]<=640'd0;
data[168]<=640'd0;
data[169]<=640'd0;
data[170]<=640'd0;
data[171]<=640'd0;
data[172]<=640'd0;
data[173]<=640'd0;
data[174]<=640'd0;
data[175]<=640'd0;
data[176]<=640'd0;
data[177]<=640'd0;
data[178]<=640'd0;
data[179]<=640'd0;
data[180]<=640'd0;
data[181]<=640'd0;
data[182]<=640'd0;
data[183]<=640'd0;
data[184]<=640'd0;
data[185]<=640'd0;
data[186]<=640'd0;
data[187]<=640'd0;
data[188]<=640'd0;
data[189]<=640'd0;
data[190]<=640'd0;
data[191]<=640'd0;
data[192]<=640'd0;
data[193]<=640'd0;
data[194]<=640'd0;
data[195]<=640'd0;
data[196]<=640'd0;
data[197]<=640'd0;
data[198]<=640'd0;
data[199]<=640'd0;
data[200]<=640'd0;
data[201]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[202]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[203]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
data[204]<=640'd716054195810719752513443498452396459210236663843313538401519604681591400367843758171127472313812864627914813743442211318145061348828617500555078533120;
data[205]<=640'd716054195810719752513443498454817318470943140646115962625272428313775499548621155214406215460569721773555602363407503836845190565799776724279529308160;
data[206]<=640'd716054195810719752513443498516942619248823106185030406280912270583849488969373445934094087849421263174083520826805540203121430985236360613379530817536;
data[207]<=640'd716054195810719752513443498599582180532793891087527193434379346215841788567102110100978117211933049057178062906913029171650412120303285071331498917888;
data[208]<=640'd716054195810719752513443498594424617992336026611211666968870954002199316658579354529295692867369532881627382597869581719349971971229802136622671593472;
data[209]<=640'd716054195810719752513443498470474108272331322421689801733046036933826550285750168652928145848503239957568531354763767237227511749508443218334678253568;
data[210]<=640'd716054195810719752513443498465308672718510340873496671745117643480671118166195844841114120965026022274926009181593149300629143946687042173319644184576;
data[211]<=640'd716054195810719752513443498506624657223461246003890533286174287434856891565124599078778989884953122375513294241757993247051690560743735994951435026432;
data[212]<=640'd716054195810719752513443498506624652298210471454580631885054205267145339708975597071443380104758889826892124014399521046811419350104215025143861215232;
data[213]<=640'd716054195810719752513443498496295652785862855443945883084174268069311714182345803205975936425142028849943491336863722245241643132224477161940351713280;
data[214]<=640'd716054195810719752513443498578928594532792639193439159305090028273801748502798542518557450139198694610470892581121084791661332217742187629441106051072;
data[215]<=640'd716054195810719752513443498578935529295615565084795285312521661142683621566827201523159863495089171062366134461495250180271803632698486581077173338112;
data[216]<=640'd716054195810719752513443498558306559719295686255939994691463852412789730990382003880051374333913264620660854005355689082322410824234160602443344248832;
data[217]<=640'd716054195810719752513443498723684029695915337013595158856156430908443933135962537296006781336619137107590586039828334070534992578101058502990789345280;
data[218]<=640'd716054195810719752513443498726074667662435116152319054365729584236292666552544995954241525497930953128181220600548079562723803871197520873352868134912;
data[219]<=640'd716054195810719752513443498764687372869500969648166995387713925429748206448310492740292313345780339563283646892842795758416380402056113891813774852096;
data[220]<=640'd716054195810719752513443498762266503828035350362723319525822871017568885791056302026571382589134451089783145982566227641658649420802696355669019197440;
data[221]<=640'd716054195810719752513443499012744741992836455529709340851102690530689620425974536127085317615947573415639164249983869881973447411020431322848130236416;
data[222]<=640'd716054195810719752513443498930112824678828498850708675602916998574373097638935264627451193163361309192489206596011604979186284746446998068957171154944;
data[223]<=640'd716054195810719752513443498930112805131814622444746571190038572981539243817399858943490253968280715111299464596629928971483814150922352367596472369152;
data[224]<=640'd716054195810719752513443499591168773883566058145757224900889316156738702612168354968539617553353773703844976370883228066977480014210530902843334852608;
data[225]<=640'd716054195810719752513443499591168931491741113896338500626710837487951928012927739405129935394457478811456723544995424280807755658899542164501228945408;
data[226]<=640'd716054195810719752513443499425904939601969561137220759507440701221919135022913033671278759931037052797222372081332600693355028792468667943584333299712;
data[227]<=640'd716054195810719752513443499425904900123006321892684327391627979833966398203541687810086025966492434445610482967791808411731173206438044431614669225984;
data[228]<=640'd716054195810719752513443500748016837703804356719440658621889048670187383705742252154792706093711491586733855110068319510099229844196759380564610383872;
data[229]<=640'd716054195810719752513443500748017152919778787986916839628238819076166832342626120149144509311646161009324757501601892866314905534279262675934774296576;
data[230]<=640'd716054195810719752513443500417489168524654615226286366532113576586219958341702119533547297296133204822806923134614207553653809644564894950407257718784;
data[231]<=640'd716054195810719752513443499756432805560279541931114698735649863252824271402368568143057938395255371826363848621175488615897430102674974581120177274880;
data[232]<=640'd818347651926401364867860531027859302980412393131277380521395508717963006741230473315177183548362701793830182762363954799343770380606623659043181297664;
data[233]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[234]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[235]<=640'd0;
data[236]<=640'd0;
data[237]<=640'd0;
data[238]<=640'd0;
data[239]<=640'd0;
data[240]<=640'd0;
data[241]<=640'd0;
data[242]<=640'd0;
data[243]<=640'd0;
data[244]<=640'd0;
data[245]<=640'd0;
data[246]<=640'd0;
data[247]<=640'd0;
data[248]<=640'd0;
data[249]<=640'd0;
data[250]<=640'd0;
data[251]<=640'd0;
data[252]<=640'd0;
data[253]<=640'd0;
data[254]<=640'd0;
data[255]<=640'd0;
data[256]<=640'd0;
data[257]<=640'd0;
data[258]<=640'd0;
data[259]<=640'd0;
data[260]<=640'd0;
data[261]<=640'd0;
data[262]<=640'd0;
data[263]<=640'd0;
data[264]<=640'd0;
data[265]<=640'd0;
data[266]<=640'd0;
data[267]<=640'd0;
data[268]<=640'd0;
data[269]<=640'd0;
data[270]<=640'd0;
data[271]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[272]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[273]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[274]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[275]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[276]<=640'd716054195810719752513443498436902329509616069993710626904859931137792284335040089646996829001874510964265422620294556570204156201562945562670748663808;
data[277]<=640'd716054195810719752513443498475636077680919698838549414484905109252737871227478442339456719349984225294518040539739236869406223673101493142261961064448;
data[278]<=640'd716054195810719752513443498764203131989230876044265778420883288506903374851972497345429589616096064986448387994971887726721704494713925516264338358272;
data[279]<=640'd716054195810719752513443501075962335346535790933735072534116409542307789640129758881856114652118974840552957684284325086262295903437522520986112491520;
data[280]<=640'd716054195810719752513443508936330964243310997934299320101161945139223999366914197463078394669438236193084646203335782881574369898171715801520548085760;
data[281]<=640'd716054195810719752513443519265330476590982933239308044822392414689331103834041171381277090042968167159521430263441464572718312641489842287878613237760;
data[282]<=640'd716054195810719752513443518284075522917920092488719067374528189671023665650908402235286529253574501650522280565529526920176121880409916046746893418496;
data[283]<=640'd716054195810719752513443498452396459210462123931259826391396994818883176722471823695822671021400764561181905809853213728717576452673555296046144290816;
data[284]<=640'd716054195810719752513443498449814209332375215341603907219393982944553470929642600182992011664860116939165064615223568375437438621237652124073396797440;
data[285]<=640'd716054195810719752513443498449814209332675828792198959741552492891738828164790680447610376885677107245592361074099645100643052151091383788153310543872;
data[286]<=640'd716054195810719752513443498470472208357296532456069495355220800717315295409424067509323404103846287738224339862431283562756427942171383677257546465280;
data[287]<=640'd716054195810719752513443498470472245296789193897524885153498362561344464051193620122991184124157306732063564090470508834172320742291097521131574263808;
data[288]<=640'd716054195810719752513443498465307865602658693133458516961066248897713390654644228328779303032332226412839833220615876792369138435907871673042136465408;
data[289]<=640'd716054195810719752513443498465307988733919250055530179090002669739408021728330603250509907113241755854240066293028306935115618068248898069690446774272;
data[290]<=640'd716054195810719752513443498506624260127372139531325437036200070719626186885047975754102994146508111398543647493240509431258382984310276384408731648000;
data[291]<=640'd716054195810719752513443498496295814704383881295676062170550081767161153415043803623859074324190431956418429410889029815587060889478067374352666460160;
data[292]<=640'd716054195810719752513443498496295662022812323782761870587916157253896573255094066940805254400867231041917333922361192552993492372979840399978975461376;
data[293]<=640'd716054195810719752513443498496296951822858908309987685876216829396839914528060514285023767266729571651450982271288846974036962317272084211347933364224;
data[294]<=640'd716054195810719752513443498578931741769841824547066520502883281936589987764275614399516277332028591823409897256980011086917888149978517610143791710208;
data[295]<=640'd716054195810719752513443498558278771426188544946502498052319976344874161232557918827616281603359197962840568093369515775553924105436891689389884702720;
data[296]<=640'd716054195810719752513443498558278475911141483705513398365213768819594491263525670780384220844274925653013265520827590983322030889469131576425356197888;
data[297]<=640'd716054195810719752513443498558272486806201980287395889563734169743938988323341750211228189541787287895625183229269806637466046417796349828133076074496;
data[298]<=640'd716054195810719752513443498723536479927252173067244483859558766269051291626509507707747657120232923303169422018570654865081928527056940318848807075840;
data[299]<=640'd716054195810719752513443498723536481158874883499457587595962191555952092861975347895139843247036184052869221329693412692250148544623692447520611368960;
data[300]<=640'd716054195810719752513443498682221130472412500164015030748316599426718847179850664840786266601969270520428233878680726559662575733659658746413042368512;
data[301]<=640'd716054195810719752513443498682219217626935783688236265452195436977737437282247049624759838328005796649578242945000593351105964490429237779900150054912;
data[302]<=640'd818347651926401364867860531027860544143832906622819285070802166648325145936293367879823861257253301713640055421807465536124401416969883210374893797376;
data[303]<=640'd818347651926401364867860531027859302980412246347505941203204878388585547550201790102400479621947948184075711318110122128264813958505529454328717246464;
data[304]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[305]<=640'd0;
data[306]<=640'd0;
data[307]<=640'd0;
data[308]<=640'd0;
data[309]<=640'd0;
data[310]<=640'd0;
data[311]<=640'd0;
data[312]<=640'd0;
data[313]<=640'd0;
data[314]<=640'd0;
data[315]<=640'd0;
data[316]<=640'd0;
data[317]<=640'd0;
data[318]<=640'd0;
data[319]<=640'd0;
data[320]<=640'd0;
data[321]<=640'd0;
data[322]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[323]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[324]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[325]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[326]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[327]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[328]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[329]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[330]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[331]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[332]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[333]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[334]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[335]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[336]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[337]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[338]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[339]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[340]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[341]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[342]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[343]<=640'd398353494612575324017191154914352288844846764696638810260114131509605650307885529420329033517687589677374404780947210779386712874022118574019139283960076830011772872351155913515597824;
data[344]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[345]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[346]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[347]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[348]<=640'd398353494612575324017191154914352186551390649015026455843081537971012733523942897776476074197443525535126815153878457074366752531570804226482521018768785698054402230421841660119875584;
data[349]<=640'd265568996408383549344794103276235029718992369583268475043220513910041109088511359234064155610167347940571714494382458401709398254602728763359583467446130040472067320563817398958817280;
data[350]<=640'd265568996408383549344794103276235029718992369583268475043220542153399150664074058595680099393109723421728823564014629987046110417936094572560149729192181541979598650754760850884526080;
data[351]<=640'd265568996903044352291003171397240071758286749653531173245644265870947140976898850940200584448743909205504922481436351689200150496414012795173930077975219068851482267557512510571544576;
data[352]<=640'd265568996903044352291003171397240071758286749653531173245644265558252819896327359178219133617954960188615259508155358968348673864571206520720809202410771322490992271206384922743799808;
data[353]<=640'd398353495107236126963400223035357228590685029085289154045505297848885066685838825189461651410739422896187426297242838665317545949164137665328712269515090178962203775974916756376387584;
data[354]<=640'd265568996903044352291003171397240071758286749653531173245644338184030641034303117242229689877502164522971427564103021196670092171290393849036582324453145440167845741598409794485485568;
data[355]<=640'd265568996903044352291003171397240071758286749653531173245644327855031128611515395969790338572991288106889471371187128308966430146066594692641115002204262128778152049673123406473592832;
data[356]<=640'd265568996903044352291003171397240071758286749653531173245644307197032103916246678722436962548896293469243128737399025663691577820885618557911557965041435887675500562447747624493645824;
data[357]<=640'd265568997892365958183421307639250155836875509794056569650491832117276525850132101038814803999664947352685383330305512689261723771658093458695782166283893464620766319316229012867514368;
data[358]<=640'd265568996903044352291003171397240071758286749653531173245644472461063818920267927613494590438064006976687019289681191333776707214442910372948086204241920481272126874592137966946091008;
data[359]<=640'd265568996903044352291003171397240071758286749653531173245644431205607106415498351048945982500342200140279227042640518206448955333946888070244009063416593263508288873275499490247180288;
data[360]<=640'd265568996903044352291003171397240071758286749653531173245644431770484387098227638060986536861113849285553400473186921434630770436779591819154968957088195460873412620290859285490958336;
data[361]<=640'd265568996903044352291003171397240071758286749653531173245644766756845724655747473510255706594824695543368075391008313367673797349528654530894869267351649187414430494941395726620426240;
data[362]<=640'd265568996903044352291003171397240071758286749653531173245644843659480909080866790552231080676368793600226952876822552707429198519299934820975122398871077385613727999725727203415031808;
data[363]<=640'd398353495107236126963400223035357228590685029085289154045505876272876844122221199281299545126859726022122334059205504615661116760422648465263434564713455934430047793314326588816359424;
data[364]<=640'd265568996903044352291003171397240071758286749653531173245645484702994982139725872965258139836562807659282043279684631898945903919829267023699733195241668281122035439496027543105961984;
data[365]<=640'd265568996903044352291003171397240071758286749653531173245645340097000579162458233375088372050565688726667460553454196218566568069607323140557732441880137923280415860907149770532847616;
data[366]<=640'd265568996903044352291003171397240071758286749653531173245645174833028082302793242040816850208002287043364119848697241519436780164328392567484269535213354364233174627674152840600748032;
data[367]<=640'd265568997892365958183421307639250155836875509794056569650493856601337324502862867062672605271651108427048876329190094906304104597697945171522775673170267909795562382300825067007770624;
data[368]<=640'd398353495107236126963400223035357228590685029085289154045507531495314049022707758805221808527669066460065147963112017655568023638169995171863509723114198942463964854009681611778424832;
data[369]<=640'd265568996903044352291003171397240071758286749653531173245646166982367429213654653607639590747946535849447754254214342759981391193928366993523644887359573947682335248412627898218840064;
data[370]<=640'd265568996903044352291003171397240071758286749653531173245646168838908693948757269410713320960433747478933289273331719673164322356616834544702525663131062790607969032125819749335564288;
data[371]<=640'd265568996903044352291003171397240071758286749653531173245648820651452948170946773728445373595175963805733747734958428812846622296264991660556917029629575456997943970807968902695354368;
data[372]<=640'd265568997892365958183421307639250155836875509794056569650496830070743775665005331346202969610616535024674669991064294781277940123279233337905270013843241342490693245972345363328139264;
data[373]<=640'd265568996903044352291003171397240174051742865335143527662682054913947799261606721964401616714338507026402603841286661204148291631905629204376219183101830592291163931199020767880675328;
data[374]<=640'd265568996903044352291003171397240174051742865335143527662679255747514454022224283900141070411542534696719932584147492194075207522237814138723162892139430987789628858278988575806586880;
data[375]<=640'd265568996903044352291003171397240174051742865335143527662676776787630872528466918948602142292013070382638162388580928377582346718311671832780261709203522302229601390475521153055064064;
data[376]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[377]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[378]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[379]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[380]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[381]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[382]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[383]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[384]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[385]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[386]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[387]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[388]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[389]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[390]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[391]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[392]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[393]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[394]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[395]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[396]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[397]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[398]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[399]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[400]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[401]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[402]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[403]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[404]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[405]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083711154225492614732989228270490262743671417864192;
data[406]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083756826325883777643510875830043263955216103374848;
data[407]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083733993150393632101736882977413894943200384122880;
data[408]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260510356823990064450203354978959320258094768848896;
data[409]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841306678842167437339742438259765413224120320;
data[410]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841295784489368253867537777416344549361451008;
data[411]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083866058175805198939743815208226653779662768963584;
data[412]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934544014703162186716804046514368768030868556417597440;
data[413]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260686614913495185286957388911191037195542417375232;
data[414]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083871185952298368884399164504508543769418921934848;
data[415]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986330444476161582688175652864;
data[416]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[417]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[418]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[419]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[420]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[421]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[422]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[423]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[424]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[425]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[426]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[427]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[428]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[429]<=640'd398353496343888134328922893337869117634725168541193386108065983048744062545919757800094946891136771680368312041868575743622909878699085669704398453847763599671125628542792319314690048;
data[430]<=640'd531137992816767098689588206552468627329593117540961209779768774219776665041523081944630313929275862236827838496002843258316710966147798256686047195211381820739689719850535202106376192;
data[431]<=640'd464745747548292448942947204772883260336491728765709340960903687623617040888630979714838395224460056055998811059991606943419003558340812870361086397939032316978126257926111479799480320;
data[432]<=640'd1731312810311731738423517647137530330245919443708482879398441392650280575745723070192214807428701314927183699982112975375459555240147258469772823085713252175416247405040893952;
data[433]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[434]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[435]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[436]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[437]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[438]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[439]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[440]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[441]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[442]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[443]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[444]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[445]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[446]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[447]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[448]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[449]<=640'd741991204419313602181507563058941570105394047303635519742189168278691675319595601510949203183729134968793014278048418018054095102920253629902638465305679503749820316446097408;
data[450]<=640'd989321605892418136242010084078576565810250724560193525292073344815707069964632683637707560663098643350035920994610962411690368371714661765920491625786887328011429868730318848;
data[451]<=640'd1799565517869652802850553672994603778697120433756232925976991265676467694158133288870091067319688664337182830767822544995324267558345195980337572361199321983483904;
data[452]<=640'd0;
data[453]<=640'd0;
data[454]<=640'd0;
data[455]<=640'd0;
data[456]<=640'd0;
data[457]<=640'd0;
data[458]<=640'd0;
data[459]<=640'd0;
data[460]<=640'd0;
data[461]<=640'd0;
data[462]<=640'd0;
data[463]<=640'd0;
data[464]<=640'd0;
data[465]<=640'd0;
data[466]<=640'd0;
data[467]<=640'd0;
data[468]<=640'd0;
data[469]<=640'd0;
data[470]<=640'd0;
data[471]<=640'd0;
data[472]<=640'd0;
data[473]<=640'd0;
data[474]<=640'd0;
data[475]<=640'd0;
data[476]<=640'd0;
data[477]<=640'd0;
data[478]<=640'd0;
data[479]<=640'd0;
end
else if(choise == 1) begin
data[0]<=640'd0;
data[1]<=640'd0;
data[2]<=640'd0;
data[3]<=640'd0;
data[4]<=640'd0;
data[5]<=640'd0;
data[6]<=640'd0;
data[7]<=640'd0;
data[8]<=640'd0;
data[9]<=640'd0;
data[10]<=640'd0;
data[11]<=640'd0;
data[12]<=640'd0;
data[13]<=640'd0;
data[14]<=640'd0;
data[15]<=640'd0;
data[16]<=640'd0;
data[17]<=640'd0;
data[18]<=640'd0;
data[19]<=640'd0;
data[20]<=640'd0;
data[21]<=640'd0;
data[22]<=640'd0;
data[23]<=640'd0;
data[24]<=640'd0;
data[25]<=640'd0;
data[26]<=640'd0;
data[27]<=640'd0;
data[28]<=640'd0;
data[29]<=640'd0;
data[30]<=640'd0;
data[31]<=640'd85070591732710495944414412407740301312;
data[32]<=640'd730750818665451459101842416358132502628711530496;
data[33]<=640'd27021597764222976;
data[34]<=640'd9007199254740992;
data[35]<=640'd9007199254740992;
data[36]<=640'd9007199254740992;
data[37]<=640'd9007199254740992;
data[38]<=640'd9007199254740992;
data[39]<=640'd9007199254740992;
data[40]<=640'd13510798882111488;
data[41]<=640'd9007199254740992;
data[42]<=640'd9007199254740992;
data[43]<=640'd9007199254740992;
data[44]<=640'd9007199254740992;
data[45]<=640'd13510798882111488;
data[46]<=640'd9007199254740992;
data[47]<=640'd9007199254740992;
data[48]<=640'd9007199254740992;
data[49]<=640'd13510798882111488;
data[50]<=640'd31525197391593472;
data[51]<=640'd309787241346054520360140800;
data[52]<=640'd599375721660670508425266668362373856774380817170532873411752110287376594018075499955962254745047801101257078721539110295345450208080468874490806272;
data[53]<=640'd5027929472167778066878457916438579271401010308215785621888644634346722099039006813346457612736872842782101791232293722601083851606530876499670384477470720;
data[54]<=640'd26396628205467732864788082285642163171681467387598851022504789516166031859271295734080499794632056350026575515206137239670386077067062433013666803051659264;
data[55]<=640'd107052979177370224261959331447169757995624348293019147030047829383530188356005728063506518606159218349527795023329677542352008354006734679382389176714395648;
data[56]<=640'd214315455403593848371243628535063509913572769065503325629120859826805569962864356697324533626196254014778770029289013968377661500181271326886728884677509120;
data[57]<=640'd428840407856041074259963789741753073154462173194139026648524031365156604373179187965892171529647976321944478726877311152888398901532830347995215140384407552;
data[58]<=640'd857890312710984452973429432205287855794666022103459363145609269421919230326598971951740951076827667545097005016360117896252295914307608837212705991216332800;
data[59]<=640'd1715990122520767163402835295025441171969567992656791332698788381890886667082526282063613182540215233834685701369746996036155842454675129901135972923267350528;
data[60]<=640'd3381910457608045116620999402357853392069290396874125430328045293723256668427299865470942285888501138062814744645993448611444427055806175678689141383990607872;
data[61]<=640'd6760678458734064500004395559042319423859994262652645444346415197021551412634851879054371547607344496682524987027586199293328324311640523138232093438226989056;
data[62]<=640'd13518213642638457425626434681613824247268059382700472661371176154298941598148001792901619029354125148973649014067957618735459638875554094018914426032008200192;
data[63]<=640'd13303689508433767673001792403097267332445570694662408114543717372905665493958789517438273337383157632243321737455198609118372135649314003991232408626193760256;
data[64]<=640'd26604027063486494151856852108440019966858802187707887285518607084327113815165657061281383825521489522527025728247401310676293068991128914079610415427673391104;
data[65]<=640'd54066572828686917512538848091696728615772215835780101081038941672982135750213955630549554187526714626306345586352280791600468548118337364405108883342695071744;
data[66]<=640'd108126854402215468636948495822802328610646555176645496568601164575687211790167285726112387578570729443792281568925608496419361685686955605409517285680324018176;
data[67]<=640'd106410661329377119006977893772893853047864231581297737945232268808300772200366709756376036593409518210486072502430351275254099497567078879082869518791243464704;
data[68]<=640'd216247436575855479282092410736678649095590945920787579121648876487916844005673158738319991589732162304852207301197122119583818767818967446770323958965500641280;
data[69]<=640'd212814617933244944225846956985053715385389454010758270613221946629202400863949106570233714202028220831395569769179299962980594675440578057599903261196493520896;
data[70]<=640'd425630075491580350373514556489764094002022545108418790299028410609512909024529356069086987000409094756423964141442302784669197120254938147435314767835038744576;
data[71]<=640'd864977176477493792998426720553126075865707973051461377546367259004900087853513061839282910684749462706454618560081417516813094727567860441403240096422265094144;
data[72]<=640'd851247682632341467128970141392075156053575187939118035919251798845312188512943540402250903746277609282808142921882505770245391633396799966707883547220447854592;
data[73]<=640'd1729955184390208237472303383221228712183658530661859015675224928698743183157140205290275958981656649640543026924220237830657450719240773284034815281766284132352;
data[74]<=640'd1702495365258689079671238639778692186686648698691038037051379820481306262388471864585215024917390711291478313796939795069715334066961525319969474466567994474496;
data[75]<=640'd3459883972158554305902524366150836688105814640052773469618604938651459850491363095953710892695995849384108774563596257108611723471560113782663469689111389929472;
data[76]<=640'd3404966402678380287026472699061892275557714108338375202607199483365135647893772515601448216130947937129818071330403331790953794098718246683046836199909150949376;
data[77]<=640'd6919769620281112346282473663417035300574804215453964264447298784452164613972549122915290026490312135640287871664655176173607558561847291296195597047089902649344;
data[78]<=640'd6809932805344772864421133650764320560533861927265129952552077886232105511571101450500741662581779928543593774435373931650172041152181291712486836710752275922944;
data[79]<=640'd13839485504582804636771634314557442765540704517288645763211024595086836483792384167084161877332950073509926851413873715336011710023323021165928452172413373775872;
data[80]<=640'd13619811979458625123224703741313646734349949348047649061338701020815318781929897902843165232488609907086914327981229207162956470717094728387741441325879816880128;
data[81]<=640'd27678971009140035495573996324079679547060880019621936630943123616759766761141886885221954464300421961469106309459060756254840548257620172840974207485516475006976;
data[82]<=640'd27239623539897679053327564100571767080268538237049088531596804344288460452819900738111875815959250704898749886308357836242488687851363195978447168975123953745920;
data[83]<=640'd55357834755792656445893429784966008765323002970073268929816810071248050828911928509004133547621889284623934433607299484814503444967508689819300071169627483275264;
data[84]<=640'd54479247079796955661475752410167943692920068694349925510592349617495011916437736470975248442430863494517913342821690832962759812414814875610540376595600097935360;
data[85]<=640'd110715669511586911227044760910989549664951290921252942767736421845620006903796688988886746286888562537833446547416159306317038729986015682962372443556378803437568;
data[86]<=640'd108958279634617483897186059353955721834531173292492643743446586046970229497852579626815538309591923960744126037655557682374053725383735175296355788649654040657920;
data[87]<=640'd108958276282663903076283488369549075760180252722079693234698334086877633526618490491310064159152584231270217074212862956664341061242741187353202903905637178015744;
data[88]<=640'd221431335671170693240215314621644771431426395490521791277898172646833623334842425363648422135228700058062154206682413788871748700324389950795583538713360416636928;
data[89]<=640'd217916552565331002823165766959398391001306435154144838499707258298812106106143536212746440113533544594240287378617390005937186876393157600823930063484681833152512;
data[90]<=640'd442862242292490821964359011659308181960156777221913368692767379022222992390025038628709715690211444402007032171733189041754440386983041800259773752932296824979456;
data[91]<=640'd442862228884679695448036652215884974418818052233948439596294440625308896041677152899905542243931370874668803798369585865243004234553139213729170333811226439581696;
data[92]<=640'd435833105130508562534745063552623256078125856084596639737079105219936424717994818075581101639306710098286409836474796876868486384501888739015930737911622812041216;
data[93]<=640'd435833078314886309308436457572871538053355971474607200970256890968555190777274628892512546854519477174740741143016318386965325376872929856817777546809377032241152;
data[94]<=640'd421773972706900460565300364381239083639546980409929178366340363577876513135139219757465394741596352353179657050576974825036112800830974047350341605563815455358976;
data[95]<=640'd421773490025814980266866852072168080722746520326731594415381246511774577959324591550086354122775601042723754080244766925928918731942453508047105353713736589770752;
data[96]<=640'd168709267295369864355395194106365450110326787925898158555921256322683905591083810756201579645300549095178113289751200261547810419468161304768314266015640158470144;
data[97]<=640'd9007199271518208;
data[98]<=640'd9007199271518208;
data[99]<=640'd9007199305072640;
data[100]<=640'd13510798898888704;
data[101]<=640'd9007199271518208;
data[102]<=640'd9007199271518208;
data[103]<=640'd9007199271518208;
data[104]<=640'd9007199305072640;
data[105]<=640'd13510798898888704;
data[106]<=640'd9007199271518208;
data[107]<=640'd9007199271518208;
data[108]<=640'd9007199271518208;
data[109]<=640'd9007199271518208;
data[110]<=640'd13510798898888704;
data[111]<=640'd9007199271518208;
data[112]<=640'd9007199271518208;
data[113]<=640'd9007199271518208;
data[114]<=640'd9007199305072640;
data[115]<=640'd13510798898888704;
data[116]<=640'd9007199271518208;
data[117]<=640'd9007199271518208;
data[118]<=640'd9007199271518208;
data[119]<=640'd9007199305072640;
data[120]<=640'd9007199271518208;
data[121]<=640'd9007199271518208;
data[122]<=640'd9007199271518208;
data[123]<=640'd9007199271518208;
data[124]<=640'd9007199271518208;
data[125]<=640'd13510798898888704;
data[126]<=640'd9007199271518208;
data[127]<=640'd9007199271518208;
data[128]<=640'd9007199271518208;
data[129]<=640'd533996758980227548388856843498274930307712532674261077271556721709290300914980308412090940391424;
data[130]<=640'd1868988656430796558311506037023396764362175874785403194374430124751192900551531866420075563057152;
data[131]<=640'd70608395103938906748405908848113786735498346477469127413701232021435384158860502965062554256599959879843061883878768640;
data[132]<=640'd320259506364294327037405639924244233692028483547307954462621785835688912818792645285933467907937828686853293558248505344;
data[133]<=640'd1636695303852802729735721062057007209171471377742890289643062904937418624395482718595003351178232432600793374821907689755208590573672079544628279246848;
data[134]<=640'd1636695303852802729735721062058147030406720677237543099851066895318485373478903061535747386712734283593220464541437540325981490295668695865160609300480;
data[135]<=640'd1636695303852802729735721062065404564732046969152611200271195788852249740197418431205925877357108034363812204308885191990930668944454828233263325118464;
data[136]<=640'd1432108391621439505026886996886717169273864967559035645802998680124266543704676409646449470163531041179254364961423359278795446832131342830488728371200;
data[137]<=640'd1432108391621439505026886996904792918420473327686627080007019763244601044180741872875958218823407205924272963993675377937932973822672338671949406273536;
data[138]<=640'd1432108391621439505026886996940944416713690047941809952687036001327029501520034157640508399872311787975085208710858581108289465131830540530627962208256;
data[139]<=640'd1432108391621439505026886997013247413300123488452175689503120333808321972122134470033220033847614419284429732306322481390539143083906703564612258758656;
data[140]<=640'd1432108391621439505026886996992589414275428219734928335071630492107686374016258216053810355123933847131021312988412579121760328376010588614750415880192;
data[141]<=640'd1432108391621439505026886997116552548875351926674048803359290596818587304240900274827643548059306807017147154621225407180839476298628368035496429879296;
data[142]<=640'd1432108391621439505026886997447224277695550190362521311331009167475215864237658663636716821857020275584059608091812043003909209505308931123163491729408;
data[143]<=640'd1432108391621439505026886997365723278023620873331869727152474194724948003708818863349359636397631083540867698410506682259627063857046814088751761850368;
data[144]<=640'd1432108391621439505026886997865358389702177150605165303145258429402837446582954197638295636923873398044756134233409858196019054312570197228487975108608;
data[145]<=640'd1432108391621439505026886997865074693978380074121854890236161915340260594625376070520270905906096337945375461411509381279946242164821610597170840338432;
data[146]<=640'd1432108391621439505026886998854409262952676980504621109721009824267732975110142491754913744821047592131340536058964915344021645435596313560973708361728;
data[147]<=640'd1432108391621439505026886998851827008149193100032196504936387199730249542554028750995786366208166543904089351905520081125512928689697626404479748276224;
data[148]<=640'd1432108391621439505026886998851844660249461589263663137068926051993840052404754591566545789242465351085204514756844446676376195612999575383996222144512;
data[149]<=640'd1432108391621439505026886998851880003851417626235672409156543054723011927644083903878583113956520208122970877229942782243849384203947466329057474379776;
data[150]<=640'd1432108391621439505026886998851960689309465379937974215348640987936299799157058308259933202125717275149084196427410320986260374569061910111429653954560;
data[151]<=640'd1432108391621439505026886999182639977407932912318160474930286812633850667917497385985339999057114568437894464897525317349637161329206581616471477059584;
data[152]<=640'd1432108391621439505026886999182942584814920873430650423032694709628170154583606385661603819914208139368650191170835502616397517265060376598406542393344;
data[153]<=640'd1432108391621439505026886998027910362682132534108847785449568960627476270656738845839804216555704037225247595403564818688043503454028482857191008632832;
data[154]<=640'd1432108391621439505026886997529374725893571591274898906303286495872453939078611570843770547722574507543904434341396434297579741388017383966642400133120;
data[155]<=640'd1432108391621439505026886997197878397791758610023294126888758972915747772504473914776023068001049077871092589863193076052654946685102377569148978855936;
data[156]<=640'd1432108391621439505026886996940944456116278685118659163126484435799439642037184193056598196011954859360205143397155628336586548693470503394095768010752;
data[157]<=640'd1432108391621439505026886996868641420127256607431444208395909635239964769402726650831033115052207720387956190202354378611678955879848565437861870960640;
data[158]<=640'd1432108391621439505026886996868641420127256607431444208396822227357362619169374914499440516468358778228318529642639369532989718702142540282232032985088;
data[159]<=640'd1432108391621439505026886996868641420127256607431444208398647411592158318702671441836255319300660893909043208523209351375611244346730489970972357033984;
data[160]<=640'd1432108391621439505026886996868641420127256607431444208402297780061749717769264496509884924965265125270492566284349315060854295635906389348453005131776;
data[161]<=640'd1432108391621439505026886996868641420127256607431444208426285915719064625921161712936593762189807217074302631571840504992451489821919442400468675854336;
data[162]<=640'd1432108391621439505026886996868641420127256607431444208657823572933147652430778323663957321487561320571947609564146773027867885878219345772098355200000;
data[163]<=640'd1432108391621439505026886996868641420127256607431444208645308023894548569916744993354370102066061098761264097240238326107034567172473405049307561721856;
data[164]<=640'd1636695303852802729735721062055718605960824492694731914513886315868436735039865809623431264300745114147225121181134921005965207090773500786651179253760;
data[165]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[166]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[167]<=640'd0;
data[168]<=640'd0;
data[169]<=640'd0;
data[170]<=640'd0;
data[171]<=640'd0;
data[172]<=640'd0;
data[173]<=640'd0;
data[174]<=640'd0;
data[175]<=640'd0;
data[176]<=640'd0;
data[177]<=640'd0;
data[178]<=640'd0;
data[179]<=640'd0;
data[180]<=640'd0;
data[181]<=640'd0;
data[182]<=640'd0;
data[183]<=640'd0;
data[184]<=640'd0;
data[185]<=640'd0;
data[186]<=640'd0;
data[187]<=640'd0;
data[188]<=640'd0;
data[189]<=640'd0;
data[190]<=640'd0;
data[191]<=640'd0;
data[192]<=640'd0;
data[193]<=640'd0;
data[194]<=640'd0;
data[195]<=640'd0;
data[196]<=640'd0;
data[197]<=640'd0;
data[198]<=640'd0;
data[199]<=640'd0;
data[200]<=640'd0;
data[201]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[202]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[203]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
data[204]<=640'd716054195810719752513443498452396459210236663843313538401519604681591400367843758171127472313812864627914813743442211318145061348828617500555078533120;
data[205]<=640'd716054195810719752513443498454817318470943140646115962625272428313775499548621155214406215460569721773555602363407503836845190565799776724279529308160;
data[206]<=640'd716054195810719752513443498516942619248823106185030406280912270583849488969373445934094087849421263174083520826805540203121430985236360613379530817536;
data[207]<=640'd716054195810719752513443498599582180532793891087527193434379346215841788567102110100978117211933049057178062906913029171650412120303285071331498917888;
data[208]<=640'd716054195810719752513443498594424617992336026611211666968870954002199316658579354529295692867369532881627382597869581719349971971229802136622671593472;
data[209]<=640'd719250854131913053886533600199418131689862005089317237406482255616901057409693253883221885703094540644270681789158137926077829791260379425268454916096;
data[210]<=640'd719250854131913053886533600194252696136041023541124107418553862163745625290138930071407860819617322961628159615987519989479461988438978380253420847104;
data[211]<=640'd719250854131913053886533600235568680640991928671517968959610506117931398689067684309072729739544423062215444676152363935902008602495672201885211688960;
data[212]<=640'd719250854131913053886533600235568675715741154122208067558490423950219846832918682301737119959350190513594274448793891735661737391856151232077637877760;
data[213]<=640'd719250854131913053886533600225239676203393538111573318757610486752386221306288888436269676279733329536645641771258092934091961173976413368874128375808;
data[214]<=640'd719250854131913053886533600307872617950323321861066594978526246956876255626741627748851189993789995297173043015515455480511650259494123836374882713600;
data[215]<=640'd719250854131913053886533600307879552713146247752422720985957879825758128690770286753453603349680471749068284895889620869122121674450422788010950000640;
data[216]<=640'd719250854131913053886533600287250583136826368923567430364900071095864238114325089110345114188504565307363004439750059771172728865986096809377120911360;
data[217]<=640'd719250854131913053886533600452628053113446019681222594529592649591518440259905622526300521191210437794292736474222704759385310619852994709924566007808;
data[218]<=640'd719250854131913053886533600455018691079965798819946490039165802919367173676488081184535265352522253814883371034942450251574121912949457080286644797440;
data[219]<=640'd719250854131913053886533600493631396287031652315794431061150144112822713572253577970586053200371640249985797327237166447266698443808050098747551514624;
data[220]<=640'd719250854131913053886533600491210527245566033030350755199259089700643392914999387256865122443725751776485296416960598330508967462554632562602795859968;
data[221]<=640'd719250854131913053886533600741688765410367138197336776524538909213764127549917621357379057470538874102341314684378240570823765452772367529781906898944;
data[222]<=640'd719250854131913053886533600659056848096359181518336111276353217257447604762878349857744933017952609879191357030405975668036602788198934275890947817472;
data[223]<=640'd719250854131913053886533600659056828549345305112374006863474791664613750941342944173783993822872015798001615031024299660334132192674288574530249031680;
data[224]<=640'd719250854131913053886533601320112797301096740813384660574325534839813209736111440198833357407945074390547126805277598755827798055962467109777111515136;
data[225]<=640'd719250854131913053886533601320112954909271796563965936300147056171026435136870824635423675249048779498158873979389794969658073700651478371435005607936;
data[226]<=640'd719250854131913053886533601154848963019500243804848195180876919904993642146856118901572499785628353483924522515726971382205346834220604150518109962240;
data[227]<=640'd716054195810719752513443499425904900123006321892684327391627979833966398203541687810086025966492434445610482967791808411731173206438044431614669225984;
data[228]<=640'd716054195810719752513443500748016837703804356719440658621889048670187383705742252154792706093711491586733855110068319510099229844196759380564610383872;
data[229]<=640'd716054195810719752513443500748017152919778787986916839628238819076166832342626120149144509311646161009324757501601892866314905534279262675934774296576;
data[230]<=640'd716054195810719752513443500417489168524654615226286366532113576586219958341702119533547297296133204822806923134614207553653809644564894950407257718784;
data[231]<=640'd716054195810719752513443499756432805560279541931114698735649863252824271402368568143057938395255371826363848621175488615897430102674974581120177274880;
data[232]<=640'd818347651926401364867860531027859302980412393131277380521395508717963006741230473315177183548362701793830182762363954799343770380606623659043181297664;
data[233]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[234]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[235]<=640'd0;
data[236]<=640'd0;
data[237]<=640'd0;
data[238]<=640'd0;
data[239]<=640'd0;
data[240]<=640'd0;
data[241]<=640'd0;
data[242]<=640'd0;
data[243]<=640'd0;
data[244]<=640'd0;
data[245]<=640'd0;
data[246]<=640'd0;
data[247]<=640'd0;
data[248]<=640'd0;
data[249]<=640'd0;
data[250]<=640'd0;
data[251]<=640'd0;
data[252]<=640'd0;
data[253]<=640'd0;
data[254]<=640'd0;
data[255]<=640'd0;
data[256]<=640'd0;
data[257]<=640'd0;
data[258]<=640'd0;
data[259]<=640'd0;
data[260]<=640'd0;
data[261]<=640'd0;
data[262]<=640'd0;
data[263]<=640'd0;
data[264]<=640'd0;
data[265]<=640'd0;
data[266]<=640'd0;
data[267]<=640'd0;
data[268]<=640'd0;
data[269]<=640'd0;
data[270]<=640'd0;
data[271]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[272]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[273]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[274]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[275]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[276]<=640'd716054195810719752513443498436902329509616069993710626904859931137792284335040089646996829001874510964265422620294556570204156201562945562670748663808;
data[277]<=640'd716054195810719752513443498475636077680919698838549414484905109252737871227478442339456719349984225294518040539739236869406223673101493142261961064448;
data[278]<=640'd716054195810719752513443498764203131989230876044265778420883288506903374851972497345429589616096064986448387994971887726721704494713925516264338358272;
data[279]<=640'd716054195810719752513443501075962335346535790933735072534116409542307789640129758881856114652118974840552957684284325086262295903437522520986112491520;
data[280]<=640'd716054195810719752513443508936330964243310997934299320101161945139223999366914197463078394669438236193084646203335782881574369898171715801520548085760;
data[281]<=640'd716054195810719752513443519265330476590982933239308044822392414689331103834041171381277090042968167159521430263441464572718312641489842287878613237760;
data[282]<=640'd716054195810719752513443518284075522917920092488719067374528189671023665650908402235286529253574501650522280565529526920176121880409916046746893418496;
data[283]<=640'd716054195810719752513443498452396459210462123931259826391396994818883176722471823695822671021400764561181905809853213728717576452673555296046144290816;
data[284]<=640'd716054195810719752513443498449814209332375215341603907219393982944553470929642600182992011664860116939165064615223568375437438621237652124073396797440;
data[285]<=640'd716054195810719752513443498449814209332675828792198959741552492891738828164790680447610376885677107245592361074099645100643052151091383788153310543872;
data[286]<=640'd716054195810719752513443498470472208357296532456069495355220800717315295409424067509323404103846287738224339862431283562756427942171383677257546465280;
data[287]<=640'd716054195810719752513443498470472245296789193897524885153498362561344464051193620122991184124157306732063564090470508834172320742291097521131574263808;
data[288]<=640'd716054195810719752513443498465307865602658693133458516961066248897713390654644228328779303032332226412839833220615876792369138435907871673042136465408;
data[289]<=640'd716054195810719752513443498465307988733919250055530179090002669739408021728330603250509907113241755854240066293028306935115618068248898069690446774272;
data[290]<=640'd716054195810719752513443498506624260127372139531325437036200070719626186885047975754102994146508111398543647493240509431258382984310276384408731648000;
data[291]<=640'd716054195810719752513443498496295814704383881295676062170550081767161153415043803623859074324190431956418429410889029815587060889478067374352666460160;
data[292]<=640'd716054195810719752513443498496295662022812323782761870587916157253896573255094066940805254400867231041917333922361192552993492372979840399978975461376;
data[293]<=640'd716054195810719752513443498496296951822858908309987685876216829396839914528060514285023767266729571651450982271288846974036962317272084211347933364224;
data[294]<=640'd716054195810719752513443498578931741769841824547066520502883281936589987764275614399516277332028591823409897256980011086917888149978517610143791710208;
data[295]<=640'd716054195810719752513443498558278771426188544946502498052319976344874161232557918827616281603359197962840568093369515775553924105436891689389884702720;
data[296]<=640'd716054195810719752513443498558278475911141483705513398365213768819594491263525670780384220844274925653013265520827590983322030889469131576425356197888;
data[297]<=640'd716054195810719752513443498558272486806201980287395889563734169743938988323341750211228189541787287895625183229269806637466046417796349828133076074496;
data[298]<=640'd716054195810719752513443498723536479927252173067244483859558766269051291626509507707747657120232923303169422018570654865081928527056940318848807075840;
data[299]<=640'd716054195810719752513443498723536481158874883499457587595962191555952092861975347895139843247036184052869221329693412692250148544623692447520611368960;
data[300]<=640'd716054195810719752513443498682221130472412500164015030748316599426718847179850664840786266601969270520428233878680726559662575733659658746413042368512;
data[301]<=640'd716054195810719752513443498682219217626935783688236265452195436977737437282247049624759838328005796649578242945000593351105964490429237779900150054912;
data[302]<=640'd818347651926401364867860531027860544143832906622819285070802166648325145936293367879823861257253301713640055421807465536124401416969883210374893797376;
data[303]<=640'd818347651926401364867860531027859302980412246347505941203204878388585547550201790102400479621947948184075711318110122128264813958505529454328717246464;
data[304]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[305]<=640'd0;
data[306]<=640'd0;
data[307]<=640'd0;
data[308]<=640'd0;
data[309]<=640'd0;
data[310]<=640'd0;
data[311]<=640'd0;
data[312]<=640'd0;
data[313]<=640'd0;
data[314]<=640'd0;
data[315]<=640'd0;
data[316]<=640'd0;
data[317]<=640'd0;
data[318]<=640'd0;
data[319]<=640'd0;
data[320]<=640'd0;
data[321]<=640'd0;
data[322]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[323]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[324]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[325]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[326]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[327]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[328]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[329]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[330]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[331]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[332]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[333]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[334]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[335]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[336]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[337]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[338]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[339]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[340]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[341]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[342]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[343]<=640'd398353494612575324017191154914352288844846764696638810260114131509605650307885529420329033517687589677374404780947210779386712874022118574019139283960076830011772872351155913515597824;
data[344]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[345]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[346]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[347]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[348]<=640'd398353494612575324017191154914352186551390649015026455843081537971012733523942897776476074197443525535126815153878457074366752531570804226482521018768785698054402230421841660119875584;
data[349]<=640'd265568996408383549344794103276235029718992369583268475043220513910041109088511359234064155610167347940571714494382458401709398254602728763359583467446130040472067320563817398958817280;
data[350]<=640'd265568996408383549344794103276235029718992369583268475043220542153399150664074058595680099393109723421728823564014629987046110417936094572560149729192181541979598650754760850884526080;
data[351]<=640'd265568996903044352291003171397240071758286749653531173245644265870947140976898850940200584448743909205504922481436351689200150496414012795173930077975219068851482267557512510571544576;
data[352]<=640'd265568996903044352291003171397240071758286749653531173245644265558252819896327359178219133617954960188615259508155358968348673864571206520720809202410771322490992271206384922743799808;
data[353]<=640'd398353495107236126963400223035357228590685029085289154045505297848885066685838825189461651410739422896187426297242838665317545949164137665328712269515090178962203775974916756376387584;
data[354]<=640'd265568996903044352291003171397240071758286749653531173245644338184030641034303117242229689877502164522971427564103021196670092171290393849036582324453145440167845741598409794485485568;
data[355]<=640'd265568996903044352291003171397240071758286749653531173245644327855031128611515395969790338572991288106889471371187128308966430146066594692641115002204262128778152049673123406473592832;
data[356]<=640'd265568996903044352291003171397240071758286749653531173245644307197032103916246678722436962548896293469243128737399025663691577820885618557911557965041435887675500562447747624493645824;
data[357]<=640'd265568997892365958183421307639250155836875509794056569650491832117276525850132101038814803999664947352685383330305512689261723771658093458695782166283893464620766319316229012867514368;
data[358]<=640'd265568996903044352291003171397240071758286749653531173245644472461063818920267927613494590438064006976687019289681191333776707214442910372948086204241920481272126874592137966946091008;
data[359]<=640'd265568996903044352291003171397240071758286749653531173245644431205607106415498351048945982500342200140279227042640518206448955333946888070244009063416593263508288873275499490247180288;
data[360]<=640'd265568996903044352291003171397240071758286749653531173245644431770484387098227638060986536861113849285553400473186921434630770436779591819154968957088195460873412620290859285490958336;
data[361]<=640'd265568996903044352291003171397240071758286749653531173245644766756845724655747473510255706594824695543368075391008313367673797349528654530894869267351649187414430494941395726620426240;
data[362]<=640'd265568996903044352291003171397240071758286749653531173245644843659480909080866790552231080676368793600226952876822552707429198519299934820975122398871077385613727999725727203415031808;
data[363]<=640'd398353495107236126963400223035357228590685029085289154045505876272876844122221199281299545126859726022122334059205504615661116760422648465263434564713455934430047793314326588816359424;
data[364]<=640'd265568996903044352291003171397240071758286749653531173245645484702994982139725872965258139836562807659282043279684631898945903919829267023699733195241668281122035439496027543105961984;
data[365]<=640'd265568996903044352291003171397240071758286749653531173245645340097000579162458233375088372050565688726667460553454196218566568069607323140557732441880137923280415860907149770532847616;
data[366]<=640'd265568996903044352291003171397240071758286749653531173245645174833028082302793242040816850208002287043364119848697241519436780164328392567484269535213354364233174627674152840600748032;
data[367]<=640'd265568997892365958183421307639250155836875509794056569650493856601337324502862867062672605271651108427048876329190094906304104597697945171522775673170267909795562382300825067007770624;
data[368]<=640'd398353495107236126963400223035357228590685029085289154045507531495314049022707758805221808527669066460065147963112017655568023638169995171863509723114198942463964854009681611778424832;
data[369]<=640'd265568996903044352291003171397240071758286749653531173245646166982367429213654653607639590747946535849447754254214342759981391193928366993523644887359573947682335248412627898218840064;
data[370]<=640'd265568996903044352291003171397240071758286749653531173245646168838908693948757269410713320960433747478933289273331719673164322356616834544702525663131062790607969032125819749335564288;
data[371]<=640'd265568996903044352291003171397240071758286749653531173245648820651452948170946773728445373595175963805733747734958428812846622296264991660556917029629575456997943970807968902695354368;
data[372]<=640'd265568997892365958183421307639250155836875509794056569650496830070743775665005331346202969610616535024674669991064294781277940123279233337905270013843241342490693245972345363328139264;
data[373]<=640'd265568996903044352291003171397240174051742865335143527662682054913947799261606721964401616714338507026402603841286661204148291631905629204376219183101830592291163931199020767880675328;
data[374]<=640'd265568996903044352291003171397240174051742865335143527662679255747514454022224283900141070411542534696719932584147492194075207522237814138723162892139430987789628858278988575806586880;
data[375]<=640'd265568996903044352291003171397240174051742865335143527662676776787630872528466918948602142292013070382638162388580928377582346718311671832780261709203522302229601390475521153055064064;
data[376]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[377]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[378]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[379]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[380]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[381]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[382]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[383]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[384]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[385]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[386]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[387]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[388]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[389]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[390]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[391]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[392]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[393]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[394]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[395]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[396]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[397]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[398]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[399]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[400]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[401]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[402]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[403]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[404]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[405]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083711154225492614732989228270490262743671417864192;
data[406]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083756826325883777643510875830043263955216103374848;
data[407]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083733993150393632101736882977413894943200384122880;
data[408]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260510356823990064450203354978959320258094768848896;
data[409]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841306678842167437339742438259765413224120320;
data[410]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841295784489368253867537777416344549361451008;
data[411]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083866058175805198939743815208226653779662768963584;
data[412]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934544014703162186716804046514368768030868556417597440;
data[413]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260686614913495185286957388911191037195542417375232;
data[414]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083871185952298368884399164504508543769418921934848;
data[415]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986330444476161582688175652864;
data[416]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[417]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[418]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[419]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[420]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[421]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[422]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[423]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[424]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[425]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[426]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[427]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[428]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[429]<=640'd398353496343888134328922893337869117634725168541193386108065983048744062545919757800094946891136771680368312041868575743622909878699085669704398453847763599671125628542792319314690048;
data[430]<=640'd531137992816767098689588206552468627329593117540961209779768774219776665041523081944630313929275862236827838496002843258316710966147798256686047195211381820739689719850535202106376192;
data[431]<=640'd464745747548292448942947204772883260336491728765709340960903687623617040888630979714838395224460056055998811059991606943419003558340812870361086397939032316978126257926111479799480320;
data[432]<=640'd1731312810311731738423517647137530330245919443708482879398441392650280575745723070192214807428701314927183699982112975375459555240147258469772823085713252175416247405040893952;
data[433]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[434]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[435]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[436]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[437]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[438]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[439]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[440]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[441]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[442]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[443]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[444]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[445]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[446]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[447]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[448]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[449]<=640'd741991204419313602181507563058941570105394047303635519742189168278691675319595601510949203183729134968793014278048418018054095102920253629902638465305679503749820316446097408;
data[450]<=640'd989321605892418136242010084078576565810250724560193525292073344815707069964632683637707560663098643350035920994610962411690368371714661765920491625786887328011429868730318848;
data[451]<=640'd1799565517869652802850553672994603778697120433756232925976991265676467694158133288870091067319688664337182830767822544995324267558345195980337572361199321983483904;
data[452]<=640'd0;
data[453]<=640'd0;
data[454]<=640'd0;
data[455]<=640'd0;
data[456]<=640'd0;
data[457]<=640'd0;
data[458]<=640'd0;
data[459]<=640'd0;
data[460]<=640'd0;
data[461]<=640'd0;
data[462]<=640'd0;
data[463]<=640'd0;
data[464]<=640'd0;
data[465]<=640'd0;
data[466]<=640'd0;
data[467]<=640'd0;
data[468]<=640'd0;
data[469]<=640'd0;
data[470]<=640'd0;
data[471]<=640'd0;
data[472]<=640'd0;
data[473]<=640'd0;
data[474]<=640'd0;
data[475]<=640'd0;
data[476]<=640'd0;
data[477]<=640'd0;
data[478]<=640'd0;
data[479]<=640'd0;
end
else if (choise == 2) begin
data[0]<=640'd0;
data[1]<=640'd0;
data[2]<=640'd0;
data[3]<=640'd0;
data[4]<=640'd0;
data[5]<=640'd0;
data[6]<=640'd0;
data[7]<=640'd0;
data[8]<=640'd0;
data[9]<=640'd0;
data[10]<=640'd0;
data[11]<=640'd0;
data[12]<=640'd0;
data[13]<=640'd0;
data[14]<=640'd0;
data[15]<=640'd0;
data[16]<=640'd0;
data[17]<=640'd0;
data[18]<=640'd0;
data[19]<=640'd0;
data[20]<=640'd0;
data[21]<=640'd0;
data[22]<=640'd0;
data[23]<=640'd0;
data[24]<=640'd0;
data[25]<=640'd0;
data[26]<=640'd0;
data[27]<=640'd0;
data[28]<=640'd0;
data[29]<=640'd0;
data[30]<=640'd0;
data[31]<=640'd85070591732710495944414412407740301312;
data[32]<=640'd730750818665451459101842416358132502628711530496;
data[33]<=640'd27021597764222976;
data[34]<=640'd9007199254740992;
data[35]<=640'd9007199254740992;
data[36]<=640'd9007199254740992;
data[37]<=640'd9007199254740992;
data[38]<=640'd9007199254740992;
data[39]<=640'd9007199254740992;
data[40]<=640'd13510798882111488;
data[41]<=640'd9007199254740992;
data[42]<=640'd9007199254740992;
data[43]<=640'd9007199254740992;
data[44]<=640'd9007199254740992;
data[45]<=640'd13510798882111488;
data[46]<=640'd9007199254740992;
data[47]<=640'd9007199254740992;
data[48]<=640'd9007199254740992;
data[49]<=640'd13510798882111488;
data[50]<=640'd31525197391593472;
data[51]<=640'd309787241346054520360140800;
data[52]<=640'd599375721660670508425266668362373856774380817170532873411752110287376594018075499955962254745047801101257078721539110295345450208080468874490806272;
data[53]<=640'd5027929472167778066878457916438579271401010308215785621888644634346722099039006813346457612736872842782101791232293722601083851606530876499670384477470720;
data[54]<=640'd26396628205467732864788082285642163171681467387598851022504789516166031859271295734080499794632056350026575515206137239670386077067062433013666803051659264;
data[55]<=640'd107052979177370224261959331447169757995624348293019147030047829383530188356005728063506518606159218349527795023329677542352008354006734679382389176714395648;
data[56]<=640'd214315455403593848371243628535063509913572769065503325629120859826805569962864356697324533626196254014778770029289013968377661500181271326886728884677509120;
data[57]<=640'd428840407856041074259963789741753073154462173194139026648524031365156604373179187965892171529647976321944478726877311152888398901532830347995215140384407552;
data[58]<=640'd857890312710984452973429432205287855794666022103459363145609269421919230326598971951740951076827667545097005016360117896252295914307608837212705991216332800;
data[59]<=640'd1715990122520767163402835295025441171969567992656791332698788381890886667082526282063613182540215233834685701369746996036155842454675129901135972923267350528;
data[60]<=640'd3381910457608045116620999402357853392069290396874125430328045293723256668427299865470942285888501138062814744645993448611444427055806175678689141383990607872;
data[61]<=640'd6760678458734064500004395559042319423859994262652645444346415197021551412634851879054371547607344496682524987027586199293328324311640523138232093438226989056;
data[62]<=640'd13518213642638457425626434681613824247268059382700472661371176154298941598148001792901619029354125148973649014067957618735459638875554094018914426032008200192;
data[63]<=640'd13303689508433767673001792403097267332445570694662408114543717372905665493958789517438273337383157632243321737455198609118372135649314003991232408626193760256;
data[64]<=640'd26604027063486494151856852108440019966858802187707887285518607084327113815165657061281383825521489522527025728247401310676293068991128914079610415427673391104;
data[65]<=640'd54066572828686917512538848091696728615772215835780101081038941672982135750213955630549554187526714626306345586352280791600468548118337364405108883342695071744;
data[66]<=640'd108126854402215468636948495822802328610646555176645496568601164575687211790167285726112387578570729443792281568925608496419361685686955605409517285680324018176;
data[67]<=640'd106410661329377119006977893772893853047864231581297737945232268808300772200366709756376036593409518210486072502430351275254099497567078879082869518791243464704;
data[68]<=640'd216247436575855479282092410736678649095590945920787579121648876487916844005673158738319991589732162304852207301197122119583818767818967446770323958965500641280;
data[69]<=640'd212814617933244944225846956985053715385389454010758270613221946629202400863949106570233714202028220831395569769179299962980594675440578057599903261196493520896;
data[70]<=640'd425630075491580350373514556489764094002022545108418790299028410609512909024529356069086987000409094756423964141442302784669197120254938147435314767835038744576;
data[71]<=640'd864977176477493792998426720553126075865707973051461377546367259004900087853513061839282910684749462706454618560081417516813094727567860441403240096422265094144;
data[72]<=640'd851247682632341467128970141392075156053575187939118035919251798845312188512943540402250903746277609282808142921882505770245391633396799966707883547220447854592;
data[73]<=640'd1729955184390208237472303383221228712183658530661859015675224928698743183157140205290275958981656649640543026924220237830657450719240773284034815281766284132352;
data[74]<=640'd1702495365258689079671238639778692186686648698691038037051379820481306262388471864585215024917390711291478313796939795069715334066961525319969474466567994474496;
data[75]<=640'd3459883972158554305902524366150836688105814640052773469618604938651459850491363095953710892695995849384108774563596257108611723471560113782663469689111389929472;
data[76]<=640'd3404966402678380287026472699061892275557714108338375202607199483365135647893772515601448216130947937129818071330403331790953794098718246683046836199909150949376;
data[77]<=640'd6919769620281112346282473663417035300574804215453964264447298784452164613972549122915290026490312135640287871664655176173607558561847291296195597047089902649344;
data[78]<=640'd6809932805344772864421133650764320560533861927265129952552077886232105511571101450500741662581779928543593774435373931650172041152181291712486836710752275922944;
data[79]<=640'd13839485504582804636771634314557442765540704517288645763211024595086836483792384167084161877332950073509926851413873715336011710023323021165928452172413373775872;
data[80]<=640'd13619811979458625123224703741313646734349949348047649061338701020815318781929897902843165232488609907086914327981229207162956470717094728387741441325879816880128;
data[81]<=640'd27678971009140035495573996324079679547060880019621936630943123616759766761141886885221954464300421961469106309459060756254840548257620172840974207485516475006976;
data[82]<=640'd27239623539897679053327564100571767080268538237049088531596804344288460452819900738111875815959250704898749886308357836242488687851363195978447168975123953745920;
data[83]<=640'd55357834755792656445893429784966008765323002970073268929816810071248050828911928509004133547621889284623934433607299484814503444967508689819300071169627483275264;
data[84]<=640'd54479247079796955661475752410167943692920068694349925510592349617495011916437736470975248442430863494517913342821690832962759812414814875610540376595600097935360;
data[85]<=640'd110715669511586911227044760910989549664951290921252942767736421845620006903796688988886746286888562537833446547416159306317038729986015682962372443556378803437568;
data[86]<=640'd108958279634617483897186059353955721834531173292492643743446586046970229497852579626815538309591923960744126037655557682374053725383735175296355788649654040657920;
data[87]<=640'd108958276282663903076283488369549075760180252722079693234698334086877633526618490491310064159152584231270217074212862956664341061242741187353202903905637178015744;
data[88]<=640'd221431335671170693240215314621644771431426395490521791277898172646833623334842425363648422135228700058062154206682413788871748700324389950795583538713360416636928;
data[89]<=640'd217916552565331002823165766959398391001306435154144838499707258298812106106143536212746440113533544594240287378617390005937186876393157600823930063484681833152512;
data[90]<=640'd442862242292490821964359011659308181960156777221913368692767379022222992390025038628709715690211444402007032171733189041754440386983041800259773752932296824979456;
data[91]<=640'd442862228884679695448036652215884974418818052233948439596294440625308896041677152899905542243931370874668803798369585865243004234553139213729170333811226439581696;
data[92]<=640'd435833105130508562534745063552623256078125856084596639737079105219936424717994818075581101639306710098286409836474796876868486384501888739015930737911622812041216;
data[93]<=640'd435833078314886309308436457572871538053355971474607200970256890968555190777274628892512546854519477174740741143016318386965325376872929856817777546809377032241152;
data[94]<=640'd421773972706900460565300364381239083639546980409929178366340363577876513135139219757465394741596352353179657050576974825036112800830974047350341605563815455358976;
data[95]<=640'd421773490025814980266866852072168080722746520326731594415381246511774577959324591550086354122775601042723754080244766925928918731942453508047105353713736589770752;
data[96]<=640'd168709267295369864355395194106365450110326787925898158555921256322683905591083810756201579645300549095178113289751200261547810419468161304768314266015640158470144;
data[97]<=640'd9007199271518208;
data[98]<=640'd9007199271518208;
data[99]<=640'd9007199305072640;
data[100]<=640'd13510798898888704;
data[101]<=640'd9007199271518208;
data[102]<=640'd9007199271518208;
data[103]<=640'd9007199271518208;
data[104]<=640'd9007199305072640;
data[105]<=640'd13510798898888704;
data[106]<=640'd9007199271518208;
data[107]<=640'd9007199271518208;
data[108]<=640'd9007199271518208;
data[109]<=640'd9007199271518208;
data[110]<=640'd13510798898888704;
data[111]<=640'd9007199271518208;
data[112]<=640'd9007199271518208;
data[113]<=640'd9007199271518208;
data[114]<=640'd9007199305072640;
data[115]<=640'd13510798898888704;
data[116]<=640'd9007199271518208;
data[117]<=640'd9007199271518208;
data[118]<=640'd9007199271518208;
data[119]<=640'd9007199305072640;
data[120]<=640'd9007199271518208;
data[121]<=640'd9007199271518208;
data[122]<=640'd9007199271518208;
data[123]<=640'd9007199271518208;
data[124]<=640'd9007199271518208;
data[125]<=640'd13510798898888704;
data[126]<=640'd9007199271518208;
data[127]<=640'd9007199271518208;
data[128]<=640'd9007199271518208;
data[129]<=640'd533996758980227548388856843498274930307712532674261077271556721709290300914980308412090940391424;
data[130]<=640'd1868988656430796558311506037023396764362175874785403194374430124751192900551531866420075563057152;
data[131]<=640'd70608395103938906748405908848113786735498346477469127413701232021435384158860502965062554256599959879843061883878768640;
data[132]<=640'd320259506364294327037405639924244233692028483547307954462621785835688912818792645285933467907937828686853293558248505344;
data[133]<=640'd1636695303852802729735721062057007209171471377742890289643062904937418624395482718595003351178232432600793374821907689755208590573672079544628279246848;
data[134]<=640'd1636695303852802729735721062058147030406720677237543099851066895318485373478903061535747386712734283593220464541437540325981490295668695865160609300480;
data[135]<=640'd1636695303852802729735721062065404564732046969152611200271195788852249740197418431205925877357108034363812204308885191990930668944454828233263325118464;
data[136]<=640'd1432108391621439505026886996886717169273864967559035645802998680124266543704676409646449470163531041179254364961423359278795446832131342830488728371200;
data[137]<=640'd1432108391621439505026886996904792918420473327686627080007019763244601044180741872875958218823407205924272963993675377937932973822672338671949406273536;
data[138]<=640'd1432108391621439505026886996940944416713690047941809952687036001327029501520034157640508399872311787975085208710858581108289465131830540530627962208256;
data[139]<=640'd1432108391621439505026886997013247413300123488452175689503120333808321972122134470033220033847614419284429732306322481390539143083906703564612258758656;
data[140]<=640'd1432108391621439505026886996992589414275428219734928335071630492107686374016258216053810355123933847131021312988412579121760328376010588614750415880192;
data[141]<=640'd1432108391621439505026886997116552548875351926674048803359290596818587304240900274827643548059306807017147154621225407180839476298628368035496429879296;
data[142]<=640'd1432108391621439505026886997447224277695550190362521311331009167475215864237658663636716821857020275584059608091812043003909209505308931123163491729408;
data[143]<=640'd1432108391621439505026886997365723278023620873331869727152474194724948003708818863349359636397631083540867698410506682259627063857046814088751761850368;
data[144]<=640'd1432108391621439505026886997865358389702177150605165303145258429402837446582954197638295636923873398044756134233409858196019054312570197228487975108608;
data[145]<=640'd1432108391621439505026886997865074693978380074121854890236161915340260594625376070520270905906096337945375461411509381279946242164821610597170840338432;
data[146]<=640'd1432108391621439505026886998854409262952676980504621109721009824267732975110142491754913744821047592131340536058964915344021645435596313560973708361728;
data[147]<=640'd1432108391621439505026886998851827008149193100032196504936387199730249542554028750995786366208166543904089351905520081125512928689697626404479748276224;
data[148]<=640'd1432108391621439505026886998851844660249461589263663137068926051993840052404754591566545789242465351085204514756844446676376195612999575383996222144512;
data[149]<=640'd1432108391621439505026886998851880003851417626235672409156543054723011927644083903878583113956520208122970877229942782243849384203947466329057474379776;
data[150]<=640'd1432108391621439505026886998851960689309465379937974215348640987936299799157058308259933202125717275149084196427410320986260374569061910111429653954560;
data[151]<=640'd1432108391621439505026886999182639977407932912318160474930286812633850667917497385985339999057114568437894464897525317349637161329206581616471477059584;
data[152]<=640'd1432108391621439505026886999182942584814920873430650423032694709628170154583606385661603819914208139368650191170835502616397517265060376598406542393344;
data[153]<=640'd1432108391621439505026886998027910362682132534108847785449568960627476270656738845839804216555704037225247595403564818688043503454028482857191008632832;
data[154]<=640'd1432108391621439505026886997529374725893571591274898906303286495872453939078611570843770547722574507543904434341396434297579741388017383966642400133120;
data[155]<=640'd1432108391621439505026886997197878397791758610023294126888758972915747772504473914776023068001049077871092589863193076052654946685102377569148978855936;
data[156]<=640'd1432108391621439505026886996940944456116278685118659163126484435799439642037184193056598196011954859360205143397155628336586548693470503394095768010752;
data[157]<=640'd1432108391621439505026886996868641420127256607431444208395909635239964769402726650831033115052207720387956190202354378611678955879848565437861870960640;
data[158]<=640'd1432108391621439505026886996868641420127256607431444208396822227357362619169374914499440516468358778228318529642639369532989718702142540282232032985088;
data[159]<=640'd1432108391621439505026886996868641420127256607431444208398647411592158318702671441836255319300660893909043208523209351375611244346730489970972357033984;
data[160]<=640'd1432108391621439505026886996868641420127256607431444208402297780061749717769264496509884924965265125270492566284349315060854295635906389348453005131776;
data[161]<=640'd1432108391621439505026886996868641420127256607431444208426285915719064625921161712936593762189807217074302631571840504992451489821919442400468675854336;
data[162]<=640'd1432108391621439505026886996868641420127256607431444208657823572933147652430778323663957321487561320571947609564146773027867885878219345772098355200000;
data[163]<=640'd1432108391621439505026886996868641420127256607431444208645308023894548569916744993354370102066061098761264097240238326107034567172473405049307561721856;
data[164]<=640'd1636695303852802729735721062055718605960824492694731914513886315868436735039865809623431264300745114147225121181134921005965207090773500786651179253760;
data[165]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[166]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[167]<=640'd0;
data[168]<=640'd0;
data[169]<=640'd0;
data[170]<=640'd0;
data[171]<=640'd0;
data[172]<=640'd0;
data[173]<=640'd0;
data[174]<=640'd0;
data[175]<=640'd0;
data[176]<=640'd0;
data[177]<=640'd0;
data[178]<=640'd0;
data[179]<=640'd0;
data[180]<=640'd0;
data[181]<=640'd0;
data[182]<=640'd0;
data[183]<=640'd0;
data[184]<=640'd0;
data[185]<=640'd0;
data[186]<=640'd0;
data[187]<=640'd0;
data[188]<=640'd0;
data[189]<=640'd0;
data[190]<=640'd0;
data[191]<=640'd0;
data[192]<=640'd0;
data[193]<=640'd0;
data[194]<=640'd0;
data[195]<=640'd0;
data[196]<=640'd0;
data[197]<=640'd0;
data[198]<=640'd0;
data[199]<=640'd0;
data[200]<=640'd0;
data[201]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[202]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[203]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
data[204]<=640'd716054195810719752513443498452396459210236663843313538401519604681591400367843758171127472313812864627914813743442211318145061348828617500555078533120;
data[205]<=640'd716054195810719752513443498454817318470943140646115962625272428313775499548621155214406215460569721773555602363407503836845190565799776724279529308160;
data[206]<=640'd716054195810719752513443498516942619248823106185030406280912270583849488969373445934094087849421263174083520826805540203121430985236360613379530817536;
data[207]<=640'd716054195810719752513443498599582180532793891087527193434379346215841788567102110100978117211933049057178062906913029171650412120303285071331498917888;
data[208]<=640'd716054195810719752513443498594424617992336026611211666968870954002199316658579354529295692867369532881627382597869581719349971971229802136622671593472;
data[209]<=640'd716054195810719752513443498470474108272331322421689801733046036933826550285750168652928145848503239957568531354763767237227511749508443218334678253568;
data[210]<=640'd716054195810719752513443498465308672718510340873496671745117643480671118166195844841114120965026022274926009181593149300629143946687042173319644184576;
data[211]<=640'd716054195810719752513443498506624657223461246003890533286174287434856891565124599078778989884953122375513294241757993247051690560743735994951435026432;
data[212]<=640'd716054195810719752513443498506624652298210471454580631885054205267145339708975597071443380104758889826892124014399521046811419350104215025143861215232;
data[213]<=640'd716054195810719752513443498496295652785862855443945883084174268069311714182345803205975936425142028849943491336863722245241643132224477161940351713280;
data[214]<=640'd716054195810719752513443498578928594532792639193439159305090028273801748502798542518557450139198694610470892581121084791661332217742187629441106051072;
data[215]<=640'd716054195810719752513443498578935529295615565084795285312521661142683621566827201523159863495089171062366134461495250180271803632698486581077173338112;
data[216]<=640'd716054195810719752513443498558306559719295686255939994691463852412789730990382003880051374333913264620660854005355689082322410824234160602443344248832;
data[217]<=640'd716054195810719752513443498723684029695915337013595158856156430908443933135962537296006781336619137107590586039828334070534992578101058502990789345280;
data[218]<=640'd716054195810719752513443498726074667662435116152319054365729584236292666552544995954241525497930953128181220600548079562723803871197520873352868134912;
data[219]<=640'd716054195810719752513443498764687372869500969648166995387713925429748206448310492740292313345780339563283646892842795758416380402056113891813774852096;
data[220]<=640'd716054195810719752513443498762266503828035350362723319525822871017568885791056302026571382589134451089783145982566227641658649420802696355669019197440;
data[221]<=640'd716054195810719752513443499012744741992836455529709340851102690530689620425974536127085317615947573415639164249983869881973447411020431322848130236416;
data[222]<=640'd716054195810719752513443498930112824678828498850708675602916998574373097638935264627451193163361309192489206596011604979186284746446998068957171154944;
data[223]<=640'd716054195810719752513443498930112805131814622444746571190038572981539243817399858943490253968280715111299464596629928971483814150922352367596472369152;
data[224]<=640'd716054195810719752513443499591168773883566058145757224900889316156738702612168354968539617553353773703844976370883228066977480014210530902843334852608;
data[225]<=640'd716054195810719752513443499591168931491741113896338500626710837487951928012927739405129935394457478811456723544995424280807755658899542164501228945408;
data[226]<=640'd716054195810719752513443499425904939601969561137220759507440701221919135022913033671278759931037052797222372081332600693355028792468667943584333299712;
data[227]<=640'd716054195810719752513443499425904900123006321892684327391627979833966398203541687810086025966492434445610482967791808411731173206438044431614669225984;
data[228]<=640'd716054195810719752513443500748016837703804356719440658621889048670187383705742252154792706093711491586733855110068319510099229844196759380564610383872;
data[229]<=640'd716054195810719752513443500748017152919778787986916839628238819076166832342626120149144509311646161009324757501601892866314905534279262675934774296576;
data[230]<=640'd716054195810719752513443500417489168524654615226286366532113576586219958341702119533547297296133204822806923134614207553653809644564894950407257718784;
data[231]<=640'd716054195810719752513443499756432805560279541931114698735649863252824271402368568143057938395255371826363848621175488615897430102674974581120177274880;
data[232]<=640'd818347651926401364867860531027859302980412393131277380521395508717963006741230473315177183548362701793830182762363954799343770380606623659043181297664;
data[233]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[234]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[235]<=640'd0;
data[236]<=640'd0;
data[237]<=640'd0;
data[238]<=640'd0;
data[239]<=640'd0;
data[240]<=640'd0;
data[241]<=640'd0;
data[242]<=640'd0;
data[243]<=640'd0;
data[244]<=640'd0;
data[245]<=640'd0;
data[246]<=640'd0;
data[247]<=640'd0;
data[248]<=640'd0;
data[249]<=640'd0;
data[250]<=640'd0;
data[251]<=640'd0;
data[252]<=640'd0;
data[253]<=640'd0;
data[254]<=640'd0;
data[255]<=640'd0;
data[256]<=640'd0;
data[257]<=640'd0;
data[258]<=640'd0;
data[259]<=640'd0;
data[260]<=640'd0;
data[261]<=640'd0;
data[262]<=640'd0;
data[263]<=640'd0;
data[264]<=640'd0;
data[265]<=640'd0;
data[266]<=640'd0;
data[267]<=640'd0;
data[268]<=640'd0;
data[269]<=640'd0;
data[270]<=640'd0;
data[271]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[272]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[273]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[274]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[275]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[276]<=640'd716054195810719752513443498436902329509616069993710626904859931137792284335040089646996829001874510964265422620294556570204156201562945562670748663808;
data[277]<=640'd716054195810719752513443498475636077680919698838549414484905109252737871227478442339456719349984225294518040539739236869406223673101493142261961064448;
data[278]<=640'd716054195810719752513443498764203131989230876044265778420883288506903374851972497345429589616096064986448387994971887726721704494713925516264338358272;
data[279]<=640'd719250854131913053886533602804906358764066473601362508207552628225382296764072844112149854506710275527255108118678695775112613945189458727919889154048;
data[280]<=640'd719250854131913053886533610665274987660841680601926755774598163822298506490857282693372134524029536879786796637730153570424687939923652008454324748288;
data[281]<=640'd719250854131913053886533620994274500008513615906935480495828633372405610957984256611570829897559467846223580697835835261568630683241778494812389900288;
data[282]<=640'd719250854131913053886533620013019546335450775156346503047964408354098172774851487465580269108165802337224430999923897609026439922161852253680670081024;
data[283]<=640'd719250854131913053886533600181340482627992806598887262064833213501957683846414908926116410875992065247884056244247584417567894494425491502979920953344;
data[284]<=640'd719250854131913053886533600178758232749905898009231342892830201627627978053585685413285751519451417625867215049617939064287756662989588331007173459968;
data[285]<=640'd719250854131913053886533600178758232750206511459826395414988711574813335288733765677904116740268407932294511508494015789493370192843319995087087206400;
data[286]<=640'd719250854131913053886533600199416231774827215123696931028657019400389802533367152739617143958437588424926490296825654251606745983923319884191323127808;
data[287]<=640'd719250854131913053886533600199416268714319876565152320826934581244418971175136705353284923978748607418765714524864879523022638784043033728065350926336;
data[288]<=640'd719250854131913053886533600194251889020189375801085952634502467580787897778587313559073042886923527099541983655010247481219456477659807879975913127936;
data[289]<=640'd719250854131913053886533600194252012151449932723157614763438888422482528852273688480803646967833056540942216727422677623965936110000834276624223436800;
data[290]<=640'd719250854131913053886533600235568283544902822198952872709636289402700694008991060984396734001099412085245797927634880120108701026062212591342508310528;
data[291]<=640'd719250854131913053886533600225239838121914563963303497843986300450235660538986888854152814178781732643120579845283400504437378931230003581286443122688;
data[292]<=640'd719250854131913053886533600225239685440343006450389306261352375936971080379037152171098994255458531728619484356755563241843810414731776606912752123904;
data[293]<=640'd719250854131913053886533600225240975240389590977615121549653048079914421652003599515317507121320872338153132705683217662887280359024020418281710026752;
data[294]<=640'd719250854131913053886533600307875765187372507214693956176319500619664494888218699629810017186619892510112047691374381775768206191730453817077568372736;
data[295]<=640'd719250854131913053886533600287222794843719227614129933725756195027948668356501004057910021457950498649542718527763886464404242147188827896323661365248;
data[296]<=640'd719250854131913053886533600287222499328672166373140834038649987502668998387468756010677960698866226339715415955221961672172348931221067783359132860416;
data[297]<=640'd716054195810719752513443498558272486806201980287395889563734169743938988323341750211228189541787287895625183229269806637466046417796349828133076074496;
data[298]<=640'd716054195810719752513443498723536479927252173067244483859558766269051291626509507707747657120232923303169422018570654865081928527056940318848807075840;
data[299]<=640'd716054195810719752513443498723536481158874883499457587595962191555952092861975347895139843247036184052869221329693412692250148544623692447520611368960;
data[300]<=640'd716054195810719752513443498682221130472412500164015030748316599426718847179850664840786266601969270520428233878680726559662575733659658746413042368512;
data[301]<=640'd716054195810719752513443498682219217626935783688236265452195436977737437282247049624759838328005796649578242945000593351105964490429237779900150054912;
data[302]<=640'd818347651926401364867860531027860544143832906622819285070802166648325145936293367879823861257253301713640055421807465536124401416969883210374893797376;
data[303]<=640'd818347651926401364867860531027859302980412246347505941203204878388585547550201790102400479621947948184075711318110122128264813958505529454328717246464;
data[304]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[305]<=640'd0;
data[306]<=640'd0;
data[307]<=640'd0;
data[308]<=640'd0;
data[309]<=640'd0;
data[310]<=640'd0;
data[311]<=640'd0;
data[312]<=640'd0;
data[313]<=640'd0;
data[314]<=640'd0;
data[315]<=640'd0;
data[316]<=640'd0;
data[317]<=640'd0;
data[318]<=640'd0;
data[319]<=640'd0;
data[320]<=640'd0;
data[321]<=640'd0;
data[322]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[323]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[324]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[325]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[326]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[327]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[328]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[329]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[330]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[331]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[332]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[333]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[334]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[335]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[336]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[337]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[338]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[339]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[340]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[341]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[342]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[343]<=640'd398353494612575324017191154914352288844846764696638810260114131509605650307885529420329033517687589677374404780947210779386712874022118574019139283960076830011772872351155913515597824;
data[344]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[345]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[346]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[347]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[348]<=640'd398353494612575324017191154914352186551390649015026455843081537971012733523942897776476074197443525535126815153878457074366752531570804226482521018768785698054402230421841660119875584;
data[349]<=640'd265568996408383549344794103276235029718992369583268475043220513910041109088511359234064155610167347940571714494382458401709398254602728763359583467446130040472067320563817398958817280;
data[350]<=640'd265568996408383549344794103276235029718992369583268475043220542153399150664074058595680099393109723421728823564014629987046110417936094572560149729192181541979598650754760850884526080;
data[351]<=640'd265568996903044352291003171397240071758286749653531173245644265870947140976898850940200584448743909205504922481436351689200150496414012795173930077975219068851482267557512510571544576;
data[352]<=640'd265568996903044352291003171397240071758286749653531173245644265558252819896327359178219133617954960188615259508155358968348673864571206520720809202410771322490992271206384922743799808;
data[353]<=640'd398353495107236126963400223035357228590685029085289154045505297848885066685838825189461651410739422896187426297242838665317545949164137665328712269515090178962203775974916756376387584;
data[354]<=640'd265568996903044352291003171397240071758286749653531173245644338184030641034303117242229689877502164522971427564103021196670092171290393849036582324453145440167845741598409794485485568;
data[355]<=640'd265568996903044352291003171397240071758286749653531173245644327855031128611515395969790338572991288106889471371187128308966430146066594692641115002204262128778152049673123406473592832;
data[356]<=640'd265568996903044352291003171397240071758286749653531173245644307197032103916246678722436962548896293469243128737399025663691577820885618557911557965041435887675500562447747624493645824;
data[357]<=640'd265568997892365958183421307639250155836875509794056569650491832117276525850132101038814803999664947352685383330305512689261723771658093458695782166283893464620766319316229012867514368;
data[358]<=640'd265568996903044352291003171397240071758286749653531173245644472461063818920267927613494590438064006976687019289681191333776707214442910372948086204241920481272126874592137966946091008;
data[359]<=640'd265568996903044352291003171397240071758286749653531173245644431205607106415498351048945982500342200140279227042640518206448955333946888070244009063416593263508288873275499490247180288;
data[360]<=640'd265568996903044352291003171397240071758286749653531173245644431770484387098227638060986536861113849285553400473186921434630770436779591819154968957088195460873412620290859285490958336;
data[361]<=640'd265568996903044352291003171397240071758286749653531173245644766756845724655747473510255706594824695543368075391008313367673797349528654530894869267351649187414430494941395726620426240;
data[362]<=640'd265568996903044352291003171397240071758286749653531173245644843659480909080866790552231080676368793600226952876822552707429198519299934820975122398871077385613727999725727203415031808;
data[363]<=640'd398353495107236126963400223035357228590685029085289154045505876272876844122221199281299545126859726022122334059205504615661116760422648465263434564713455934430047793314326588816359424;
data[364]<=640'd265568996903044352291003171397240071758286749653531173245645484702994982139725872965258139836562807659282043279684631898945903919829267023699733195241668281122035439496027543105961984;
data[365]<=640'd265568996903044352291003171397240071758286749653531173245645340097000579162458233375088372050565688726667460553454196218566568069607323140557732441880137923280415860907149770532847616;
data[366]<=640'd265568996903044352291003171397240071758286749653531173245645174833028082302793242040816850208002287043364119848697241519436780164328392567484269535213354364233174627674152840600748032;
data[367]<=640'd265568997892365958183421307639250155836875509794056569650493856601337324502862867062672605271651108427048876329190094906304104597697945171522775673170267909795562382300825067007770624;
data[368]<=640'd398353495107236126963400223035357228590685029085289154045507531495314049022707758805221808527669066460065147963112017655568023638169995171863509723114198942463964854009681611778424832;
data[369]<=640'd265568996903044352291003171397240071758286749653531173245646166982367429213654653607639590747946535849447754254214342759981391193928366993523644887359573947682335248412627898218840064;
data[370]<=640'd265568996903044352291003171397240071758286749653531173245646168838908693948757269410713320960433747478933289273331719673164322356616834544702525663131062790607969032125819749335564288;
data[371]<=640'd265568996903044352291003171397240071758286749653531173245648820651452948170946773728445373595175963805733747734958428812846622296264991660556917029629575456997943970807968902695354368;
data[372]<=640'd265568997892365958183421307639250155836875509794056569650496830070743775665005331346202969610616535024674669991064294781277940123279233337905270013843241342490693245972345363328139264;
data[373]<=640'd265568996903044352291003171397240174051742865335143527662682054913947799261606721964401616714338507026402603841286661204148291631905629204376219183101830592291163931199020767880675328;
data[374]<=640'd265568996903044352291003171397240174051742865335143527662679255747514454022224283900141070411542534696719932584147492194075207522237814138723162892139430987789628858278988575806586880;
data[375]<=640'd265568996903044352291003171397240174051742865335143527662676776787630872528466918948602142292013070382638162388580928377582346718311671832780261709203522302229601390475521153055064064;
data[376]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[377]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[378]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[379]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[380]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[381]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[382]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[383]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[384]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[385]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[386]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[387]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[388]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[389]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[390]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[391]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[392]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[393]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[394]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[395]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[396]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[397]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[398]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[399]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[400]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[401]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[402]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[403]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[404]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[405]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083711154225492614732989228270490262743671417864192;
data[406]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083756826325883777643510875830043263955216103374848;
data[407]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083733993150393632101736882977413894943200384122880;
data[408]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260510356823990064450203354978959320258094768848896;
data[409]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841306678842167437339742438259765413224120320;
data[410]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841295784489368253867537777416344549361451008;
data[411]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083866058175805198939743815208226653779662768963584;
data[412]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934544014703162186716804046514368768030868556417597440;
data[413]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260686614913495185286957388911191037195542417375232;
data[414]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083871185952298368884399164504508543769418921934848;
data[415]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986330444476161582688175652864;
data[416]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[417]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[418]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[419]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[420]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[421]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[422]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[423]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[424]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[425]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[426]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[427]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[428]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[429]<=640'd398353496343888134328922893337869117634725168541193386108065983048744062545919757800094946891136771680368312041868575743622909878699085669704398453847763599671125628542792319314690048;
data[430]<=640'd531137992816767098689588206552468627329593117540961209779768774219776665041523081944630313929275862236827838496002843258316710966147798256686047195211381820739689719850535202106376192;
data[431]<=640'd464745747548292448942947204772883260336491728765709340960903687623617040888630979714838395224460056055998811059991606943419003558340812870361086397939032316978126257926111479799480320;
data[432]<=640'd1731312810311731738423517647137530330245919443708482879398441392650280575745723070192214807428701314927183699982112975375459555240147258469772823085713252175416247405040893952;
data[433]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[434]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[435]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[436]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[437]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[438]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[439]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[440]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[441]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[442]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[443]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[444]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[445]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[446]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[447]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[448]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[449]<=640'd741991204419313602181507563058941570105394047303635519742189168278691675319595601510949203183729134968793014278048418018054095102920253629902638465305679503749820316446097408;
data[450]<=640'd989321605892418136242010084078576565810250724560193525292073344815707069964632683637707560663098643350035920994610962411690368371714661765920491625786887328011429868730318848;
data[451]<=640'd1799565517869652802850553672994603778697120433756232925976991265676467694158133288870091067319688664337182830767822544995324267558345195980337572361199321983483904;
data[452]<=640'd0;
data[453]<=640'd0;
data[454]<=640'd0;
data[455]<=640'd0;
data[456]<=640'd0;
data[457]<=640'd0;
data[458]<=640'd0;
data[459]<=640'd0;
data[460]<=640'd0;
data[461]<=640'd0;
data[462]<=640'd0;
data[463]<=640'd0;
data[464]<=640'd0;
data[465]<=640'd0;
data[466]<=640'd0;
data[467]<=640'd0;
data[468]<=640'd0;
data[469]<=640'd0;
data[470]<=640'd0;
data[471]<=640'd0;
data[472]<=640'd0;
data[473]<=640'd0;
data[474]<=640'd0;
data[475]<=640'd0;
data[476]<=640'd0;
data[477]<=640'd0;
data[478]<=640'd0;
data[479]<=640'd0;
end
else if(choise == 3) begin
data[0]<=640'd0;
data[1]<=640'd0;
data[2]<=640'd0;
data[3]<=640'd0;
data[4]<=640'd0;
data[5]<=640'd0;
data[6]<=640'd0;
data[7]<=640'd0;
data[8]<=640'd0;
data[9]<=640'd0;
data[10]<=640'd0;
data[11]<=640'd0;
data[12]<=640'd0;
data[13]<=640'd0;
data[14]<=640'd0;
data[15]<=640'd0;
data[16]<=640'd0;
data[17]<=640'd0;
data[18]<=640'd0;
data[19]<=640'd0;
data[20]<=640'd0;
data[21]<=640'd0;
data[22]<=640'd0;
data[23]<=640'd0;
data[24]<=640'd0;
data[25]<=640'd0;
data[26]<=640'd0;
data[27]<=640'd0;
data[28]<=640'd0;
data[29]<=640'd0;
data[30]<=640'd0;
data[31]<=640'd85070591732710495944414412407740301312;
data[32]<=640'd730750818665451459101842416358132502628711530496;
data[33]<=640'd27021597764222976;
data[34]<=640'd9007199254740992;
data[35]<=640'd9007199254740992;
data[36]<=640'd9007199254740992;
data[37]<=640'd9007199254740992;
data[38]<=640'd9007199254740992;
data[39]<=640'd9007199254740992;
data[40]<=640'd13510798882111488;
data[41]<=640'd9007199254740992;
data[42]<=640'd9007199254740992;
data[43]<=640'd9007199254740992;
data[44]<=640'd9007199254740992;
data[45]<=640'd13510798882111488;
data[46]<=640'd9007199254740992;
data[47]<=640'd9007199254740992;
data[48]<=640'd9007199254740992;
data[49]<=640'd13510798882111488;
data[50]<=640'd31525197391593472;
data[51]<=640'd309787241346054520360140800;
data[52]<=640'd599375721660670508425266668362373856774380817170532873411752110287376594018075499955962254745047801101257078721539110295345450208080468874490806272;
data[53]<=640'd5027929472167778066878457916438579271401010308215785621888644634346722099039006813346457612736872842782101791232293722601083851606530876499670384477470720;
data[54]<=640'd26396628205467732864788082285642163171681467387598851022504789516166031859271295734080499794632056350026575515206137239670386077067062433013666803051659264;
data[55]<=640'd107052979177370224261959331447169757995624348293019147030047829383530188356005728063506518606159218349527795023329677542352008354006734679382389176714395648;
data[56]<=640'd214315455403593848371243628535063509913572769065503325629120859826805569962864356697324533626196254014778770029289013968377661500181271326886728884677509120;
data[57]<=640'd428840407856041074259963789741753073154462173194139026648524031365156604373179187965892171529647976321944478726877311152888398901532830347995215140384407552;
data[58]<=640'd857890312710984452973429432205287855794666022103459363145609269421919230326598971951740951076827667545097005016360117896252295914307608837212705991216332800;
data[59]<=640'd1715990122520767163402835295025441171969567992656791332698788381890886667082526282063613182540215233834685701369746996036155842454675129901135972923267350528;
data[60]<=640'd3381910457608045116620999402357853392069290396874125430328045293723256668427299865470942285888501138062814744645993448611444427055806175678689141383990607872;
data[61]<=640'd6760678458734064500004395559042319423859994262652645444346415197021551412634851879054371547607344496682524987027586199293328324311640523138232093438226989056;
data[62]<=640'd13518213642638457425626434681613824247268059382700472661371176154298941598148001792901619029354125148973649014067957618735459638875554094018914426032008200192;
data[63]<=640'd13303689508433767673001792403097267332445570694662408114543717372905665493958789517438273337383157632243321737455198609118372135649314003991232408626193760256;
data[64]<=640'd26604027063486494151856852108440019966858802187707887285518607084327113815165657061281383825521489522527025728247401310676293068991128914079610415427673391104;
data[65]<=640'd54066572828686917512538848091696728615772215835780101081038941672982135750213955630549554187526714626306345586352280791600468548118337364405108883342695071744;
data[66]<=640'd108126854402215468636948495822802328610646555176645496568601164575687211790167285726112387578570729443792281568925608496419361685686955605409517285680324018176;
data[67]<=640'd106410661329377119006977893772893853047864231581297737945232268808300772200366709756376036593409518210486072502430351275254099497567078879082869518791243464704;
data[68]<=640'd216247436575855479282092410736678649095590945920787579121648876487916844005673158738319991589732162304852207301197122119583818767818967446770323958965500641280;
data[69]<=640'd212814617933244944225846956985053715385389454010758270613221946629202400863949106570233714202028220831395569769179299962980594675440578057599903261196493520896;
data[70]<=640'd425630075491580350373514556489764094002022545108418790299028410609512909024529356069086987000409094756423964141442302784669197120254938147435314767835038744576;
data[71]<=640'd864977176477493792998426720553126075865707973051461377546367259004900087853513061839282910684749462706454618560081417516813094727567860441403240096422265094144;
data[72]<=640'd851247682632341467128970141392075156053575187939118035919251798845312188512943540402250903746277609282808142921882505770245391633396799966707883547220447854592;
data[73]<=640'd1729955184390208237472303383221228712183658530661859015675224928698743183157140205290275958981656649640543026924220237830657450719240773284034815281766284132352;
data[74]<=640'd1702495365258689079671238639778692186686648698691038037051379820481306262388471864585215024917390711291478313796939795069715334066961525319969474466567994474496;
data[75]<=640'd3459883972158554305902524366150836688105814640052773469618604938651459850491363095953710892695995849384108774563596257108611723471560113782663469689111389929472;
data[76]<=640'd3404966402678380287026472699061892275557714108338375202607199483365135647893772515601448216130947937129818071330403331790953794098718246683046836199909150949376;
data[77]<=640'd6919769620281112346282473663417035300574804215453964264447298784452164613972549122915290026490312135640287871664655176173607558561847291296195597047089902649344;
data[78]<=640'd6809932805344772864421133650764320560533861927265129952552077886232105511571101450500741662581779928543593774435373931650172041152181291712486836710752275922944;
data[79]<=640'd13839485504582804636771634314557442765540704517288645763211024595086836483792384167084161877332950073509926851413873715336011710023323021165928452172413373775872;
data[80]<=640'd13619811979458625123224703741313646734349949348047649061338701020815318781929897902843165232488609907086914327981229207162956470717094728387741441325879816880128;
data[81]<=640'd27678971009140035495573996324079679547060880019621936630943123616759766761141886885221954464300421961469106309459060756254840548257620172840974207485516475006976;
data[82]<=640'd27239623539897679053327564100571767080268538237049088531596804344288460452819900738111875815959250704898749886308357836242488687851363195978447168975123953745920;
data[83]<=640'd55357834755792656445893429784966008765323002970073268929816810071248050828911928509004133547621889284623934433607299484814503444967508689819300071169627483275264;
data[84]<=640'd54479247079796955661475752410167943692920068694349925510592349617495011916437736470975248442430863494517913342821690832962759812414814875610540376595600097935360;
data[85]<=640'd110715669511586911227044760910989549664951290921252942767736421845620006903796688988886746286888562537833446547416159306317038729986015682962372443556378803437568;
data[86]<=640'd108958279634617483897186059353955721834531173292492643743446586046970229497852579626815538309591923960744126037655557682374053725383735175296355788649654040657920;
data[87]<=640'd108958276282663903076283488369549075760180252722079693234698334086877633526618490491310064159152584231270217074212862956664341061242741187353202903905637178015744;
data[88]<=640'd221431335671170693240215314621644771431426395490521791277898172646833623334842425363648422135228700058062154206682413788871748700324389950795583538713360416636928;
data[89]<=640'd217916552565331002823165766959398391001306435154144838499707258298812106106143536212746440113533544594240287378617390005937186876393157600823930063484681833152512;
data[90]<=640'd442862242292490821964359011659308181960156777221913368692767379022222992390025038628709715690211444402007032171733189041754440386983041800259773752932296824979456;
data[91]<=640'd442862228884679695448036652215884974418818052233948439596294440625308896041677152899905542243931370874668803798369585865243004234553139213729170333811226439581696;
data[92]<=640'd435833105130508562534745063552623256078125856084596639737079105219936424717994818075581101639306710098286409836474796876868486384501888739015930737911622812041216;
data[93]<=640'd435833078314886309308436457572871538053355971474607200970256890968555190777274628892512546854519477174740741143016318386965325376872929856817777546809377032241152;
data[94]<=640'd421773972706900460565300364381239083639546980409929178366340363577876513135139219757465394741596352353179657050576974825036112800830974047350341605563815455358976;
data[95]<=640'd421773490025814980266866852072168080722746520326731594415381246511774577959324591550086354122775601042723754080244766925928918731942453508047105353713736589770752;
data[96]<=640'd168709267295369864355395194106365450110326787925898158555921256322683905591083810756201579645300549095178113289751200261547810419468161304768314266015640158470144;
data[97]<=640'd9007199271518208;
data[98]<=640'd9007199271518208;
data[99]<=640'd9007199305072640;
data[100]<=640'd13510798898888704;
data[101]<=640'd9007199271518208;
data[102]<=640'd9007199271518208;
data[103]<=640'd9007199271518208;
data[104]<=640'd9007199305072640;
data[105]<=640'd13510798898888704;
data[106]<=640'd9007199271518208;
data[107]<=640'd9007199271518208;
data[108]<=640'd9007199271518208;
data[109]<=640'd9007199271518208;
data[110]<=640'd13510798898888704;
data[111]<=640'd9007199271518208;
data[112]<=640'd9007199271518208;
data[113]<=640'd9007199271518208;
data[114]<=640'd9007199305072640;
data[115]<=640'd13510798898888704;
data[116]<=640'd9007199271518208;
data[117]<=640'd9007199271518208;
data[118]<=640'd9007199271518208;
data[119]<=640'd9007199305072640;
data[120]<=640'd9007199271518208;
data[121]<=640'd9007199271518208;
data[122]<=640'd9007199271518208;
data[123]<=640'd9007199271518208;
data[124]<=640'd9007199271518208;
data[125]<=640'd13510798898888704;
data[126]<=640'd9007199271518208;
data[127]<=640'd9007199271518208;
data[128]<=640'd9007199271518208;
data[129]<=640'd533996758980227548388856843498274930307712532674261077271556721709290300914980308412090940391424;
data[130]<=640'd1868988656430796558311506037023396764362175874785403194374430124751192900551531866420075563057152;
data[131]<=640'd70608395103938906748405908848113786735498346477469127413701232021435384158860502965062554256599959879843061883878768640;
data[132]<=640'd320259506364294327037405639924244233692028483547307954462621785835688912818792645285933467907937828686853293558248505344;
data[133]<=640'd1636695303852802729735721062057007209171471377742890289643062904937418624395482718595003351178232432600793374821907689755208590573672079544628279246848;
data[134]<=640'd1636695303852802729735721062058147030406720677237543099851066895318485373478903061535747386712734283593220464541437540325981490295668695865160609300480;
data[135]<=640'd1636695303852802729735721062065404564732046969152611200271195788852249740197418431205925877357108034363812204308885191990930668944454828233263325118464;
data[136]<=640'd1432108391621439505026886996886717169273864967559035645802998680124266543704676409646449470163531041179254364961423359278795446832131342830488728371200;
data[137]<=640'd1432108391621439505026886996904792918420473327686627080007019763244601044180741872875958218823407205924272963993675377937932973822672338671949406273536;
data[138]<=640'd1432108391621439505026886996940944416713690047941809952687036001327029501520034157640508399872311787975085208710858581108289465131830540530627962208256;
data[139]<=640'd1432108391621439505026886997013247413300123488452175689503120333808321972122134470033220033847614419284429732306322481390539143083906703564612258758656;
data[140]<=640'd1432108391621439505026886996992589414275428219734928335071630492107686374016258216053810355123933847131021312988412579121760328376010588614750415880192;
data[141]<=640'd1432108391621439505026886997116552548875351926674048803359290596818587304240900274827643548059306807017147154621225407180839476298628368035496429879296;
data[142]<=640'd1432108391621439505026886997447224277695550190362521311331009167475215864237658663636716821857020275584059608091812043003909209505308931123163491729408;
data[143]<=640'd1432108391621439505026886997365723278023620873331869727152474194724948003708818863349359636397631083540867698410506682259627063857046814088751761850368;
data[144]<=640'd1432108391621439505026886997865358389702177150605165303145258429402837446582954197638295636923873398044756134233409858196019054312570197228487975108608;
data[145]<=640'd1432108391621439505026886997865074693978380074121854890236161915340260594625376070520270905906096337945375461411509381279946242164821610597170840338432;
data[146]<=640'd1432108391621439505026886998854409262952676980504621109721009824267732975110142491754913744821047592131340536058964915344021645435596313560973708361728;
data[147]<=640'd1432108391621439505026886998851827008149193100032196504936387199730249542554028750995786366208166543904089351905520081125512928689697626404479748276224;
data[148]<=640'd1432108391621439505026886998851844660249461589263663137068926051993840052404754591566545789242465351085204514756844446676376195612999575383996222144512;
data[149]<=640'd1432108391621439505026886998851880003851417626235672409156543054723011927644083903878583113956520208122970877229942782243849384203947466329057474379776;
data[150]<=640'd1432108391621439505026886998851960689309465379937974215348640987936299799157058308259933202125717275149084196427410320986260374569061910111429653954560;
data[151]<=640'd1432108391621439505026886999182639977407932912318160474930286812633850667917497385985339999057114568437894464897525317349637161329206581616471477059584;
data[152]<=640'd1432108391621439505026886999182942584814920873430650423032694709628170154583606385661603819914208139368650191170835502616397517265060376598406542393344;
data[153]<=640'd1432108391621439505026886998027910362682132534108847785449568960627476270656738845839804216555704037225247595403564818688043503454028482857191008632832;
data[154]<=640'd1432108391621439505026886997529374725893571591274898906303286495872453939078611570843770547722574507543904434341396434297579741388017383966642400133120;
data[155]<=640'd1432108391621439505026886997197878397791758610023294126888758972915747772504473914776023068001049077871092589863193076052654946685102377569148978855936;
data[156]<=640'd1432108391621439505026886996940944456116278685118659163126484435799439642037184193056598196011954859360205143397155628336586548693470503394095768010752;
data[157]<=640'd1432108391621439505026886996868641420127256607431444208395909635239964769402726650831033115052207720387956190202354378611678955879848565437861870960640;
data[158]<=640'd1432108391621439505026886996868641420127256607431444208396822227357362619169374914499440516468358778228318529642639369532989718702142540282232032985088;
data[159]<=640'd1432108391621439505026886996868641420127256607431444208398647411592158318702671441836255319300660893909043208523209351375611244346730489970972357033984;
data[160]<=640'd1432108391621439505026886996868641420127256607431444208402297780061749717769264496509884924965265125270492566284349315060854295635906389348453005131776;
data[161]<=640'd1432108391621439505026886996868641420127256607431444208426285915719064625921161712936593762189807217074302631571840504992451489821919442400468675854336;
data[162]<=640'd1432108391621439505026886996868641420127256607431444208657823572933147652430778323663957321487561320571947609564146773027867885878219345772098355200000;
data[163]<=640'd1432108391621439505026886996868641420127256607431444208645308023894548569916744993354370102066061098761264097240238326107034567172473405049307561721856;
data[164]<=640'd1636695303852802729735721062055718605960824492694731914513886315868436735039865809623431264300745114147225121181134921005965207090773500786651179253760;
data[165]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[166]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
data[167]<=640'd0;
data[168]<=640'd0;
data[169]<=640'd0;
data[170]<=640'd0;
data[171]<=640'd0;
data[172]<=640'd0;
data[173]<=640'd0;
data[174]<=640'd0;
data[175]<=640'd0;
data[176]<=640'd0;
data[177]<=640'd0;
data[178]<=640'd0;
data[179]<=640'd0;
data[180]<=640'd0;
data[181]<=640'd0;
data[182]<=640'd0;
data[183]<=640'd0;
data[184]<=640'd0;
data[185]<=640'd0;
data[186]<=640'd0;
data[187]<=640'd0;
data[188]<=640'd0;
data[189]<=640'd0;
data[190]<=640'd0;
data[191]<=640'd0;
data[192]<=640'd0;
data[193]<=640'd0;
data[194]<=640'd0;
data[195]<=640'd0;
data[196]<=640'd0;
data[197]<=640'd0;
data[198]<=640'd0;
data[199]<=640'd0;
data[200]<=640'd0;
data[201]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[202]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[203]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
data[204]<=640'd716054195810719752513443498452396459210236663843313538401519604681591400367843758171127472313812864627914813743442211318145061348828617500555078533120;
data[205]<=640'd716054195810719752513443498454817318470943140646115962625272428313775499548621155214406215460569721773555602363407503836845190565799776724279529308160;
data[206]<=640'd716054195810719752513443498516942619248823106185030406280912270583849488969373445934094087849421263174083520826805540203121430985236360613379530817536;
data[207]<=640'd716054195810719752513443498599582180532793891087527193434379346215841788567102110100978117211933049057178062906913029171650412120303285071331498917888;
data[208]<=640'd716054195810719752513443498594424617992336026611211666968870954002199316658579354529295692867369532881627382597869581719349971971229802136622671593472;
data[209]<=640'd716054195810719752513443498470474108272331322421689801733046036933826550285750168652928145848503239957568531354763767237227511749508443218334678253568;
data[210]<=640'd716054195810719752513443498465308672718510340873496671745117643480671118166195844841114120965026022274926009181593149300629143946687042173319644184576;
data[211]<=640'd716054195810719752513443498506624657223461246003890533286174287434856891565124599078778989884953122375513294241757993247051690560743735994951435026432;
data[212]<=640'd716054195810719752513443498506624652298210471454580631885054205267145339708975597071443380104758889826892124014399521046811419350104215025143861215232;
data[213]<=640'd716054195810719752513443498496295652785862855443945883084174268069311714182345803205975936425142028849943491336863722245241643132224477161940351713280;
data[214]<=640'd716054195810719752513443498578928594532792639193439159305090028273801748502798542518557450139198694610470892581121084791661332217742187629441106051072;
data[215]<=640'd716054195810719752513443498578935529295615565084795285312521661142683621566827201523159863495089171062366134461495250180271803632698486581077173338112;
data[216]<=640'd716054195810719752513443498558306559719295686255939994691463852412789730990382003880051374333913264620660854005355689082322410824234160602443344248832;
data[217]<=640'd716054195810719752513443498723684029695915337013595158856156430908443933135962537296006781336619137107590586039828334070534992578101058502990789345280;
data[218]<=640'd716054195810719752513443498726074667662435116152319054365729584236292666552544995954241525497930953128181220600548079562723803871197520873352868134912;
data[219]<=640'd716054195810719752513443498764687372869500969648166995387713925429748206448310492740292313345780339563283646892842795758416380402056113891813774852096;
data[220]<=640'd716054195810719752513443498762266503828035350362723319525822871017568885791056302026571382589134451089783145982566227641658649420802696355669019197440;
data[221]<=640'd716054195810719752513443499012744741992836455529709340851102690530689620425974536127085317615947573415639164249983869881973447411020431322848130236416;
data[222]<=640'd716054195810719752513443498930112824678828498850708675602916998574373097638935264627451193163361309192489206596011604979186284746446998068957171154944;
data[223]<=640'd716054195810719752513443498930112805131814622444746571190038572981539243817399858943490253968280715111299464596629928971483814150922352367596472369152;
data[224]<=640'd716054195810719752513443499591168773883566058145757224900889316156738702612168354968539617553353773703844976370883228066977480014210530902843334852608;
data[225]<=640'd716054195810719752513443499591168931491741113896338500626710837487951928012927739405129935394457478811456723544995424280807755658899542164501228945408;
data[226]<=640'd716054195810719752513443499425904939601969561137220759507440701221919135022913033671278759931037052797222372081332600693355028792468667943584333299712;
data[227]<=640'd716054195810719752513443499425904900123006321892684327391627979833966398203541687810086025966492434445610482967791808411731173206438044431614669225984;
data[228]<=640'd716054195810719752513443500748016837703804356719440658621889048670187383705742252154792706093711491586733855110068319510099229844196759380564610383872;
data[229]<=640'd716054195810719752513443500748017152919778787986916839628238819076166832342626120149144509311646161009324757501601892866314905534279262675934774296576;
data[230]<=640'd716054195810719752513443500417489168524654615226286366532113576586219958341702119533547297296133204822806923134614207553653809644564894950407257718784;
data[231]<=640'd716054195810719752513443499756432805560279541931114698735649863252824271402368568143057938395255371826363848621175488615897430102674974581120177274880;
data[232]<=640'd818347651926401364867860531027859302980412393131277380521395508717963006741230473315177183548362701793830182762363954799343770380606623659043181297664;
data[233]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[234]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[235]<=640'd0;
data[236]<=640'd0;
data[237]<=640'd0;
data[238]<=640'd0;
data[239]<=640'd0;
data[240]<=640'd0;
data[241]<=640'd0;
data[242]<=640'd0;
data[243]<=640'd0;
data[244]<=640'd0;
data[245]<=640'd0;
data[246]<=640'd0;
data[247]<=640'd0;
data[248]<=640'd0;
data[249]<=640'd0;
data[250]<=640'd0;
data[251]<=640'd0;
data[252]<=640'd0;
data[253]<=640'd0;
data[254]<=640'd0;
data[255]<=640'd0;
data[256]<=640'd0;
data[257]<=640'd0;
data[258]<=640'd0;
data[259]<=640'd0;
data[260]<=640'd0;
data[261]<=640'd0;
data[262]<=640'd0;
data[263]<=640'd0;
data[264]<=640'd0;
data[265]<=640'd0;
data[266]<=640'd0;
data[267]<=640'd0;
data[268]<=640'd0;
data[269]<=640'd0;
data[270]<=640'd0;
data[271]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[272]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[273]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[274]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[275]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
data[276]<=640'd716054195810719752513443498436902329509616069993710626904859931137792284335040089646996829001874510964265422620294556570204156201562945562670748663808;
data[277]<=640'd716054195810719752513443498475636077680919698838549414484905109252737871227478442339456719349984225294518040539739236869406223673101493142261961064448;
data[278]<=640'd716054195810719752513443498764203131989230876044265778420883288506903374851972497345429589616096064986448387994971887726721704494713925516264338358272;
data[279]<=640'd716054195810719752513443501075962335346535790933735072534116409542307789640129758881856114652118974840552957684284325086262295903437522520986112491520;
data[280]<=640'd716054195810719752513443508936330964243310997934299320101161945139223999366914197463078394669438236193084646203335782881574369898171715801520548085760;
data[281]<=640'd716054195810719752513443519265330476590982933239308044822392414689331103834041171381277090042968167159521430263441464572718312641489842287878613237760;
data[282]<=640'd716054195810719752513443518284075522917920092488719067374528189671023665650908402235286529253574501650522280565529526920176121880409916046746893418496;
data[283]<=640'd716054195810719752513443498452396459210462123931259826391396994818883176722471823695822671021400764561181905809853213728717576452673555296046144290816;
data[284]<=640'd716054195810719752513443498449814209332375215341603907219393982944553470929642600182992011664860116939165064615223568375437438621237652124073396797440;
data[285]<=640'd716054195810719752513443498449814209332675828792198959741552492891738828164790680447610376885677107245592361074099645100643052151091383788153310543872;
data[286]<=640'd716054195810719752513443498470472208357296532456069495355220800717315295409424067509323404103846287738224339862431283562756427942171383677257546465280;
data[287]<=640'd716054195810719752513443498470472245296789193897524885153498362561344464051193620122991184124157306732063564090470508834172320742291097521131574263808;
data[288]<=640'd716054195810719752513443498465307865602658693133458516961066248897713390654644228328779303032332226412839833220615876792369138435907871673042136465408;
data[289]<=640'd716054195810719752513443498465307988733919250055530179090002669739408021728330603250509907113241755854240066293028306935115618068248898069690446774272;
data[290]<=640'd716054195810719752513443498506624260127372139531325437036200070719626186885047975754102994146508111398543647493240509431258382984310276384408731648000;
data[291]<=640'd716054195810719752513443498496295814704383881295676062170550081767161153415043803623859074324190431956418429410889029815587060889478067374352666460160;
data[292]<=640'd716054195810719752513443498496295662022812323782761870587916157253896573255094066940805254400867231041917333922361192552993492372979840399978975461376;
data[293]<=640'd716054195810719752513443498496296951822858908309987685876216829396839914528060514285023767266729571651450982271288846974036962317272084211347933364224;
data[294]<=640'd716054195810719752513443498578931741769841824547066520502883281936589987764275614399516277332028591823409897256980011086917888149978517610143791710208;
data[295]<=640'd716054195810719752513443498558278771426188544946502498052319976344874161232557918827616281603359197962840568093369515775553924105436891689389884702720;
data[296]<=640'd716054195810719752513443498558278475911141483705513398365213768819594491263525670780384220844274925653013265520827590983322030889469131576425356197888;
data[297]<=640'd716054195810719752513443498558272486806201980287395889563734169743938988323341750211228189541787287895625183229269806637466046417796349828133076074496;
data[298]<=640'd716054195810719752513443498723536479927252173067244483859558766269051291626509507707747657120232923303169422018570654865081928527056940318848807075840;
data[299]<=640'd716054195810719752513443498723536481158874883499457587595962191555952092861975347895139843247036184052869221329693412692250148544623692447520611368960;
data[300]<=640'd716054195810719752513443498682221130472412500164015030748316599426718847179850664840786266601969270520428233878680726559662575733659658746413042368512;
data[301]<=640'd716054195810719752513443498682219217626935783688236265452195436977737437282247049624759838328005796649578242945000593351105964490429237779900150054912;
data[302]<=640'd818347651926401364867860531027860544143832906622819285070802166648325145936293367879823861257253301713640055421807465536124401416969883210374893797376;
data[303]<=640'd818347651926401364867860531027859302980412246347505941203204878388585547550201790102400479621947948184075711318110122128264813958505529454328717246464;
data[304]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
data[305]<=640'd0;
data[306]<=640'd0;
data[307]<=640'd0;
data[308]<=640'd0;
data[309]<=640'd0;
data[310]<=640'd0;
data[311]<=640'd0;
data[312]<=640'd0;
data[313]<=640'd0;
data[314]<=640'd0;
data[315]<=640'd0;
data[316]<=640'd0;
data[317]<=640'd0;
data[318]<=640'd0;
data[319]<=640'd0;
data[320]<=640'd0;
data[321]<=640'd0;
data[322]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[323]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[324]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[325]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[326]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[327]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[328]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[329]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[330]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[331]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[332]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[333]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[334]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[335]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[336]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[337]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[338]<=640'd398353494612575324017191154914351470497194838295273942399583103650302669895639182054371876698921964251666997114684875761509934503239530429557139984074940513957873453126544914273796096;
data[339]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[340]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[341]<=640'd265568996408383549344794103276234313664796558863515961599722069100201779930426121369581251132614642834444664743123250507673289668826353619704759989383293675971915635417696609515864064;
data[342]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[343]<=640'd398353494612575324017191154914352288844846764696638810260114131509605650307885529420329033517687589677374404780947210779386712874022118574019139283960076830011772872351155913515597824;
data[344]<=640'd265568996408383549344794103276235132012448485264880829460253096959504760342672468735538407951380268260152072409385585525550068039608941764166759289268429992025815054642307608757665792;
data[345]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[346]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[347]<=640'd265568996408383549344794103276235029718992369583268475043220503420911843558729837091685448631136204117904482782316831820530107697157627416630141024077138860068444412712993355361943552;
data[348]<=640'd398353494612575324017191154914352186551390649015026455843081537971012733523942897776476074197443525535126815153878457074366752531570804226482521018768785698054402230421841660119875584;
data[349]<=640'd265568996408383549344794103276235029718992369583268475043220513910041109088511359234064155610167347940571714494382458401709398254602728763359583467446130040472067320563817398958817280;
data[350]<=640'd265568996408383549344794103276235032915650690776569848133322271097422568194756726223115772829328406496235947507099860280785965009236781274710584123562870392297640402690967784661188608;
data[351]<=640'd265568996903044352291003171397240074954945070846832546335745994814970558507581518567636257884962592280012046424521581982940005087714699497324364472345907919169524019493719444348207104;
data[352]<=640'd265568996903044352291003171397240074954945070846832546335745994502276237427010026805654807054173643263122383451240589262088528455871893222871243596781460172809034023142591856520462336;
data[353]<=640'd398353495107236126963400223035357231787343350278590527135607026792908484216521492816897324846958105970694550240328068959057400540464824367479146663885779029280245527911123690153050112;
data[354]<=640'd265568996903044352291003171397240074954945070846832546335746067128054058564985784869665363313720847597478551507188251490409946762591080551187016718823834290485887493534616728262148096;
data[355]<=640'd265568996903044352291003171397240074954945070846832546335746056799054546142198063597226012009209971181396595314272358602706284737367281394791549396574950979096193801609330340250255360;
data[356]<=640'd265568996903044352291003171397240074954945070846832546335746036141055521446929346349872635985114976543750252680484255957431432412186305260061992359412124737993542314383954558270308352;
data[357]<=640'd265568997892365958183421307639250159033533830987357942740593561061299943380814768666250477435883630427192507273390742983001578362958780160846216560654582314938808071252435946644176896;
data[358]<=640'd265568996903044352291003171397240074954945070846832546335746201405087236450950595240930263874282690051194143232766421627516561805743597075098520598612609331590168626528344900722753536;
data[359]<=640'd265568996903044352291003171397240074954945070846832546335746160149630523946181018676381655936560883214786350985725748500188809925247574772394443457787282113826330625211706424023842816;
data[360]<=640'd265568996903044352291003171397240074954945070846832546335746160714507804628910305688422210297332532360060524416272151728370625028080278521305403351458884311191454372227066219267620864;
data[361]<=640'd265568996903044352291003171397240074954945070846832546335746495700869142186430141137691380031043378617875199334093543661413651940829341233045303661722338037732472246877602660397088768;
data[362]<=640'd265568996903044352291003171397240074954945070846832546335746572603504326611549458179666754112587476674734076819907783001169053110600621523125556793241766235931769751661934137191694336;
data[363]<=640'd398353495107236126963400223035357231787343350278590527135607605216900261652903866908735218563078409096629458002290734909400971351723335167413868959084144784748089545250533522593021952;
data[364]<=640'd265568996903044352291003171397240074954945070846832546335747213647018399670408540592693813272781490733789167222769862192685758511129953725850167589612357131440077191432234476882624512;
data[365]<=640'd265568996903044352291003171397240074954945070846832546335747069041023996693140901002524045486784371801174584496539426512306422660908009842708166836250826773598457612843356704309510144;
data[366]<=640'd265568996903044352291003171397240074954945070846832546335746903777051499833475909668252523644220970117871243791782471813176634755629079269634703929584043214551216379610359774377410560;
data[367]<=640'd265568997892365958183421307639250159033533830987357942740595585545360742033545534690108278707869791501556000272275325200043959188998631873673210067540956760113604134237032000784433152;
data[368]<=640'd398353495107236126963400223035357228590685029085289154045507531495314049022707758805221808527669066460065147963112017655568023638169995171863509723114198942463964854009681611778424832;
data[369]<=640'd265568996903044352291003171397240071758286749653531173245646166982367429213654653607639590747946535849447754254214342759981391193928366993523644887359573947682335248412627898218840064;
data[370]<=640'd265568996903044352291003171397240071758286749653531173245646168838908693948757269410713320960433747478933289273331719673164322356616834544702525663131062790607969032125819749335564288;
data[371]<=640'd265568996903044352291003171397240071758286749653531173245648820651452948170946773728445373595175963805733747734958428812846622296264991660556917029629575456997943970807968902695354368;
data[372]<=640'd265568997892365958183421307639250155836875509794056569650496830070743775665005331346202969610616535024674669991064294781277940123279233337905270013843241342490693245972345363328139264;
data[373]<=640'd265568996903044352291003171397240174051742865335143527662682054913947799261606721964401616714338507026402603841286661204148291631905629204376219183101830592291163931199020767880675328;
data[374]<=640'd265568996903044352291003171397240174051742865335143527662679255747514454022224283900141070411542534696719932584147492194075207522237814138723162892139430987789628858278988575806586880;
data[375]<=640'd265568996903044352291003171397240174051742865335143527662676776787630872528466918948602142292013070382638162388580928377582346718311671832780261709203522302229601390475521153055064064;
data[376]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[377]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[378]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[379]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[380]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[381]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[382]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[383]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[384]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[385]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[386]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[387]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[388]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[389]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[390]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[391]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[392]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[393]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[394]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[395]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[396]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[397]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[398]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[399]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[400]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[401]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[402]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[403]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[404]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[405]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083711154225492614732989228270490262743671417864192;
data[406]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083756826325883777643510875830043263955216103374848;
data[407]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083733993150393632101736882977413894943200384122880;
data[408]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260510356823990064450203354978959320258094768848896;
data[409]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841306678842167437339742438259765413224120320;
data[410]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083791841295784489368253867537777416344549361451008;
data[411]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083866058175805198939743815208226653779662768963584;
data[412]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934544014703162186716804046514368768030868556417597440;
data[413]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260686614913495185286957388911191037195542417375232;
data[414]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083871185952298368884399164504508543769418921934848;
data[415]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986330444476161582688175652864;
data[416]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[417]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[418]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[419]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[420]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[421]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[422]<=640'd265568997892365958183421307639249439782679699074304056206993108584580116487809472008772454154513049201902934680709279063770125704934543825545267249188570606583274642917337242408058880;
data[423]<=640'd398353495107236126963400223035356512536489218365536640602006783478428782081433632267435611039554766374153087093880218613542213181942260498170642404010032824161659788959758458571194368;
data[424]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[425]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[426]<=640'd265568996903044352291003171397239355704090938933778659802145748928327892116220571582644985473247444956930754722318593359705568347529083688318262409318385986175701971250910153813262336;
data[427]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[428]<=640'd398353496096557732855818359277366596615077978506062037006854143134681006453022532693563079720820370619125267052270904317606770539347720635397647243880217444569232460626185547165990912;
data[429]<=640'd398353496343888134328922893337869117634725168541193386108065983048744062545919757800094946891136771680368312041868575743622909878699085669704398453847763599671125628542792319314690048;
data[430]<=640'd531137992816767098689588206552468627329593117540961209779768774219776665041523081944630313929275862236827838496002843258316710966147798256686047195211381820739689719850535202106376192;
data[431]<=640'd464745747548292448942947204772883260336491728765709340960903687623617040888630979714838395224460056055998811059991606943419003558340812870361086397939032316978126257926111479799480320;
data[432]<=640'd1731312810311731738423517647137530330245919443708482879398441392650280575745723070192214807428701314927183699982112975375459555240147258469772823085713252175416247405040893952;
data[433]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[434]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[435]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[436]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[437]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[438]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[439]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[440]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[441]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[442]<=640'd1483982408838627204363015126117883140210788094607271039484378336557383350639191203021898406367458269937586028556096836036108190205840507259805276930611359007499640632892194816;
data[443]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[444]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[445]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[446]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[447]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[448]<=640'd494660802946209068121005042039294380070262698202423679828126112185794450213063734340632802122486089979195342852032278678702730068613502419935092310203786335833213544297398272;
data[449]<=640'd741991204419313602181507563058941570105394047303635519742189168278691675319595601510949203183729134968793014278048418018054095102920253629902638465305679503749820316446097408;
data[450]<=640'd989321605892418136242010084078576565810250724560193525292073344815707069964632683637707560663098643350035920994610962411690368371714661765920491625786887328011429868730318848;
data[451]<=640'd1799565517869652802850553672994603778697120433756232925976991265676467694158133288870091067319688664337182830767822544995324267558345195980337572361199321983483904;
data[452]<=640'd0;
data[453]<=640'd0;
data[454]<=640'd0;
data[455]<=640'd0;
data[456]<=640'd0;
data[457]<=640'd0;
data[458]<=640'd0;
data[459]<=640'd0;
data[460]<=640'd0;
data[461]<=640'd0;
data[462]<=640'd0;
data[463]<=640'd0;
data[464]<=640'd0;
data[465]<=640'd0;
data[466]<=640'd0;
data[467]<=640'd0;
data[468]<=640'd0;
data[469]<=640'd0;
data[470]<=640'd0;
data[471]<=640'd0;
data[472]<=640'd0;
data[473]<=640'd0;
data[474]<=640'd0;
data[475]<=640'd0;
data[476]<=640'd0;
data[477]<=640'd0;
data[478]<=640'd0;
data[479]<=640'd0;
end
else if(choise == 4) begin
data[0]<=640'd0;
data[1]<=640'd0;
data[2]<=640'd0;
data[3]<=640'd0;
data[4]<=640'd0;
data[5]<=640'd0;
data[6]<=640'd0;
data[7]<=640'd0;
data[8]<=640'd0;
data[9]<=640'd0;
data[10]<=640'd0;
data[11]<=640'd0;
data[12]<=640'd0;
data[13]<=640'd0;
data[14]<=640'd0;
data[15]<=640'd0;
data[16]<=640'd0;
data[17]<=640'd0;
data[18]<=640'd0;
data[19]<=640'd0;
data[20]<=640'd0;
data[21]<=640'd0;
data[22]<=640'd0;
data[23]<=640'd0;
data[24]<=640'd0;
data[25]<=640'd0;
data[26]<=640'd0;
data[27]<=640'd0;
data[28]<=640'd0;
data[29]<=640'd0;
data[30]<=640'd0;
data[31]<=640'd0;
data[32]<=640'd0;
data[33]<=640'd0;
data[34]<=640'd0;
data[35]<=640'd0;
data[36]<=640'd0;
data[37]<=640'd0;
data[38]<=640'd0;
data[39]<=640'd0;
data[40]<=640'd0;
data[41]<=640'd0;
data[42]<=640'd0;
data[43]<=640'd0;
data[44]<=640'd0;
data[45]<=640'd0;
data[46]<=640'd1813962041959816781742757536418579403841941399081541595129205241096870139782246321354582145161712086162960596136900452777307423468626143427956283140613483479487741952;
data[47]<=640'd235872539078501470947974175555756220337744249944214030294279290980879917074599726974611327609305069787197239149552864111379733307796815443384959153605941188750095679488;
data[48]<=640'd3773962417791988548370103677149226631423652920863738510150696305360178916026613975223128338121084635473847781346621983765795421484438944250461034188410988560694361718784;
data[49]<=640'd30191699396814942617348174385333510972188244553048511608955201082071946107807859465551661882290367936120823902904785617779867557794976058645826975830061622645348785717248;
data[50]<=640'd120766797592531935072373005808156236018699915384542436169994929481159710550049086976932592010968789430178493407509161014415555214689087071746011741590890871100866723577856;
data[51]<=640'd483067190375399904889198940887168656892272868257506581535269944593274630081815226910258451595332557556953559505940254062790538522602779284378577852475168448031372523601920;
data[52]<=640'd966134380752557197985938099077450768744950267098787140186707701875476249819238594259240373277263892395246441606794325463355060020865034315301789976562838767992925784637440;
data[53]<=640'd3864537523013743568319552143621061928998588228176918439051889623776060063734170847070580804534859188081601159522807586342582631818176906787765234696674808217954998173040640;
data[54]<=640'd7729075046031001913041091159416230316783282707350963113123850225361022052280555797284156131167359408651648383816513631847174627801028373488254335546045482258813656481398784;
data[55]<=640'd15458148278103476642667387245335357040445284495097406982111484393174517134483113913382054231209645811926413776466261025858223266560933455671195932505963555179946191873900544;
data[56]<=640'd61832482432168273979091049387078064708532896633687211582111721653882661806661580989944292406531425412583824780140896631593018964257391714335488947692270391455018065718149120;
data[57]<=640'd123664728991270252996413132759771591613332600921374623926934903150805625840852920278508866471806135706536356880945086387264347151305418943905302445167747742736369752351965184;
data[58]<=640'd123661426774127445489736955804160157862165140287603956803514519725263277474525124592918247762007910033884974760296979536106444854753703436098601802390684907787631275248975872;
data[59]<=640'd247322853548254890979473911608283734966354826077350774408876733221179808776098672080183140498755123168458374504633306698886538314465940811478067648667588064102593928166899712;
data[60]<=640'd494630611246810495791862881006982401468569899805904430997584682961315378238158224790263059700483537161373044204668161281352966869769619201791150026315285783330674196487340032;
data[61]<=640'd989261222493620991583725762013955658305858076246370669137571076607226144026600761195660719317639482079900796423432250439597526522933522010843891362561922308716712798464245760;
data[62]<=640'd989200839094823846922089487966832334880656033253902573193918916542764079402351243671184621125641618921880401742665153674044856909389402522459630298414994460754584577536688128;
data[63]<=640'd1978401678189647693844178975933663145656098445946898780911571451282571834493621670775928655675341490544492568104068167350003542921918583024843650661985671161560704858919534592;
data[64]<=640'd3956803356379295387681655684597656654675523745518033665298526632071289086585961776349611600877686093664389338859594047827884205879731271964821350382654816926568621689265979392;
data[65]<=640'd3956320289188918230395271032880957125663518011641079276869682931273281822054764176299227030148139799816873600246619044596582092026589079441100544328090620856947507157150990336;
data[66]<=640'd7913606712758590775363311369195312166225619597260468715494691828759637423759239875231714712566710199303137630229043630766106190458105057001722903511310894763762761095608008704;
data[67]<=640'd7912640578377836460790542065761913679857357433104196928178508442616073615078459121392433718661052188226891973051492611024757433184816709901033036672147463274944218227902775296;
data[68]<=640'd15825281156755672921554275062445157767309411140678122587929197619963059058916317002734003088456879506431386007740783148363280077830514087898856060469048491623081533388967903232;
data[69]<=640'd15825281156755672921554268515663941975025671113605561509200689471784363426750967110292157627345332553289656346046531994331460655917571902188889503356968004839916318859152326656;
data[70]<=640'd15821416619232655663236388779632895086635576643789706608577930939865217363157271878512622177156541575089711669550334813391274428545187334519493585044647838222703199765697396736;
data[71]<=640'd31650562313511345843108550124890315248883982986267264363077966529810639769975311377412871845076096454423962640815162143522716372994498646622871048004920263337660513437154803712;
data[72]<=640'd31650562313511345843108537031327883664316502932122142205620950233453248505644607320555109081032837758097089252886666282953283385933269469990938464870503870437647677653327544320;
data[73]<=640'd31642833238465311326419146327546019641993802442025836156578107232408941810620616269612104332208138888985146249276515137118598274636909989131969193489327365853096022827688001536;
data[74]<=640'd63301124627022691686217100249780630354900546324990038319765718704413307032680147796501621312292324036638843155784649904598250407537216012062788963066685970039325258086338265088;
data[75]<=640'd63301124627022691686217100249780630354900546324990038319765718704413307032680147796501621312292324036638843155784598482776801987136624207038407671960251046398770473964836749312;
data[76]<=640'd63301124627022691686217074062655767185765586216699794004851686111698524504018748226734239467846136224086052383781118876919205043799980906898025133021505914042061940449897086976;
data[77]<=640'd63285666476930622652838292655092039212571339189662521675334292905422016599079881883480611381282330188772793233894949578858805293644896841232344797606300948624365242354413600768;
data[78]<=640'd63285666476930622652838292655092039212571339189662521675334292905422016599079881883480611381282330189112000263347012220829404756228684219151548413222767935656791717551680782336;
data[79]<=640'd63285666476930622652838292655092039212571339189662521675334292905422016599079881883480611381282330192278134989459089759428020327590891647614041218251279567894318467731582615552;
data[80]<=640'd126602249254045383372434200499561260638361568116413466581211935024952943623444677646277644904545844801482504370375670593386838186605878406243538999330167338578882721217721139200;
data[81]<=640'd126602249254045383372434200499561260638361568116413466581211935024952943623444677646799126114487473239566784754842270385058542970434750952764854141947926373869146829743041019904;
data[82]<=640'd126602249254045383372434200499561260638367382826207831436336330231072394478383244469544626223713690865528505699572614178639797002847017585442798125569072689065002106613326151680;
data[83]<=640'd126602249257730893333250461852180142904442913594389304363027330732322760342844031121693327218354055327662904588583280420189033139164021828760212824963920630369576961290125967360;
data[84]<=640'd126602249257730893333250461852180142904442913594389304363027330732322760342844031121693327218354055327665996570946642592759673927626858380729477533674851726811814815653653643264;
data[85]<=640'd126602249257730893333250461852180142904442913594389304363027330732322760342844031121693327218354055327666327854771286932883426536917972135989102845742913383163468834023560708096;
data[86]<=640'd126602249257730893333250461852180142904442913594389304363027330732322760342844031121693327218354055327666410675727448419636615789661392349427665482833376954333180871336777482240;
data[87]<=640'd126602249257730893333250461852180142904442913594389304363027330732322760342844031121693327218354055327666424479220141197295168529677979132497524214470020034004794304988807430144;
data[88]<=640'd126602249257730893333250461852180142904437098884594939507902935526203309487905464298426345899186194443134541390099694368187133365584563781003623807797225138701269642539780014080;
data[89]<=640'd126602249257730893333250461852180142904437098884594939507902935526203309487905464298426345899186194442342997355952151182081198737882087388562597973698949089488239363685103960064;
data[90]<=640'd126602249257730893333250461852180142904437098884594939507902935526203309487905464298426345899186194442258190422279375431853107459227684425591774754557352528219241404744238891008;
data[91]<=640'd126602249257730893333250461852180142904437098884594939507902935526203309487905464298426345899186194442236989120220327967851325786189467745284764961538141306744727302795151015936;
data[92]<=640'd63285666476931072324544221850550809387001282217243825692424193492499553574014312373301296661344368424809977348064927311154220550609374416812820879186142872588584420338558828544;
data[93]<=640'd63285666476931072324544221850550809387001282217243825692424193492499553574014314509288332582254450819829917101911410203939396324433642837652691995703303794920172534757117132800;
data[94]<=640'd63285666476931072324544221850550809410818333534962272281946957757770255402384020474856779972841846769894415083397982046269896400415623175426888816737746548047245985114941816832;
data[95]<=640'd63301124627023141357923029445239400529330489352571342336855619291490844007614578286322306592354362272772300161105078777852697042113343314704305698259446184935727968394749673472;
data[96]<=640'd63301124627023141357923029445239400529330489352571342336855619291490844007614578285279344172471105396602856184319050496599463581892504650535647177287158339781479423657732210688;
data[97]<=640'd63301124627023141357923029445239400529318859932982612626606828879251942297737448911762415795838834934717084381002062365768724531332633238653102143710870272322498739198400397312;
data[98]<=640'd31642833238465760998125075523004789864057848105044033352713536350027882442294462961500793815381876939128189805508034215360713845605000113844378918938265617849019132743916716032;
data[99]<=640'd31650562313511795514814479320349085423313926013848568380167867116888176744909741867233557125138134690567574056127777177234509990829045913112044230673334341032790525934143799296;
data[100]<=640'd31650562313511795514814479320349085423313926013848568380167867116888176744909750409095775969011950518315510457244819019738454960994267328705590393961928702799623755065133629440;
data[101]<=640'd31654426851034812773159174672240017505903171372874601752760000588744632157776596540812101288223245737293979985497092410922856751020398570116425806925331734387565595810882125824;
data[102]<=640'd15825281156756122593260204257903927941739354168259426605019098207040596033850747492554688368518917742576764377957346472148072039707963526584044286463447548534889341840114319360;
data[103]<=640'd15827213425517631222432551933849393935411503631924279822518426824666321793421909356491394153149840359361618196319872571039432305241616183107919095397817625284350299763619397632;
data[104]<=640'd7912640578378286132496474534611291940919063337614435359819615576992966193544711871638345035196581309413670275800806854244296355581680274145607875990481420267484113370827718656;
data[105]<=640'd7913606712759040447069240564654082340655562624841772732584592415837174398693704532501275368124011746440260202995725282213767128070588240916572791414992024398468929005060882432;
data[106]<=640'd7914089779949417604362329120335753168124320724311434057015456553708295321526122837417109728524211051344563610583824057249457588267280434475742978768434669937720075877754077184;
data[107]<=640'd3956803356379745059387584880056427591158073583379790865126560409900070890334050686915511852230075979122292184497629806280031234220314593285996575440993757986594748001373126656;
data[108]<=640'd3957044889974933638034129157897262814216489056302292288174393409803196206267247599481870428231013250344641858375667076171724527690345140490437504953211799474631344330668769280;
data[109]<=640'd1978522444987691654870029176678018780574071829492995382836869868755548089401107224622376542313920143777512400000835085397573982761563094480410264884678774127853208247096836096;
data[110]<=640'd989261222494070663289655162059641874455095220795504950890270306320326672721925710123607624898786371450195771923344656246454135643186343235041228912426116897182202297438961664;
data[111]<=640'd989306510043168521784206187016833502963910067119849478360109736164807967781799979114113451491072138955820130877299902960708401728910539237983238159650136127347751430119227392;
data[112]<=640'd494653255021809096745067691237820129075914274599505317324081314735845844444591023020226043289185535985016251701333380707972508015250036961288947053878592512514687618248605696;
data[113]<=640'd247328514492341794996593570910163772220114163811772491727985820399731419975138933321454737516596797631332582126307672354590867970972337650051912062418048649794375228808232960;
data[114]<=640'd123664964864800278769719248114573399258207930383252715016342337134013817956261794850132671422770737934734057017082123647682630271794541687912302854959748408882824013001261056;
data[115]<=640'd61832585640631716025202323909265334608151247552105920196560177086088338680637563965386486056796938672331991992121916092500874699838130650053946584111149357181169831312883712;
data[116]<=640'd30916300184137847084142439447397672056354963475599197500694383314880789386424484155769343204241563806662955519379816509962597645921965137779885231197036102214559216632332288;
data[117]<=640'd15458150092068813705308657633943360592187719857838238155235991608807827124748321432197963197647928166233906958927728602065826409920642968445404463846404333195023724413190144;
data[118]<=640'd3864537523017038671196414836284181790228194141581439199703162598267084297051051358025388996263287562768746452719219606897026342645281488609401857746332894743524863981387776;
data[119]<=640'd1932268761508409498829098547170715998653378385258627423793039353647114750930204168707142744792705548682858130008070844923058918901272860478236406329751020042623822310932480;
data[120]<=640'd483067190376937619565068197462752993439641857620026388700135548161098116543389634949150693228362295380351831025359417428458207669866236734478706838706296502244757500592128;
data[121]<=640'd120766797593410629172051376197032374105894483628191533227184431631830770855068527991461178137110769897616482638331877312768727736206323067018960348362134910978876696952832;
data[122]<=640'd15095849685227059801223316528469321319352992936396013180872667584106411252611270037761649744678199803674906338243973938194733855754507362449340466862942108600451351969792;
data[123]<=640'd1886980987465080948986531416536755472144091188229835651778731242562566076001477634045308530923586981390001209161136942831943944646906003643053215641577048825283951460352;
data[124]<=640'd7313434264409420040290151715434147130932702532991568418954792092702091966541137789583202805543600955543863425285056377617172288154729263647986750313658269605394644992;
data[125]<=640'd0;
data[126]<=640'd0;
data[127]<=640'd0;
data[128]<=640'd0;
data[129]<=640'd0;
data[130]<=640'd0;
data[131]<=640'd0;
data[132]<=640'd0;
data[133]<=640'd0;
data[134]<=640'd0;
data[135]<=640'd0;
data[136]<=640'd0;
data[137]<=640'd0;
data[138]<=640'd0;
data[139]<=640'd0;
data[140]<=640'd0;
data[141]<=640'd0;
data[142]<=640'd0;
data[143]<=640'd0;
data[144]<=640'd0;
data[145]<=640'd0;
data[146]<=640'd0;
data[147]<=640'd0;
data[148]<=640'd0;
data[149]<=640'd0;
data[150]<=640'd0;
data[151]<=640'd0;
data[152]<=640'd0;
data[153]<=640'd0;
data[154]<=640'd0;
data[155]<=640'd0;
data[156]<=640'd0;
data[157]<=640'd0;
data[158]<=640'd0;
data[159]<=640'd0;
data[160]<=640'd0;
data[161]<=640'd0;
data[162]<=640'd0;
data[163]<=640'd0;
data[164]<=640'd0;
data[165]<=640'd0;
data[166]<=640'd7214722814281215676076484393336843348098096790246358642812797864546946125152077138320483323038009455714104246272;
data[167]<=640'd241297722551031487448653655127651147668736199768482553359071186336407315063274642552448991132676384547940425377358337692000562661887128504912223566292631510221054057381888;
data[168]<=640'd241297722551031487448653655127651147668736199768482553363380808946651192104516644453612440992450620450936566618149368819315923153392580196932899610645776161253333091221504;
data[169]<=640'd241297722551031487448653655127651147668736199768482553378156568315926870130821216944225671857591138089362151354333594516751919611513644670771912946616549732426580379041792;
data[170]<=640'd482949254065385807159370696891556240090260311663272754577321532838133668965558001292702124553721874536734782135922242580324178442799524478372411283568289922842510166589440;
data[171]<=640'd482949254065385807159370696891556240090260311663272754695527551720884929449132618778677106622637576323631165566254773446013170873699890083221821026989242270507009212153856;
data[172]<=640'd482949254065385807159370696891556240090260311663272754853118742300013434885040015975105846201982546500732399114458542527788028643601077900859443741491585524292495800795136;
data[173]<=640'd966075412605430936829918457548382599829046804770646136881891733085991734711288357200008409700961778649217711474909133859901269953731709948516311503514925286375143543668736;
data[174]<=640'd958527487755787854125434948826885016851635058189106052083835471813395818673069421293051132678656452977801345448527378008075595348328083253180401792029187972360813225705472;
data[175]<=640'd958527487755787854125434948826885016851635058189106052713036201897048172021618876785704915163836127010122885098999115201551984921420802051643767989501563239537040657743872;
data[176]<=640'd1920917390166724817238845754124057554886160257842332866648217061092929340044868549565594826722121029175276304477673101362980524006632274563683865990863297558117264971005952;
data[177]<=640'd1905821540467438651829879535800104479322492572960667104929786985126571527957591861001920147357674969328724617494086491534627677529542564629947344198669940376777619048235008;
data[178]<=640'd1905821540467438651829879535800104479322492572960667107451515376998733031995717222037778917438223621559127529094516661353362023406360600477482020819188536907259130591313920;
data[179]<=640'd3838105044016789783323462674838680136897311382037401858490705843387298732264959194487635963667633188832644065732742411839498422117692651934169352814746859357235096282202112;
data[180]<=640'd3836218062804379012647341897548186002451852921427193643300273530277472019749340732829903660452711116433217781708634438958378062691272042493172019595447887212058340348657664;
data[181]<=640'd3836218062804379012647341897548186002451852921427193643300273529103200728362424118887152655003681749313998036247061786965134401528356920805629653771171026007724122334822400;
data[182]<=640'd3806026363405806681829409460900279851324517551663862129920775458784121432810432225118695982392896080083151754562798775412332877422493151251295542100883071398175190386999296;
data[183]<=640'd7669627766837220620759654559973311121113393223176951644331128330351373690600628477633235505866810952555968191711295992551883015815560115882326954113841178718103409845600256;
data[184]<=640'd7669627766837220620759654559973311121113393223176951644331128330351373690600628477633235505866810952555968191711295992551883015815560115882326954113841178718103409845600256;
data[185]<=640'd7609244368040075959123789686677498818858722483650288617572132189708628102264664286331498958898704598838252698005828327411742845976784902021102064030122804787376631142416384;
data[186]<=640'd15338323099584773138300970266934619003812915929119037927816708528458210396922397103755868984695469488018710849993126361592333970244774311295753405982192599622388854070181888;
data[187]<=640'd15337851354281670445631940072611995470201551313966485872763161502670679693902164834743834442840883076370618394720836852771090093325589779284583410437755079078389752927354880;
data[188]<=640'd15337851354281670445631940072611995470201551313966485872763161502670679693902164313262531253105618156653118027748500094687662479317635113735608288720474872258503119969714176;
data[189]<=640'd30675236491511504746034856288944892991066088546766839430149116824938378831672663790371727003786838104951976189488292024883136068517876937425291998869046457096641812772159488;
data[190]<=640'd30675000618859953399700341191783581224260494964610198373197205843715275413912765865834699402572914665386108863285018769216463155141012926722283843763092149315396542486544384;
data[191]<=640'd30675000618859953399700341191783581224260494964610198373039597818929697497064181616268265408359442124842404533438639355026434317328790193270762194788546689232888639248138240;
data[192]<=640'd61349768129186986633166316025654517143722315340668996043461583431468818673273112852868123460605516012647747987966178462485446101304388804853400244962619494514349647778021376;
data[193]<=640'd61349768129186986633166316025654517143722315340668996043461583431468818682013563460157128451710935478740015516107497701154328780252800458430642807311196794581161980326838272;
data[194]<=640'd61349650192861210959999058477073861260319474186880858029698196675021936006258472018106782628140754965796450395594882656155094751072265562018311928674768776055113561891930112;
data[195]<=640'd60866583002484053666912139490707362842282108270667553654866042268590496113472176840647449614657902376908665745835572882233438648141043920985977398540939423435744112942252032;
data[196]<=640'd122699183831448959743261079345418303538109487894227498547498069521332173025557178394797162743758280192489871777484346296911172276536136477459991336738023379901112149614788608;
data[197]<=640'd122699124863286071906677450571127975596407978591913794570041513611438069753929855636906808932145446869018557050394271157414910356170141864936376114103715830794902966848454656;
data[198]<=640'd122699124863286071906677450571127975596407978591913794529851467291115700957405284796956477247294168946465039797964697885971516883292282675081507867395924860935033579909414912;
data[199]<=640'd245398191449428410631366527908118145371421192484221598194276818139460119034084453455372444239444665103646664240086575730305704826465366495984130243961359521272498250418487296;
data[200]<=640'd247330401242774151967130575079293811101869235572180746686723742386962437267347432659942244522895764803850853833242709220979137957015491669652752930619925432538073661825875968;
data[201]<=640'd247330401242774151967130575079293811101869235572180746686723742386962437267345300844756003145840874459921454143534580349864051532082985930860570988667046707301624963336765440;
data[202]<=640'd494660802831050879167938923498890786933761720260456832829315864287239005032739142086744533232210163502925646736531393649172373155158895231044860105944667543573368449133445120;
data[203]<=640'd494660802831050879167938923498890786933761720260456832829315864287531426106277344293640772435354333171339051315824935733021961682906961788752006502928600706614190865446338560;
data[204]<=640'd494660802831050879167938923498890786933761720260456832809220841127370241708015033842567529394763666143401673515171306096856643579443384376930730712937293729802810590389862400;
data[205]<=640'd494660802831050879167938872352162538556545001304367819877984087742338272285127431167760412778912797942648482270061788166538893515242701503603643416451937620274791261870751744;
data[206]<=640'd985457083053862477920743409649724264699896435768186221171690574180774650734913763814498510168990043276456800959806793962700370525944855521103891545410554566952966483043418112;
data[207]<=640'd981592545530845219576048057758792277355597508438479786173072740935517232573220492358550849195317898350824006225454071797803513580215922821183474418183902383291966004532346880;
data[208]<=640'd981592545530845247035251791843662721850680757522839965637335894491820327023275744614503942485421980799730788879100992147484103405138683805990715346557972270306180069100355584;
data[209]<=640'd1970914144081036070582765379175452637447683760252341628224879874646069743189258307517738447477951547043468599710843098266405463093698651512747244149282089297480466373606899712;
data[210]<=640'd1970914144081032555806363290009822069960041192666836360406499088214395342241597719021869428807062122982426462680998490094504019705513897889543605185723341225931170383451389952;
data[211]<=640'd1963185069034998052846594093614040694370205041687784545741272951139159378435345089566041998239314350094765562137415506303002178626341373493318007175274459902103243168547864576;
data[212]<=640'd3941828277148720675848216047778154845631315647776348875372767390542368033107751429261675549059974582769039254258454722141331533631525119378691412458380847586630663687156793344;
data[213]<=640'd3941828277148718918460014849755154816755844207115329202672386002950818447430674648086787016727654832392964305910512936720004614110597577803017224265107945594472494275781197824;
data[214]<=640'd3926370127056649888513736611582358414391705567758786451034191984652620038250311526655733189248845391294005501581072306554379803036919108980792604671954798850059255590072352768;
data[215]<=640'd7883656548790764729188979940537664928491879604618321010416934801777886039777346218556158265064761841216488817188437546887136343220196733316756244599876123291614977761289961472;
data[216]<=640'd7883656548790764290605335937842097817971757008447076262156329004649676628631719766784566843548990789850516076572029415109315063125580336938470126772796203330772226250515677184;
data[217]<=640'd7883656548790764290699188956656392049597840176839668771248950865882221232237954018644790958221835538636237264753758055548134044236911685206883779776726740627251929797521047552;
data[218]<=640'd7852740247685248459145651124759219088906664089711223541210299832170481701714148275957569895644698752891621890466395046633646801489847941472987410168124682590795258096141729792;
data[219]<=640'd15767313094828192515362215964578328648987656842104267306490148420715782734974350173392734672855698186215676330983281590889805487261050268505962115280990153815908536194403663872;
data[220]<=640'd15767313094828192487902986043368595035357613487502332506222565844678639304940996432830437793424830493847412315223171819443386858439947933359724544815042153044477864221060628480;
data[221]<=640'd15705480494459916330360911479907370220602417220336705561041716437331795894373752662739660023573619804611726925940389367608297883456027908334290851645146137787875099033213075456;
data[222]<=640'd93854655509598179697018174987440922892355575173592382206496282259021134884201525033806700579885609619425952101197652660130553820650272065643946971251081216;
data[223]<=640'd0;
data[224]<=640'd0;
data[225]<=640'd0;
data[226]<=640'd0;
data[227]<=640'd0;
data[228]<=640'd0;
data[229]<=640'd0;
data[230]<=640'd0;
data[231]<=640'd0;
data[232]<=640'd0;
data[233]<=640'd0;
data[234]<=640'd0;
data[235]<=640'd0;
data[236]<=640'd0;
data[237]<=640'd0;
data[238]<=640'd0;
data[239]<=640'd0;
data[240]<=640'd0;
data[241]<=640'd0;
data[242]<=640'd0;
data[243]<=640'd0;
data[244]<=640'd0;
data[245]<=640'd0;
data[246]<=640'd0;
data[247]<=640'd0;
data[248]<=640'd0;
data[249]<=640'd0;
data[250]<=640'd0;
data[251]<=640'd11116040566782354760662814560834039153924126998909122301691829302982613491777536;
data[252]<=640'd189012119257413592134515284333917086950981151340247970757227920207850702247198916291224333625963632600111436613438956721511635782798643837272064;
data[253]<=640'd192060701826081553298053956646462627203301470031508405129734080619546080592526520452416785201696333400475709238857389842717133079938950041174016;
data[254]<=640'd192060701826081553298051375027016639437023481508801043720157571795029079696460836428810921605718176085893492280031706033102119941319938524839936;
data[255]<=640'd157122749371075511586714658745776114159588285093117234717130498115241725821626951852549106870928098175151189917444542644369811846227810714886176812040192;
data[256]<=640'd196403436665829214026911752483424994763789988301900347966313463049152771929259604897829805964465390899141370800476363169662645070069808927716408907792384;
data[257]<=640'd15829145694278690166142978472212890152219855198965399491626527148227007960710927247178222179401240160022762731119997456680786202796522419513164193828117248311415698841237716992;
data[258]<=640'd15829145694278690166143402376296614226883306331816652877463904757716381803755671751959479362129220439779595859975161515970162064384365265021384833722495262092803666734728871936;
data[259]<=640'd15829145694278690166142984226219723588585477957577490935583332074802863409787266102796372931245503104808339702293796255753326617565362294530780522511571709786697503302158909440;
data[260]<=640'd15829145694278690166142670389895191545983690398912572414885390350202979531667788809044033102395615863102816073057643098081642042513531591207328075064843485880374266018163326976;
data[261]<=640'd15829145694278690166142618220232378201222637041563744636028020753023969968805272474462551794616781303999570648551217039614682096346555270820402001283008322609251769595715387392;
data[262]<=640'd3714994261933704794416304691966621394795572027862286710809865341136366841636183442709137153527969773283742062168353131570094750774649961051007813467578668935536611164160;
data[263]<=640'd3656026099045868197693168802425603460734971862117062168612314202745354213369433848136649178188533777031800240093940041253228854988383333927814406908256630602698634297344;
data[264]<=640'd3656026099045868190737213760646301986955557421511353562722160647811769993865721472394676952541015111565417156642772787465163754051763416302306434324571570136825804619776;
data[265]<=640'd7429988523867409538887030081764393540355125061613882296183946136071018455746432227774581489533089910633855847107467177919125991520330576555190863140222086247617986035712;
data[266]<=640'd7312052198091736369992786197160439202507029841350303854831421364393792420467102337464401154097054486758973086561328025987684821886102373833552516145551942523111056867328;
data[267]<=640'd7312052198091736369992786197160439202507029841350303854831421364393792420467102337464401154097054486758973086561328025987684821886102373833552516145551942523111056867328;
data[268]<=640'd14624104396183472739960798197872844281294004296194552777022737236555257410322223523575041835033480175481145841856357539565608338238463505673189240129267237821825756954624;
data[269]<=640'd14624104396183472739960798198539721718190120811117913054529405630268169127319864085010299861912287785421275648916389844652170606275618900910422704613560852486940499378176;
data[270]<=640'd29719954095469638148902242337453130739324883525709560395859555277939194931188320687830482070652177116304271063611506135214565745939192650126463429691379049722533055037440;
data[271]<=640'd29248208792366945479872048783072404432286481564722448611724550045727566082347046238065374262811296120538283080358736351311399496138414142976753533408976277279585660305408;
data[272]<=640'd59439908190939277973780875477192404400041394157055378175785068041560324825180807745704747538432147611740595368395748712317539455634843763898914660330520911608084695089152;
data[273]<=640'd58496417584733893892702480264063815262687546439490873784154344535659823320951536834040685599939542350761665214720052070814153349104964428252671505848729967643904842924032;
data[274]<=640'd118879816381878559194764834397475709583671286678266843293616592552123450201681081675268866462908210455736029743883908799145624040121304506515114842044112542997317351899136;
data[275]<=640'd116992835169467795274922265567212505087966708281380978141629355588012313252532169862030132047606312530579499511355502686469467995697242057413796796175820621226558229577728;
data[276]<=640'd237759632763757118585932693210093711406193883877409321305131808092971515333795433046728614465079030743297292400417683860804338022498953135277561731944647080666764199067648;
data[277]<=640'd233985670338935570539607345481495318337594229371927911985804400033402749531859341597424538603695531436117146125566263015047531950405880324009684898189290163558643044188160;
data[278]<=640'd475519265527514212055138864936270615015485460570116605144080365003619707207561530816802495295124691135120508248440279344365405796780288951004197461060793027903980956549120;
data[279]<=640'd966134380747285033785585222684485626331227247675230555317475235131409134786060191930397508801699825128533696632605017918114613905689871373627936496134745144944522206117888;
data[280]<=640'd966134380747285033468066333718559864939914574877553761778012159265137150919873058929496147196947080580603118259847062634797658851083374080645989853852601905790229338390528;
data[281]<=640'd1932268761501599619589530069212212539323037883499698431014063988271495572461358911104158755212681295671788151582221047226557494937453128077934626027967968116333949453598720;
data[282]<=640'd3864537523010228791897925327383452509032343271990984740516081909444738366132339626955102032946786489994420718490061285929430855384462863497740311236827677740448680534605824;
data[283]<=640'd7729075046027487136586730437099647569591244222303764540868883876804171378842933468755103531935899718847117794336911654792494160677250731011464785397202987703039004294250496;
data[284]<=640'd15427958393113322874613821420596769957830361697840272726586536392615320227384100885077950838330227673242102365063239996555019207871497081366074772363262981248946871354785792;
data[285]<=640'd30886108485182356253395228971839202535226654313698700205583811505393597793739712083018820507949490831424771171469850208361173625260813572856391319809736748102761336971198464;
data[286]<=640'd61802408669320423010958044099295100638370575982486406262647561649353688151193536303471388628389652989271677950117328325512912815017002731659115229982977965645334124251054080;
data[287]<=640'd123635009037596556526083674354206898147153413257789366241163325672577994427826503096050488893700414236671095806569941142934464923450328784752039727527063967857030263553916928;
data[288]<=640'd247300209774148823556334934864030493164719087808226133340202621081521853009397065951778039000181968929348234934517149927354038434684116320354357136604604879643711043706814464;
data[289]<=640'd493664476866499043030676711473376270931255768926477451384469673243397107161849289927181077658231452654593145998670957675418322219836735376185844319519475804017434366264213504;
data[290]<=640'd986393011051199481979340624348420449613109035388780957150758395860209794508353317024947221860737597200107327118701958494034682852603956572806555296879177523339538799758671872;
data[291]<=640'd3950493291205436632360704985208725807967216420142600358574611029911942554533292801696693443228971785733372573014170398656554326537158100948142970524312421322648530401225605120;
data[292]<=640'd7900050639729074660639357072784172795947122661682770671164061480001918237736049858741631576031946219475176916880855128856249714420679581025770544306796088812184871380902215680;
data[293]<=640'd15799165336776350717196655519501502953658662641793489730975520836614433442607903101192828177501844875911181438542339986601888961348531529103489853502195648121871844793934413824;
data[294]<=640'd63255686119428283190055629114396033879919410461623660756072805190711825198960336847159177169268596608083112775730663936806446541493085455754889984120968426175162763002261798912;
data[295]<=640'd63193853519060007056540503586047480282265788972128346787645175730118066578294160929443800229932802429497751744152901690808882653261534425235880884885443302572167477545524002816;
data[296]<=640'd31411896929766074429765927998327512414680475606092761390844454743443812850340750164431753268938225055719583841490645183036016904128574015219613444747914445283140489991642152960;
data[297]<=640'd15335420834014279715833368880549897738936778379582332020441630361808043875176616337053033427374548392021857830071377978056075574230126925282281300515784567774601143358312153088;
data[298]<=640'd5936865578036307421534269808412696621459917100546585276108082013635903278063615901289642090913516277742591432664917126951514843878206523332174711802975253175165019278423359488;
data[299]<=640'd935942681798604082209303941164060616764722117501118170568667406369875506851089202048467386352090217976389359991689630600989697251333345093125332342226884070741952063078400;
data[300]<=640'd935942681798604082418698646612916944919571968532698082109827468058603523696423905487051212397217995478215468535143173842525098539795505882170069877505376658064582891274240;
data[301]<=640'd935942681798604082412151865397124661179542729823420841259696629832189013328175763599486898744524921814445222657577940765933638501965209280159118463301414476609676145328128;
data[302]<=640'd935942681798604082831145863207830820541231011017353532743426811725701306382037058715792024684323264839504214078955887868502500409268332935356693435358484126451476199374848;
data[303]<=640'd966134380747285034181665117873637489418504261307676934101576774160824368117015824339361024744935356653396394737923728851976178091996278875477814146021160821312394107027456;
data[304]<=640'd966134380747285035019653116616917443714639098235294365167345195564428455034476069498132466795448007647300253724658854499040154586980864972309200827528781188883846508052480;
data[305]<=640'd966134380747285035019653193880402463234471315955788281038113844341031496161944101673342475050443277339811843007966802758131418332875061366793051475716902941766126292434944;
data[306]<=640'd966134380747285036669442160546614194575222467963473795042492388722853627632519207374822363708417363419166174586752386989556415957396224712599245563182966606877209187581952;
data[307]<=640'd966134380747285036669442359167486868457705730555379193273558482639571497298808006344067292822181110722465134125704660227158348303849713141365352724775017091847374589919232;
data[308]<=640'd935942681798604088657781941309033844012369389162468039473175703539187541233103710188647061303637464504603079777421075483582492973692581645214800996129206720075161065750528;
data[309]<=640'd935942681798604088605410079720193942625088983199403619587894457380736017914349484262780158812858356116356453336942395607691644816030765587683735367580372240838563358310400;
data[310]<=640'd935942681798604095309323622216021091342616906831477830537243923026985864474952921405084315891741705744733582530639314529026977223760427192396509695408047360439587210002432;
data[311]<=640'd935942681798604095309361907340224338771113048088802880608764615471167063745539308141792353861254595936035199552155024408688456542237001156764692637810601130819334640238592;
data[312]<=640'd935942681798604088500862783205037781920184934045247752601511384321003798687828726202882664546777853718303257737263966086777727057825920022195559909754228769612128308953088;
data[313]<=640'd935942681798604083472934210100840697084604423298418744343716446475886280398891241901527933592890044982566800554797788131479848471546357492710085073476556601081794335342592;
data[314]<=640'd935942681355742255984495629587131852612497185659254309952120522796230955426282866554528844422672973667223031105363157494881595514822404675414198035277641745087379009437696;
data[315]<=640'd209541752292570688851543356687898631514366531843470583351631868362460900406088972371085122980747456632022133445622865739316080926720488353839733545107456;
data[316]<=640'd332306998946228968225951765070086144;
data[317]<=640'd0;
data[318]<=640'd0;
data[319]<=640'd0;
data[320]<=640'd0;
data[321]<=640'd0;
data[322]<=640'd0;
data[323]<=640'd0;
data[324]<=640'd0;
data[325]<=640'd0;
data[326]<=640'd0;
data[327]<=640'd0;
data[328]<=640'd0;
data[329]<=640'd0;
data[330]<=640'd0;
data[331]<=640'd0;
data[332]<=640'd0;
data[333]<=640'd0;
data[334]<=640'd0;
data[335]<=640'd0;
data[336]<=640'd12486994201263968925526388919172665222994392570659884603436627838501486955279062480481224412253967884639307724485626491581791902717153141225160704;
data[337]<=640'd24583769833738438822130078184621184657770210373486647813015861057049802443205654258447410561624999272883637082581077155301652808474395246787035136;
data[338]<=640'd103194285053714021350404760941418638612197208826611871551409759305240008668127137988274057003664046939532693258265023287268461665189253466598997919925001439490607153152;
data[339]<=640'd1879610192049791103167229671742809209658532758605963596345746412613391819799528292038446745933603180298896651916523211813861195166022236609980848880060967327858019008512;
data[340]<=640'd936119585844405765106890194035409463806946713658222731621010377972732752497117110739029164244074899722046452979955500587464316282706200606151093622819742107439244247040;
data[341]<=640'd936119585844406131726638278403298905284192758349327779884919534795989174625750337506014361567625046648296793481221101486772938569434153638483826761983764080234334257152;
data[342]<=640'd468059792922204532342462101034805702346815108358041542638130231405978830658686520594423926552723367672095607727257610740782268951981730241129018772842980134521944408064;
data[343]<=640'd468059792922204532342661892936071664439800802323225451520314977185615739561326776552944137710863728696199252753061667253277437312531366067164274460739954129467579826176;
data[344]<=640'd469902548012448587593465051899033040579389063548152353131568013914982496765588538365555049338399168177069712532008739582342922351965525066432768883521332835915562745856;
data[345]<=640'd234029896461102266172704518837077598373465627564580942651463794537186310983916629732286004362121917110875684556946174311654407971227039521499301577126676964396066930688;
data[346]<=640'd234029896461101847180280069352643394134363865456664729665630929325396162368650452136203510226641677539044854814052802252046183384233006663641509246486603781806015643648;
data[347]<=640'd221130610829387594514632418835439030514932696987211060503791470006224685845667929043407116481322261338083940923498286422264986210957293474723930288476416220228499800064;
data[348]<=640'd412459803496882007156636985350405067566321749952983352020423717238038891664052742141534630254119475087655947664758319185403766769199937102740173398999040;
data[349]<=640'd412472390387036881236604112508740665005120516188641965329873093458215428325433795107271476648408634421137394222904077470094261604036295837392689602494464;
data[350]<=640'd63316582777114760705759253061333735025836994473930064820872926394046776640011934453215000944887200638147412984890393696895381057226689788826285116181267727796631768018341330944;
data[351]<=640'd63316582777114760705759256487365383664744527809453356600519334875711798513342299474937601448303053561331914986187539578399364620239951705204431888671426070349836376796720791552;
data[352]<=640'd63316582777114760705759256386670215172629032683900685066159455911796310150105431646612870428031272054109058601459298303382969163425852149149007197436098940356557902721587347456;
data[353]<=640'd63316582777114760705759141741278846435097757143827162580792273199247150688703468727900345623595262037265077806929424107849090199168001025306832710553590384073612136535734353920;
data[354]<=640'd63316582777114760705759050067161802249983940504907118028166797350750474494355780444863378571910678743068901105347678285310595303534868788814922161400774736709059418415115010048;
data[355]<=640'd55402024789952463460478806407744010249878908104347936016961931089382957058403315461468049761437378524394127064830161389720731897547423459018783483143627821353153126233691652096;
data[356]<=640'd14859977047734819074457314900780139040054779592552525880950949644047727865446154033267378431106796597527803394570532705323638554668826104470815819442654932662412547981312;
data[357]<=640'd14624104396183472739942217739468372234372818599327207487244635453103478932726803244818012804890808015219389653520179876983971544105029611938827618855719352581139724238848;
data[358]<=640'd14624104396183472739942217739468372234372818599327207487244635453103478932726803244818012804890808015219389653520179876983971544105029611938827618855719352581139724238848;
data[359]<=640'd29719954095469638148908436063421447798040503480992969200749460654085975582295398653162519705601443085385263153643235256583053882624728782469073355861450136755737305546752;
data[360]<=640'd29719954095469638148908436063421447798040503480992969200749460654085975582295398653162519705601443085385263153643235256583053882624728782469073355861450136755737305546752;
data[361]<=640'd29719954095469638148908436063421447798040503480992969200749460654085975582295398653162519705601443085385263153643235256583053882624728782469073355861450136755737305546752;
data[362]<=640'd29719954095469651553442975398122405502052138699477726914550412747453610189707628309170014360136359615971800404937832520335208078233216477369538394006632026462865189765120;
data[363]<=640'd29719954095469651553442975398122405502052138699477726914550412747453610189707628309170014360136359615971800404937832520335208078233216477369538394006632026462865189765120;
data[364]<=640'd29719954095469651553442975398122405502052138699477726914550412747453610189707628309170014360136359615971800404937832520335208078233216477369538394006632026462865189765120;
data[365]<=640'd30191699384513238614525880627355130111572562025028350433097291531880716919566759057677364606154575885462403714198168556237991816093339911519138308542710567793198624669696;
data[366]<=640'd30191699384513238614525880627355130111572562025028350433097291531880716919566759057677364606154575885462403714198168556237991816093339911519138308542710567793198624669696;
data[367]<=640'd30191699384513225311466450137434570377969634117665395824664016412865412459470639114989616017557184839852748501723673895034507521689211330060207706064473199066062501445632;
data[368]<=640'd30191699384513225311466450137434570377969634117665395824664016412865412459470639114989616017557184839852748501723673895034507521689211330060207706064473199066062501445632;
data[369]<=640'd30191699384513225311466250723554565800708724770131668637603790105901300754666709683070151057256603271083166341470339077936807750965448883807674904904498787257889503313920;
data[370]<=640'd29248209228199219427725500347164134975847830730021206464952146357092675231548179701090627581219300058126941546150035138882956890957575235820236230363108211037011332562944;
data[371]<=640'd59439909076662929699977575666342705661280415303022095446299248287707993624990522442323048367716106161318476776426499844369707475296166572605985535206418257383758543978496;
data[372]<=640'd59439909076662929699971382117227810126937498631589255895299970868711083867267343639239890581753819441900495522799854111930097105358432351731658765217117822610523281162240;
data[373]<=640'd58496418470457544361910994264649424900562105898514942794340917444788581425364328383737592978536996541272648886387935613466457456057468924724409579511794195022287193767936;
data[374]<=640'd58496418470457544361910994251692948983723270953815930854281389320343716087155219603316287237904350164335145091943305791181456599192952853175602795033616561587741087760384;
data[375]<=640'd118879817253543100389828380412073520791407393117176191375232756704194390862149526002168819433802967497244918520317009386880161025300028419090608190700053805595971685449728;
data[376]<=640'd118879817253543100389828380363296571834147027143100466526852398288176812274051946374501757685245900281906085588956895805459881729623302818573892633497283818996318672519168;
data[377]<=640'd118879817253543100389828383485033213624480399301402936198750266970484104878969596214559065375194263507575255797687222554776958587192086406826518463885996467371520756285440;
data[378]<=640'd237759633635421652985437358932105025698692605224856472086528013895809092172854222588696729111795184024598532043798695045915653883107286688788305243370022602197186853732352;
data[379]<=640'd237759634535204411894076647981196508539906400704801899813466681077348283552559528767909946233594822879604790282378485151684685032580785294003909331036773203474413030211584;
data[380]<=640'd237759634535204411894076647786087224145156886243452072951393786968060899635998831839212636257009089203369439024859353710216436835091602098915995400071274723518895198568448;
data[381]<=640'd475519267298961517085294660920094826326076451534208408215953959594478298982748055579528558384030843944438855829556306748757600641328939414906978269994145126710678313238528;
data[382]<=640'd475519267298961517085294760035611365727992433095754384686774492808886489130587278591023572386681876090811801081884025024204350632082034109719242976955742829297086620499968;
data[383]<=640'd958586457676118810172213944633142728830865042040482851384989314276308441142450411214514729420527613391236630725259341703115154113722533776007660422085583557690326171779072;
data[384]<=640'd1917172913580790313641569204666228914347421520306679341727371313058642959426826936008052548911902973734446200808356754066373017052689421280269286018777687888251099969224704;
data[385]<=640'd1917172913580790313641571595925618549432827468447839353606208926149400638060822662098995337977400404796740091477765886453677416841855052055345189533997833715506653050175488;
data[386]<=640'd3834345825362015109364395923200027280842975694711999959487904121864719935967664676554894669863429448340274898454516908112472099198504243156676153324987586112753689440550912;
data[387]<=640'd7698883348379273454059786149204592828250024412511538095205794211802058753066785454837503287445967197615894655988732674395675301602522464039753826514796798103104013889175552;
data[388]<=640'd15397766696814783330449797637538519338922430093153095428327735304701983912433417159739433177984753124200863204397205470105253924853731706723395426350485955549881591381622784;
data[389]<=640'd30795533390086672047595333634941764513117285412848291201975735632293567521978713492224130850904906492412107416957703442731418120634450438424045898855353805140780175513878528;
data[390]<=640'd61591066776630449481991163918992571283597959499466981980311272633135452107854486107534006838962963964416016050353958639543829136033764690447237989968232051509000884619051008;
data[391]<=640'd123423667144906582997328743818262377007243887290128880121408330705113009239115693467567291641617848417627674023890057259761395769882259319456579181135675887945165889167425536;
data[392]<=640'd246847334289869402417928697695322252626625356686373858834957546020890676257887611593209603760989454205741184775211553075245715963676143335337117421394959935945043498718199808;
data[393]<=640'd493694668594191565400827797370885223038317322265034216567301205121426030372491224145644035640017338419132178829647412014835658831130512831212170903340121265986952744799305728;
data[394]<=640'd1976710946708725350963299286672164676148107795911199862787115217498413976215782181343775414149695720218456777283633729430514315285638738475562364842023535963634835240005926912;
data[395]<=640'd3953421889732052994281626587983486276523919167846695155758435086437208502460703576078368598563950909143727347111603769081434235989671333980848456512290590087747394990275297280;
data[396]<=640'd7906843773935953190673326155371278243852477584136084343978658466003304993138157831379940295403592696708817048500736091030857739965444739548752116190216099701277375518528765952;
data[397]<=640'd1963185062613919838544452729233429772571284765570758674377004907073851016543271405661708395754259159332723819893632272015785646419324897255714309813876233407283959487723995136;
data[398]<=640'd463744503682998655109367497244512719043213053988414209533545644510821127240487781337190104336047914036294990087310415077078494950507592422189309980023956366328937837720764416;
data[399]<=640'd185497802022606814633026942452041918168985500270727925295288624660160480823578481261124053430602171029983405472221956992371000276205777865844086562071806131222053244993798144;
data[400]<=640'd123665201168447991307236101280230692290600533995862163865656013411966737612432679706145085286312986608093570464020812102345842109380638305970259318910986728819962665955753984;
data[401]<=640'd41275650395045429487781333014985642928738891032254619587902570652204414333175445970408237443837203149358264764501885714432;
data[402]<=640'd0;
data[403]<=640'd0;
data[404]<=640'd0;
data[405]<=640'd0;
data[406]<=640'd0;
data[407]<=640'd0;
data[408]<=640'd0;
data[409]<=640'd0;
data[410]<=640'd0;
data[411]<=640'd0;
data[412]<=640'd0;
data[413]<=640'd0;
data[414]<=640'd0;
data[415]<=640'd0;
data[416]<=640'd0;
data[417]<=640'd0;
data[418]<=640'd0;
data[419]<=640'd0;
data[420]<=640'd0;
data[421]<=640'd0;
data[422]<=640'd0;
data[423]<=640'd0;
data[424]<=640'd0;
data[425]<=640'd0;
data[426]<=640'd0;
data[427]<=640'd0;
data[428]<=640'd0;
data[429]<=640'd0;
data[430]<=640'd0;
data[431]<=640'd0;
data[432]<=640'd0;
data[433]<=640'd0;
data[434]<=640'd0;
data[435]<=640'd0;
data[436]<=640'd0;
data[437]<=640'd0;
data[438]<=640'd0;
data[439]<=640'd0;
data[440]<=640'd0;
data[441]<=640'd0;
data[442]<=640'd0;
data[443]<=640'd0;
data[444]<=640'd0;
data[445]<=640'd0;
data[446]<=640'd0;
data[447]<=640'd0;
data[448]<=640'd0;
data[449]<=640'd0;
data[450]<=640'd0;
data[451]<=640'd0;
data[452]<=640'd0;
data[453]<=640'd0;
data[454]<=640'd0;
data[455]<=640'd0;
data[456]<=640'd0;
data[457]<=640'd0;
data[458]<=640'd0;
data[459]<=640'd0;
data[460]<=640'd0;
data[461]<=640'd0;
data[462]<=640'd0;
data[463]<=640'd0;
data[464]<=640'd0;
data[465]<=640'd0;
data[466]<=640'd0;
data[467]<=640'd0;
data[468]<=640'd0;
data[469]<=640'd0;
data[470]<=640'd0;
data[471]<=640'd0;
data[472]<=640'd0;
data[473]<=640'd0;
data[474]<=640'd0;
data[475]<=640'd0;
data[476]<=640'd0;
data[477]<=640'd0;
data[478]<=640'd0;
data[479]<=640'd0;
end
end

//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n) begin
        red <= 4'b0000;  
        green <= 4'b0000;  
        blue <= 4'b0000; 
    end  
    else begin
        if(data[pixel_y][pixel_x] == 1'b1) begin  // 有字部分
            if(choise != 4) begin
                if(pixel_y >= 50 && pixel_y <= 100 && pixel_x >= 0 && pixel_x <= 300) begin
                    red <= pixel_x[3:0];  
                    green <= pixel_x[5:2];  
                    blue <= pixel_x[8:5]; 
                end
                else if(((pixel_x >= 438 && pixel_y <= 60) || (pixel_x >= 560 && pixel_y <= 170)) ||
                        ((pixel_x <= 100 && pixel_y >= 300) || (pixel_x <= 200 && pixel_y >= 400))) begin
                            red <= `ONES;  
                            green <= `ONES; 
                            blue <= `ONES; 
                        end
                else begin
                    case(choise)
                        0: begin
                            if(pixel_y >= 125 && pixel_y <= 180) begin
                                red <= `ONES;   
                                green <= `ZEROS;  
                                blue <= `ZEROS; 
                            end
                            else begin
                                red <= `ZEROS; 
                                green <= `ZEROS;  
                                blue <= `ONES;  
                            end
                        end
                        1: begin
                            if(pixel_y >= 190 && pixel_y <= 240) begin
                                red <= `ONES;   
                                green <= `ZEROS; 
                                blue <= `ZEROS; 
                            end
                            else begin
                                red <= `ZEROS; 
                                green <= `ZEROS;  
                                blue <= `ONES; 
                            end
                        end
                        2: begin
                            if(pixel_y >= 250 && pixel_y <= 320) begin
                                red <= `ONES;  
                                green <= `ZEROS;  
                                blue <= `ZEROS; 
                            end
                            else begin
                                red <= `ZEROS;  
                                green <= `ZEROS; 
                                blue <= `ONES; 
                            end
                        end
                        3: begin
                            if(pixel_y >= 330 && pixel_y <= 400) begin
                                red <= `ONES;  
                                green <= `ZEROS;  
                                blue <= `ZEROS; 
                            end
                            else begin
                                red <= `ZEROS;  
                                green <= `ZEROS; 
                                blue <= `ONES; 
                            end
                        end
    //                    3: begin
    //                        red <= `ONES;  
    //                        green <= `ONES;  
    //                        blue <= `ZEROS; 
    //                    end
                    endcase
                end
            end 
            else begin
                red <= `ONES;  
                green <= `ONES;  
                blue <= `ZEROS; 
            end 
        end   
        else begin // 背景颜色 黑色
            red <= `ZEROS;  
            green <= `ZEROS;    
            blue <= `ZEROS;  
        end
    end
end  
endmodule