`timescale 1ns / 1ps
`include "Definition.h"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:22:56 11/26/2014 
// Design Name: 
// Module Name:    tetris_vga2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tetris_vga2(
	clk,
	GridA, GridB,
	HSync, VSync,
	R, G, B
    );
	
input clk; // 100Mhz clock
input [199:0] GridA; // blue grid
input [199:0] GridB; // red grid
output reg HSync;
output reg VSync;
output wire [3:0] R;
output wire [3:0] G;
output wire [3:0] B;

reg [11:0] RGB;
assign R = RGB[11:8];
assign G = RGB[7:4];
assign B = RGB[3:0];

parameter HPULSE_END  = 96,
			LMARGIN_END = 336,
			LBORDER_END = 352,
			RGAME_END   = 512,
			RBORDER_END = 528;

parameter 	VPULSE_END  = 2,
			TMARGIN_END = 76,
			TBORDER_END = 92,
			BGAME_END   = 412,
			BBORDER_END = 428;

reg [9:0] HorizontalCounter;
reg [9:0] VerticalCounter;

wire [5:0] ShiftedHorizontalCounter = HorizontalCounter[9:4];
parameter SHIFTED_HGAME_START = 22; // gamestart/16

reg [199:0] GridA_Buff;
reg [199:0] GridB_Buff;
wire [9:0] a = GridA_Buff[199:190];
wire [9:0] b = GridB_Buff[199:190];

reg [1:0] clock_divider;
wire pxl_clk = clock_divider[1];

always @(posedge clk) begin
	clock_divider <= clock_divider + 1'b1;
end

// HorizontalCounter should count 25MHz clock pulses from 0 to 799
always @(posedge pxl_clk) begin
	if (HorizontalCounter < 799)
		HorizontalCounter <= HorizontalCounter + 1'b1;
	else
		HorizontalCounter <= 0;
end

// HSync is active for 96 clock pulses
always @(posedge pxl_clk) begin
	if (HorizontalCounter < 96)
		HSync <= 1'b0;
	else
		HSync <= 1'b1;
end

// VerticalCounter should count HSync pulses from 0 to 524
always @(negedge HSync) begin
	if (VerticalCounter < 524)
		VerticalCounter <= VerticalCounter + 1'b1;
	else
		VerticalCounter <= 0;
end

// VSync is active for 2 lines
always @(posedge pxl_clk) begin
	if (VerticalCounter < 2)
		VSync <= 1'b0;
	else
		VSync <= 1'b1;
end


// 存储图片
reg [0:639] data [479:0];
always @(posedge clk) begin
data[0]<=640'd0;
data[1]<=640'd0;
data[2]<=640'd0;
data[3]<=640'd0;
data[4]<=640'd0;
data[5]<=640'd0;
data[6]<=640'd0;
data[7]<=640'd0;
data[8]<=640'd0;
data[9]<=640'd0;
data[10]<=640'd0;
data[11]<=640'd0;
data[12]<=640'd0;
data[13]<=640'd0;
data[14]<=640'd0;
data[15]<=640'd0;
data[16]<=640'd0;
data[17]<=640'd0;
data[18]<=640'd0;
data[19]<=640'd0;
data[20]<=640'd0;
data[21]<=640'd0;
data[22]<=640'd0;
data[23]<=640'd0;
data[24]<=640'd0;
data[25]<=640'd0;
data[26]<=640'd0;
data[27]<=640'd0;
data[28]<=640'd0;
data[29]<=640'd0;
data[30]<=640'd0;
data[31]<=640'd0;
data[32]<=640'd0;
data[33]<=640'd0;
data[34]<=640'd0;
data[35]<=640'd0;
data[36]<=640'd0;
data[37]<=640'd0;
data[38]<=640'd0;
data[39]<=640'd0;
data[40]<=640'd0;
data[41]<=640'd0;
data[42]<=640'd0;
data[43]<=640'd0;
data[44]<=640'd0;
data[45]<=640'd0;
data[46]<=640'd0;
data[47]<=640'd0;
data[48]<=640'd0;
data[49]<=640'd0;
data[50]<=640'd0;
data[51]<=640'd0;
data[52]<=640'd185610707941024670611867973754967943496578310864896;
data[53]<=640'd1122433257470133446534986086890146351018105410420736;
data[54]<=640'd294239143846250660804807983768994727295789833808469032960;
data[55]<=640'd882717619341712379435433039071355923020125151743096913920;
data[56]<=640'd98079903149150447092893500239687948245382190378176742400;
data[57]<=640'd98079717539184093128501146813124149863244567699483853824;
data[58]<=640'd11694867681144940833069543012628525652481719403520;
data[59]<=640'd46819522602305280187712041018123711678985061662720;
data[60]<=640'd561273807846106679845714843837175089682921099233280;
data[61]<=640'd196159803421014103305810932127573547686497280029448345600;
data[62]<=640'd214549749934240722076850218749538070761618950704546856960;
data[63]<=640'd687133062325836809285545039454565675358892958818194491392;
data[64]<=640'd3139125553566837060302816234439929309539207229673440282624;
data[65]<=640'd176266286834233558213347784143678105190400;
data[66]<=640'd9223372036854779904;
data[67]<=640'd9223372036854775808;
data[68]<=640'd122880;
data[69]<=640'd0;
data[70]<=640'd0;
data[71]<=640'd0;
data[72]<=640'd0;
data[73]<=640'd2787593315969827365807629488677645134594048;
data[74]<=640'd392318858461675910519186287934157228081341079131978203136;
data[75]<=640'd5444517870735015416594585339625702686720;
data[76]<=640'd5444517870735170157918904391442653773824;
data[77]<=640'd784637716923335095479473677901113044518858024596973551616;
data[78]<=640'd795365232477448712162278388377722457166639424699319189504;
data[79]<=640'd871606932415181052160261366418047227472046871227624587264;
data[80]<=640'd11769565848493753646853800856673919055261502021971013009408;
data[81]<=640'd24520024040039994183870494074304220983351112404685553664;
data[82]<=640'd1619081588981253807811950154973809763985643760056635752448;
data[83]<=640'd1618315297371480734226510033318457735685567803283965214720;
data[84]<=640'd1618315314539118826135215037068739474491222550194836996096;
data[85]<=640'd42909922189189629062283024313458242811705956638639783936;
data[86]<=640'd93811563615648108505258443605164303419450564018176;
data[87]<=640'd374144419156711147060460229976541273862918572605440;
data[88]<=640'd0;
data[89]<=640'd5137934733362173992501248;
data[90]<=640'd0;
data[91]<=640'd0;
data[92]<=640'd0;
data[93]<=640'd0;
data[94]<=640'd0;
data[95]<=640'd0;
data[96]<=640'd0;
data[97]<=640'd0;
data[98]<=640'd0;
data[99]<=640'd0;
data[100]<=640'd0;
data[101]<=640'd0;
data[102]<=640'd0;
data[103]<=640'd0;
data[104]<=640'd0;
data[105]<=640'd0;
data[106]<=640'd0;
data[107]<=640'd0;
data[108]<=640'd46402676985256167673249403042541230250612785938432;
data[109]<=640'd93627448641510968846460666912887908465609896099840;
data[110]<=640'd882717455014122032042036011285265715417263690190847737856;
data[111]<=640'd3187590725183736530051724681248103706164086704188560506880;
data[112]<=640'd73559833094997449037266686166583376797466849876759281664;
data[113]<=640'd49039904812400458224906611002570703601236969308551118848;
data[114]<=640'd49039906999477758342595859178561834462660427395744399360;
data[115]<=640'd98079778922918986813801685606764021612684995811848716288;
data[116]<=640'd196159475998908480518349073309746515843398397693830103040;
data[117]<=640'd11440293223736796032436189862207349359370043392;
data[118]<=640'd1569275433863819472215298320071369763955930664912845537280;
data[119]<=640'd12548839736397469741716468429177477100311317350418265145344;
data[120]<=640'd18831305252939512678612015704954464893649289513096846508032;
data[121]<=640'd12554203517541413988105112824283269426702568884163177349120;
data[122]<=640'd0;
data[123]<=640'd0;
data[124]<=640'd0;
data[125]<=640'd0;
data[126]<=640'd0;
data[127]<=640'd0;
data[128]<=640'd0;
data[129]<=640'd0;
data[130]<=640'd3138550867693340381917894711603833208069624466305726808064;
data[131]<=640'd3138550867694054005764247691544362351644645024232623833088;
data[132]<=640'd3138550867694054005764247691544362351644645024232623833088;
data[133]<=640'd3138838210607252736078836901671462576667780788762215186432;
data[134]<=640'd294623027712326907953429844294149609519652397092192649216;
data[135]<=640'd767007752869800195825281488732725841423417885241376768;
data[136]<=640'd11713444114796345417654357581738937491162277085184;
data[137]<=640'd1534003812027463533315142096340281850679823428879384576;
data[138]<=640'd1573108204352550835891144337281044203514971762128247062528;
data[139]<=640'd10206421798744587020501226269911623980920209113455974678528;
data[140]<=640'd6681707122431982035149763662740426199350800087901347512320;
data[141]<=640'd6498451560073430133808531084818851995792305231004937748480;
data[142]<=640'd23386880692679858611100302060311768371943471841280;
data[143]<=640'd0;
data[144]<=640'd46768052394588893382517914646921056628989841375232;
data[145]<=640'd0;
data[146]<=640'd0;
data[147]<=640'd0;
data[148]<=640'd0;
data[149]<=640'd0;
data[150]<=640'd0;
data[151]<=640'd383123886643719949830842502963171198276005845899673600;
data[152]<=640'd3138550867693340381960430007468950515984099548160988282880;
data[153]<=640'd3138550867693340381960430007468950515984099548160988282880;
data[154]<=640'd3139317115466627821775021100744642242514807907994845577216;
data[155]<=640'd766247773421244626064643935479404303718857434661388288;
data[156]<=640'd294239706892700142262611992250434331888545500364623839232;
data[157]<=640'd392319001688828009145725346667416355209245948235724357632;
data[158]<=640'd786173302078662307567016816416583468884417689659807629312;
data[159]<=640'd7846383249085871242123050343055842839240805026049743126528;
data[160]<=640'd9476970389494926441912203448650212961697772718390180315136;
data[161]<=640'd6326141785615822218157936416370519179917100513290071572480;
data[162]<=640'd6474033772843262703984869594755675905635893045564299804672;
data[163]<=640'd392321857103517053741231290641865528154775280155984134144;
data[164]<=640'd2353913150770005286438421195962151735251746683252023230464;
data[165]<=640'd7729075046034516689390703781863974688597854659412869997314470502903038284579120849072387533163845155924927232063004354354730157322085975311485817346934161497393961629646848;
data[166]<=640'd246364267092350219474328683046914193199056617268785231164398747280034345320959477064182352619597564345107055522008263795057023764641490463053610427933526397729432526944993280;
data[167]<=640'd14183349061011450654150588248978885130701596693501525615317193411479683556692524573464857490742551226803348524756297036301811056513318292405303509311456934775901580358875369963520;
data[168]<=640'd31912300073170651499092428594791257763536706108506497228570095062614055087400406815030704079997171982928060435065548413491817686659473312841262670480229657914314842180372154810368;
data[169]<=640'd49135152398600089336961536738399769954196170839157165120996735411585050945903793590612541767762748612251073442825700274910885435634435871110962700627801144593418344663775843450880;
data[170]<=640'd98017038194366425043894141533883491354641007030816361447937759410644121515613558857007962190637660133641367607125437020923278240690259535628333564448354684479735968850114955444224;
data[171]<=640'd98016048812377133828613237887934539470068564250749217073915056304400449122783146131264899291655387558618868935776238955873699316833792954544697012142751328884141165724636035416064;
data[172]<=640'd195274277259544825665578930642498661625916410484184636188667661691427435946857381971951353722114619526678975536137290960688570671603387684862354292336024720096055064124810875371520;
data[173]<=640'd130182851491267367411099788352699556093324531425788739244112679414113465430255757998398973739731906117075348620592320473669325068136509451388537024360437409724972591908609668939776;
data[174]<=640'd130190766071662431605832807137855293965382193410793820463822810288660850741950415342932721568738119344870333281160889740189712001617148436687105571102523538809211315412617217966080;
data[175]<=640'd390544597149638908312538983495346808115050343266611386138735008949680846932709327861400707635917471210729624623619461412470907133571273599847003666017216256369904149580980674363392;
data[176]<=640'd260365702959890960273270328591949784700719449506075951165726716257969693059037771022445054366947051883084744635935830697154067066874395394997525292925506213941349007555322965917696;
data[177]<=640'd262407662758226873731295378757729546482637762815172477336473661277448858849762922280195335426194801187696521778770488318570515781497402517616942146614588878187101209109832021311488;
data[178]<=640'd261394604189185777990342580944015771561255179550542898185614025793101629255393818434212164681614787743428323615837917516903814960906228552226293889848258833835840705903528584937472;
data[179]<=640'd265438974584366311812007279426759374371132131201975808643803151661898599820890574049738778755955054329374014759085781620331723693308319346899982596001800615903482645610711604002816;
data[180]<=640'd263412837414091569377360186101160108642635691685698812371618086872301098928379312380246330393634370197824880323106505353703833324143708200477886788833047520596211039507114335666176;
data[181]<=640'd782133964519762194298163688470438126584941615284886442011889870266069693477481427710375006161496562262403430180935378252413955100314408511746174466494734480423451489193900346703872;
data[182]<=640'd530893764180937621357522066870242100361359514326424124385791399090494550644325477980379006699033442423295279326343763783370566724337994886809054706014956481354265270587855225225216;
data[183]<=640'd530877919577093250598308815927489279213247888724372328002296904425963599415842090782638408304590456540725633225518034624444139527515484610559666160089395266323195612966514449186816;
data[184]<=640'd526825720111958274188395057748733634563509805483535348520104873830701594504002949303886736968703315802377312376292042701543041600634661375423360375770744624133341906763323199717376;
data[185]<=640'd526825720111958274188395057748733634563509805483535348520104873830701594504002949303886736968703315802377312376292042701543041600634661375423360375770744624133341906763323199717376;
data[186]<=640'd530941267076170549497095062135685436349795636741160875884794893826205392717622501257117405592812267415623593929112023008132430895884896427213319097848370738710828253876031034753024;
data[187]<=640'd782149932909574099203933292936181204148272862961954268054630415670167292762437341370597952980896133972180651641923808420394495009612094649528761360435339142446951378515407847555072;
data[188]<=640'd782149932788807301609643969664451457556648258452612789001304321962128691154577368174049189714140078766495571080596820419410051972819435941371167996193373246401105105118627197091840;
data[189]<=640'd267386053461331119061225060677968885335030993449771251735307560893493937691988339823041331001320109602524804340948045435107780263546857039032484499584229842589722876816412223995904;
data[190]<=640'd261117711766396757749995684785246946950780624538150138864525546799875550418888396181476832132823965870308440956327092399691259268139309260927030553642947553840091994436607965921280;
data[191]<=640'd259345095503639803120120002847477615089546465215190627927818019125089365653709721468759754086954368200978477813178762734952786256000021553857578409868547467075100364623752443461632;
data[192]<=640'd389017457031170833073632748587826401058685409972766781052682310677922266010363101043750599366551361772484661769781912396910432064137956860372837157813642117540488137170052731371520;
data[193]<=640'd129672611763883570170633647468866832977296025894954594057363335465567844443009091148812631702315633201348424561205224451777446475056385919446288960817341194377871264566761375137792;
data[194]<=640'd129673105458552135625387182300070899538679260082920964054434413927371217374579518640156866201069314041957759265932172476180678963113397615963394304272314908897926704856668670263296;
data[195]<=640'd194509042756453700514867839363076163808046041629287269111461644297966826107200244185345543060660516166588439609025937322518244865331433015495196292435458122556102973501287010664448;
data[196]<=640'd64837668633355651170148328694101729285626640811311540862405271382245496814670216242611762186915391177011560132042557209500761061756766186768247684504019965600396468926024786116608;
data[197]<=640'd32419585973000014866643748945235205495340055437938319553226314951755362028053907603200602235231422497624852532736065106953109657695072046840058687799809232068636314202722818588672;
data[198]<=640'd48630115176541931636609535995837358272528785448065315728205359201205682357951212540414670610276427953754333253671761911778987584006834433019330688658616492805230196318945262174208;
data[199]<=640'd24319515400235089872593118426672851641454881573212056204369558432237103910727472201215717142198247277768704144363404044204629350805239937524725928408712908002315865453377754234880;
data[200]<=640'd12186469549530986918122912984234949280735066172653492679218876874729662066482704687516802234203313795560214392520320266504610578355988207685589006691245515255443801404170792075264;
data[201]<=640'd4044354393579852578329364978552179419616854163686935892481709553682257524050307072815481229162951832672516767421953972989306735926286224600631143020662415231768963145192106360832;
data[202]<=640'd981408723780445111202599807622412332803864324014315327344314119117038699262343200614501213995785282109851418796264054692912148754751202372611932092669100931323692651604929937408;
data[203]<=640'd93536104833244358554723857261783579261867076354048;
data[204]<=640'd144115188075855872;
data[205]<=640'd0;
data[206]<=640'd288230376151711744;
data[207]<=640'd0;
data[208]<=640'd0;
data[209]<=640'd0;
data[210]<=640'd0;
data[211]<=640'd1859015392949051632321347814954666316631744243705237457551454034012587162912871030435312937044214054582604819112781738467628392088522652910089393092722167001407708882622540743322894336;
data[212]<=640'd8465133328356180339480442389377213774379722311148627005162018011484832773364218454943728286662653879289748041687118174195144370759851084167453451901823286939147573264429270591682379776;
data[213]<=640'd12797300522971284902484470585366208237565080853459484514579955750524587648366844440438546201667343755455335074561489162968124662980811275749746206292275377271602502292103436376299536384;
data[214]<=640'd25519715257160401765358663452360603843460079024977014216124200290475272415746220326051723229441459816489499439594202299664598134650333979302558104684083524810787702757369616727329996800;
data[215]<=640'd17004844473635842335957438170464147107966845281077600367717159226024490618379904605761818065653789075176694212005218549421679825101275912947077366754458684292563069430501634515541164032;
data[216]<=640'd50997935358631987940188565593772267713078162105228267687866613382992995739068861202203205800170170465846029133834140279234809771644146499965170219844331089399642780572716679537778229248;
data[217]<=640'd34001389916133913251091789471347531289745213199018488569331276096288528990621232781170430736837553727447999084090295643594057283384640109842617058023561033491921930436898619878522486784;
data[218]<=640'd34001519588495440782121742984093271638531182337963246145484400960580081823521589434550005727682833324441570590274252246743719232840936125915000311223624887794254859209056008444628172800;
data[219]<=640'd50997935358631991714150990415313619954632743093497158604787833799433424115275161447827368192319022551972754311492907820703184802407991583885162209171801736537401944331619775341970587648;
data[220]<=640'd17004844473635840448976225759693470987189554786943154909256549017804276430276754482949736869579363032113331623175834778687492322668964727160093654407397515787906213658760218212634198016;
data[221]<=640'd25519715257160409313283513095443308326569241001514796049966641123356129168158820817300048013739163988742949794911737382601348196574198205775495040495507255866396204685086765675551129600;
data[222]<=640'd12863595517802246463435478441250018279055546103773468073628703868902258597293084217618747447763093976798943144085605147637921615528502290407736724638128837206036857843138311213818052608;
data[223]<=640'd8465076596697974305030589512137429956240050930171386396382821718952994646907309962848540306679323194337808731143961745633416963201267843134534843282475533433011152068713814441135702016;
data[224]<=640'd531146097092032167905855767038574878109068998875947922607802602304562555824227308468854072022742859419744503633146117286184324418034818358895216398861863818084469003003434454671687680;
data[225]<=640'd42535376994755722540756460814769061888;
data[226]<=640'd36893488147419103232;
data[227]<=640'd85070591730234618227026893292764659712;
data[228]<=640'd1190988284223284623154828794138923630592;
data[229]<=640'd0;
data[230]<=640'd0;
data[231]<=640'd0;
data[232]<=640'd15195979866507542572677274891447123355758470088778455444320034166347605510545317918944239681202772684160880932414431601009747867707806794340406035769460316236796320080816074915840;
data[233]<=640'd64582914432657055933878418288650274261973497877308435638360145206977323419817601155513018645111783907683743962761334304291428461703421701976239063869378643267744286249224264220672;
data[234]<=640'd227306532169841990982964236917896553529887115077977729354620511071616265761907047204207585231324808067239843947365872698437478545074519547246682483410783475237081783803481629392896;
data[235]<=640'd129862311275862374235671211676491875011085925633685883817918291979912245425535196048977648275612028230058194968258330056962470319452965652509315367189946898296160114694278411714560;
data[236]<=640'd129862311275862374235671211676491875011085925633685883817918291979912245425535196048977648275612028230058194968258330056962470319452965563300890055196719316569048428619334280019968;
data[237]<=640'd389080401165370204621257725866427387588065827898098369605610874800858482759587410882968136837462658934035888873694509117520425540711437657630489807270268758607097354610365473751040;
data[238]<=640'd389080401165370204621257725866427387588065827898098369605610874800858482759587410882968136837462658934035888873694509117523561026611479142775002645383652023467324703330012527329280;
data[239]<=640'd129767336401696702094591978708420330490112435195631018471391291766372572891094287811984246777604510900782189462430739859462436545092736508380746261521080821979691989644804502847488;
data[240]<=640'd194540200582685102310628862933213693794032913949049184802805437400429241379793705441484068418731329467017944436847254558766541952959544136136904537655658639775952159863904208420864;
data[241]<=640'd97285929437036829845494303627952104317178705380867069959157218735804566112303670760240934459033584288388306469394892312304247549735808973184426491855694559084785131036529121034240;
data[242]<=640'd113510803773672487279863269006840959983483321881906566657519755215498624079292161246613690368651128039705913714941551052962681144575566324525400757828811138094414921987842434400256;
data[243]<=640'd24329396932106346806463511987660654789375800548388006268666554701746114239279326709809683739592355849536743742834355594533756482301672638724688328028427136392501631657563310260224;
data[244]<=640'd14190829114920845746255392646023277175455696286031130526909281906386071187712372410764073827289880949323155995739102010736242286389037322735319600184034048691096661718714980237312;
data[245]<=640'd3053046475784002368442843119466524913793661373305358951899194364410723346715029368350385654699984147351593656082743224008134722863041122771150017187089895292762181863318667395072;
data[246]<=640'd763756219365548004034170149043797227016183351353802634991579863195565827198983807547555413099090920085337328700043837793972598564996931255460420169010629801502688605502154211328;
data[247]<=640'd190444401586365641583504236702019174350513356974090675900947696439118262840781212936845924644903694286672671915095677254881268218421752227168582967136255505302726712426433085440;
data[248]<=640'd16193216071664837027760010521889222892898001924772990125768619407147611223894223544119997374884591717802550116394407300041359485824525707628468730294761189249864950891665397121024;
data[249]<=640'd60783919469804132715530640918030048004022149246030742997696577093766628342426895838169107576897217461821182497199194779069755315730997761991548935710402700407543795981542869696512;
data[250]<=640'd97254271151309216102366871333623921348336611904557496674272879307188984717858470924831357237826935266396126118764564809008532120679619360723485817873388177710497131811955321864192;
data[251]<=640'd194508542293183526142679889286643956244202551581822690297504657543437453685102881443682342345438553719848105318675458680440154629109812259872159654165372764956709245056270456586240;
data[252]<=640'd129672361529418011165923516416469563259633079203034613735072511767021003506776191656186919705640056934095013340373883849465230393556503270686427234882342082346378279378121870278656;
data[253]<=640'd389017084584480071072949007897167135197910968718186919984801094872686804220082950806168610264834044077107381253580183173364927335769739227429356912014464812787702142090716215508992;
data[254]<=640'd389017084584480071072949007897167135197910968718186919984801094872686804220082950806168610264834044077107381253580183173364927335769739227429356912014464812787702142090716215508992;
data[255]<=640'd129672361529418011165923516416469563259633079203034613735072511767021003506776191656186919705640056934095013340373883849465233458594353054861465737718248085855282620415921642012672;
data[256]<=640'd194508542295070507355090659962764733534696686027281150907712877757625556835225693524878416771481617082436934702446192867955536551606466318208279555779479510951290826650374513885184;
data[257]<=640'd64836180775087402251220996926899056727534279051538840223681467061545069079063562274671869196056876961286068280925979956067215770252621456702075409096023099586573230752386290548736;
data[258]<=640'd113463316389425125156825231454186951856832341135716031070086421105995676015510445401607073548853143527555133707608313204636811240815078915896701089536531281795843931407305706307584;
data[259]<=640'd32418090351691058089805855617154759844378585062058668517884549461198574687198351594610520503210234591455275848819040415241351361571645170831657375541325202876969522033633020346368;
data[260]<=640'd13469200516990017663830868635516060651055665096163328;
data[261]<=640'd6681706001460045199136663066773394254253884949852955082752;
data[262]<=640'd6289363202875178113486973655552699949053063789152615530496;
data[263]<=640'd7858686614890462707953169810936694490535412800739380035584;
data[264]<=640'd12360329298116717340094278156246619881087592628421132288;
data[265]<=640'd24313567892083016011286797689078925636885081087719322882572386660689945223749985217290951348335984599631854983024205062486412447027281160549569285212755734140094488237794511552512;
data[266]<=640'd127646231357956585562824860822833267973881297892188020725176221401098086419774939142934517537041384644514063310047709077395167564728411554803646070429651385973149160673790570528768;
data[267]<=640'd67875376989922505954335098448647974581935182087977489419197661310891793396892572251558243665809541909488405590062842278244339246677211220748791533983298654975451814408469279145984;
data[268]<=640'd197547738994859782647772825247553415046090141546544176926741667053314790734617408369155918734301566215968423640661741381579526268400635411600289038088419894081369680778938002964480;
data[269]<=640'd195521608100684552691349000699659417501084867625107170207097034653348367150579128757807011391209626054865819626144372791111909967460967545458560180184533703555880759982114130100224;
data[270]<=640'd195521608100684552691349000699659417501084867625107170207097034653348367150579128757807011391209626054865819626144372791111909967460967545458560180184533703555880759982114130100224;
data[271]<=640'd195521608100684552691349000699659417501084867625107170207097034653348367150579128757807011391209626054865819626144372791111910021337763904024965356845171376808937996578411394367488;
data[272]<=640'd195521608100684552691349000699659417501084867625107170207097034653348367150579128757807011391209626054865819626144372791111909967460967545458560180184533703555880759982114130100224;
data[273]<=640'd195521609066818933445663586873497390234081703699839002633705784317657180013458914330197117525258067700346464116760276798987454261802237210719307094120260871922650947156359333806080;
data[274]<=640'd16535252224444826591873994903048945965403480550973523278996372648091587099828621631375997973398105005108701423484378336291713484076563448775328036537655972323224915251452911145713664;
data[275]<=640'd132721688146350632255547418368522652773266244268461362882193620741886798180924952637601662638191693685341172151858374472437406595088929212385492784693455005740933472610486373731794944;
data[276]<=640'd232372871857337492657907251137381145233987483140021924860367018682890745542272979010464790815463855543501670479616614928401643842145509302533979953106698247192551897338506358024044544;
data[277]<=640'd398353494612577210998403565685027591274485332429719400860193311870516857998789304866453072773348007315029585944068646495697449885161980314849454946471256794674999169474566738971459584;
data[278]<=640'd265568996408385436326006514046910434442087052997961420060332277320415968033576244181662447207040685897807253572507021241860805050748803504997074951779609956689041351765718434213527552;
data[279]<=640'd265568996408389210288431335588262675996668041266852336981552693760844344239876489805824839355892772024532431231274562710235835814593703275581704876572242518123292784461762083608854528;
data[280]<=640'd796706989225156308978019542140731303326261158993884260180996831961247904100728732544987341621122057693421760717521063725582415152246410514991224855338829870067124055297155302640582656;
data[281]<=640'd796706989225154421996807131370055182548970664859438801720386623741033715997578609732906145546696014630059171888137292991394899770323960629698909892942513589349998338949133477942919168;
data[282]<=640'd796706989225161969921656774452759665658132641397220635562827456621890468410179100981230929844400186883509527205672375928144961298013760170868169742527778712218501204341220776733573120;
data[283]<=640'd265568996408406193119343032524347762992282488476861463127044567742772037168227595114555604025727159594795730695728499317923474251895752243212539538139089044577424231593958505887825920;
data[284]<=640'd398353494612620611566289013410578369152166697521964945454228100935443184371242129544320582485146997772369129019895373382010303669378327676572699081586531251168890645479068707017719808;
data[285]<=640'd199176747306740537499574162419444721798316011414547001746241524676556479703849065926672996211711317332854817609447414085758658913007737684934160967153377629089108650088510384576135168;
data[286]<=640'd124487493196957889630120970224115297733562530158775602648208969801567058754847457127850521937103851476464806301902018611684338055607921641434360705797279539424621180671325947203420160;
data[287]<=640'd33133314497068508302448271828615955873963780837273616921088967497647083803741492048176459776358331793962462207073963046810152073572736855718778332735988364849243615555514388931674112;
data[288]<=640'd195521607615730381101780936936619653844092315142282793383584439607005857569016423890415883898142341869536667997065686599658755897840447420513224326900389402246779318373166830583808;
data[289]<=640'd195521607615730381101780936936619653844092315142282793383584439607005857569016423890415883898142341869536667997065686599658755897840447420513224326900389402246779318373166830583808;
data[290]<=640'd195521607615730381101780936936619653844092315142282793383584439607005857569016423890415883898142341869536667997065686599658755897840447420513224326900389402246779318373166830583808;
data[291]<=640'd65849246088199351148268191196270867874953370384706640258720148054172957212363044315425038618545348298030484040462536937708907426733829442141759488334328037026117387016869657968640;
data[292]<=640'd65849246088199351148268191196270867874953370384706640258720148054172957212363044315425038618545348298030484040462536937708907426733829442141759488334328037026117387016869657968640;
data[293]<=640'd128659296203097193782000927414252311078755046751657589428576289275076393322617025047061229300850142059228791894442187555215865279926097525415437769514764010804875510017576100954112;
data[294]<=640'd62810050114897842633732736217981443203801676366950949169856141220903436110253980731636190682304793761198307853979650617506957853192268083273678281180435973778758123000706442985472;
data[295]<=640'd0;
data[296]<=640'd0;
data[297]<=640'd0;
data[298]<=640'd0;
data[299]<=640'd31163630585611171291623317648475545944426549986752691829171945067705050363423015263459866533716623668689306599678033556758271994322650652455910815542838539157492453290736091136;
data[300]<=640'd126509500353492969171947039501549537702969685065269856116043253191516930641991050057616839142825817512179208934407255272078223215047903243898399858334618355389344363954059608064;
data[301]<=640'd475246272181552319367180132112351512837038707359071450340574972572014076991999956883487465309592553585616135597500019123886423858360733631902871751772508065998810388538603864064;
data[302]<=640'd886619211553230504948423535745667631645220161462111954705394031326009028897795016404118778188501778721872479729381868171443904512211993928945725694812423123959826110010923941888;
data[303]<=640'd1519786405498775897541279500998722755888494927086696055636830527110506614086463382318013220083158488207716368591534946016695252716988913059237576839112468652462307247792702095360;
data[304]<=640'd3039260711852943903255811329916706943916248806622306112483115198712395515545945258710256621658398234390674592831391597924944984206170100597974026112735212323827196777890653929472;
data[305]<=640'd6078456688928414842612807660447686196056211715294918421763562460358122917900633004891253409985079496400509546855746293157658402647502044095980025899188709822619156837703264239616;
data[306]<=640'd12156848627983507022040634912543426376383061968972458158658695270144752521627511847684651578293935119709544384738582183500029859931083592572292854941849967814472292782730903552000;
data[307]<=640'd8104585397979400827364189260481581348853797795834538520289186830501098659722522591185975395209645779638687154862925740813008506526462450226690750865206213417786233079356209496064;
data[308]<=640'd16209107995337071411869506545374157762419116288641508700801425266741258082136170895818977651227521240446653035921356782200255958420511366189869699591865765869793951810949480448000;
data[309]<=640'd48627198856513056852583444715138786040214001624484541974905432558727683302493784413369593186064863730885862502838627826594726378468030108783184573568683257106911832193496980127744;
data[310]<=640'd32447832347614069898167025626279572723879013216947835828478334017045905562045110218166069360194147054365696738218452047696173189042550006371200660350810645267708896412372473741312;
data[311]<=640'd32669440628867566749263882428572669789399699924425479743693521931382344691460509164248199389057131234046537374470138510513118085698606271770518310189713733637854722873779009093632;
data[312]<=640'd97731186235709362683926140510997994644782794056227945290822918382801110707644463228407897519599260854089820183804288056627758618992568185429367674598333758633940540341004607160320;
data[313]<=640'd65724653641877851140224630270887491076716516431738323511223846419931466601058387361631592691065920888075964719906391497000977172633000124849887461758907967560188291170785749368832;
data[314]<=640'd66611085799813967184092085968161517960555359964187836440371738305874358680778791532971969459447884280024268082411866246635521503691012875028929949020652794111143235831254338240512;
data[315]<=640'd196030180875469740500437553855256438615473725710942869587837935581229530671063109279431647477602109767776023462147787380917431140209842032003794656081923924682012288456090592477184;
data[316]<=640'd195523648213252822414681644692208201170281776707983587739693934442351277154044932015466839488228684011637327431067306327550439544619581805525781121556275247474119077786730056646656;
data[317]<=640'd132713598098354979780948908474226757966480100341032638569837793221447841043790951283830648805923890250439019577087655710043481691427313722252102840375839273695360954786023613661184;
data[318]<=640'd132713598098354979780948908474226757966480100341032638569837793221447841043790951283830648805923890250439019577087655710043481691427313722252102840375839273695360954786023613661184;
data[319]<=640'd132713598098354979780948908474226757966480100341032638569837793221447841043790951283830648805923890250439019577087655710043481691427313722252102840375839273695360954786023613661184;
data[320]<=640'd132713598098354979780948908474226757966480100341032638569837793221447841043790951283830648805923890250439019577087655710043481691427313722252102840375839273695360954786023613661184;
data[321]<=640'd130687467570254105032214595093763554777336908838536990230587882373973428583578215424520180115186242431569316014092719497559958345858931524497642066515210460909634385505362120802304;
data[322]<=640'd131194000232471023117970504256811792222528857841496272078731883512851682100596392688484988104559668187708012045173200550926949941449191750975655601040859138117527596174722656632832;
data[323]<=640'd131194000715538213495127797343730778589027275878862188292036258345006088532036285474680041171583889010448334290481152554864722088619826583606029058008722722300912689761845258485760;
data[324]<=640'd65598020717857216807364299523584924898667738199681461155840033551289106437523789438737917227234674860411451834790247235628115347320752484545570806611427590349907535297006916337664;
data[325]<=640'd65218123636530480128833833085893678647265866634291580836253906857902448456959620421739576570325709657009041038019646465291732386481231477838927940556509003360913095230599523729408;
data[326]<=640'd65079660155483914025287157149155503739710144292263696550078267111769379114730742188898763149814404307482579438504949765910100278736615303373463413945920182957997843930740011565056;
data[327]<=640'd97315725023226274119742675467151967230097384556037567183205086233781360475013535352310182939016994274053226447645229381599242735260716681683262648974552214559278575927964899213312;
data[328]<=640'd32424026315292074422017179847833222605833848232689388585790450829930660922811525820951947765610844951133955100806480177862370395437248441251830223381799220992628177445255257260032;
data[329]<=640'd48627135576598098657388821004872349319415373175007978642240549760688543933990641503013715831934999314492477751267649498261957021564752326519224107094834446209180920302260835057664;
data[330]<=640'd16209045198489303593832175922026707408118905876530861581440917300856525145072920771658153364121877646793590529658330457805258748687868416556282690085880539155448133506835937230848;
data[331]<=640'd24313567793959992965926722530798506531190089923879371151744935522908581417363756995095081194096689745012727026946027311677124278132032040204499242496259374481739504216604510519296;
data[332]<=640'd8104522610566539071380712017738017447024259611016194451969779935556881473273332873005523238319318998929771567453570353994920909043245962167915722940624572332022154884366154596352;
data[333]<=640'd12156783938493583156000316140056353656466002762025819000453312473592560011383744283861177969995738849460609956429165781176964432963492451031422340206305464006629408588445603856384;
data[334]<=640'd6078392037178115224787902410376159286021841417517491467722583947567993410113107064989268322548150477928162793961013641142231424677616748854357437489258548529103233079911917813760;
data[335]<=640'd3039196154451704905969439885884044558588600781767909668853147395327423513899023378611992836374637345359797028473368321678614128730549421104471253516840907316128674111334190678016;
data[336]<=640'd1772864680059606083013651885858070833045635038381923628482285110189692133143540013523117763075155763540677792762647689737799694943886917145827463565668058365165057533103826796544;
data[337]<=640'd379901187397854884367457676502630366638424883000168132673312766699112647803257699656291726614842196695149881888192803807446211789917084064817250281759052547767735556949508358144;
data[338]<=640'd237443948354845632900185637044670433411578618259990352578748184010871376260769599214246683357884841554525198880303548894587370821822137986797241858987996008591252720979177111552;
data[339]<=640'd63308853702068726202799254677247816674305027515250818148002827889278786588987578874751926284145055672181078957828068666519594718625206223776380329888737716825153939708437331968;
data[340]<=640'd3833621222833120277937789075804531445544535911068783518667977369439906989151243941139904216449267197338763907103250159759946158031754643754496965404079344102707404968304836608;
data[341]<=640'd0;
data[342]<=640'd0;
data[343]<=640'd0;
data[344]<=640'd0;
data[345]<=640'd0;
data[346]<=640'd24897093413285957751074447182146966906074677393454621399973943978143916868477448878398242293682622765729187319667804735094370906452470651847321249004683782122367090820409057142112256;
data[347]<=640'd264531617516163301105166001310311523377043447305455352374723154767779116727572894332981324370377866885872615271470425310377690881057500675877788270674765185050150339966846232134942720;
data[348]<=640'd399909562950905696376633307863235655928824505632364856237081475148936664699919022609271766842277128174525071322164113557453332684892809845297597562137733250340521396302820480345178112;
data[349]<=640'd797225678671260772154196360811664336138266232369578189411665664466816671392704977627043716778962316477620018965196164121667668400363487331027765827504145273376629553978515017238052864;
data[350]<=640'd797485023394315834214103386303145033710204510259093341717915393049922337193418284386193698469521510464763031333109370420991568097305700566984508757181277396107070877841227611583283200;
data[351]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[352]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[353]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[354]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[355]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[356]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[357]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[358]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[359]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[360]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[361]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[362]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[363]<=640'd531656682262862126959702971370021056255145720430498560127061929604901386637077873760812897050939329136274643587002747740494255676157534628984486138950321351667708187776643810140880896;
data[364]<=640'd531137992816793516426561957341934318211660035609268341647987053283402193304953962108299247307193888555965573097619291293971794684567005633501929452315015281983591299707698764799016960;
data[365]<=640'd531137992816772759633225438864496989661464600130368298581274762861046124170302611175406090488507414858977095974397813217909125483420056895286464865955536194095208419879458693124718592;
data[366]<=640'd531137992816769929161406822708482808495528858928700110890359450530724842015577426957284296376868350263933212730322157116627852410536382067347992422361061773019519845357425956078223360;
data[367]<=640'd531137992816768042180194411937806687718238364794254652429749242310510653912427304145203100302442307200570623900938386382440337028613932182055677459964745492302394129009404131380559872;
data[368]<=640'd531137992816768042180194411937806687718238364794254652429749242310510653912427304145203100302442307200570623900938386382440337028613932182055677459964745492302394129009404131380559872;
data[369]<=640'd531137992816767570434891309245137657523915741260643287814596690255457106886639773442182801283835796434729976693592443698893458183133319710732598719365666422123112699922398675206144000;
data[370]<=640'd531137992816767570434891309245137657523915741260643287814596690255457106886639773442182801283835796434729976693592443698893458183133319710732598719365666422123112699922398675206144000;
data[371]<=640'd531137992816767570434891309245137657523915741260643287814596690255457106886639773442182801283835796434729976693592443698893458183133319710732598719365666422123112699922398675206144000;
data[372]<=640'd531137992816768042180194411937806687718238364794254652429749242310510653912427304145203100302442307200570623900938386382440337028613932182055677459964745492302394129009404131380559872;
data[373]<=640'd531137992816768042180194411937806687718238364794254652429749242310510653912427304145203100302442307200570623900938386382440337028613932182055677459964745492302394129009404131380559872;
data[374]<=640'd531137992816768042180194411937806687718238364794254652429749242310510653912427304145203100302442307200570623900938386382440337028613932182055677459964745492302394129009404131380559872;
data[375]<=640'd531137992816768985670800617323144748106883611861477381660054346420617747964002365551243698339655328732251918315630271749534094719575157124701834941162903632660956987183415043729391616;
data[376]<=640'd531137992816772759633225438864496989661464600130368298581274762861046124170302611175406090488507414858977095974397813217909125483420056895286464865955536194095208419879458693124718592;
data[377]<=640'd531154201861950492143482752562981687818677283557344786376143913355990911560796333163284591823185063039635412441705993472304261541021796025487556562286142986745980988184725457387651072;
data[378]<=640'd531656674348304375670057167599349349844759592381859056573164718116597096489567652848442716196222839683397914554947427981477919872293452613506967119159374634144132545229401698963816448;
data[379]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[380]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[381]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[382]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[383]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[384]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[385]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[386]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[387]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[388]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[389]<=640'd531397337539822160749495232043949324901531395616547075505693866783509225661565549498312483955788479656032341854159707314670479034594920475366262908443719474674272594698105813376958464;
data[390]<=640'd796966333948205710094289335320183638566327954480063037105415935883711005591991670867893735088403122490477006597282957822343768703421274095071022897827013150646188230115802422892822528;
data[391]<=640'd796966333948205710094289335320183638566327954480063037105415935883711005591991670867893735088403122490477006597282957822343768703421274095071022897827013150646188230115802422892822528;
data[392]<=640'd399131528781740510196912231388793563213009671963819399318332289399619667297779102331821821770599546213096034218424494659481633594066170137427368773106336882149197424714682697309487104;
data[393]<=640'd466301812053001583712831833682294234345023645348243846637011992423987109682525552951667079625430788883136237507944926184371655102099398250223787559483556669333500305157244632724144128;
data[394]<=640'd131747119311971526432768949672194366544645167873697371574862120217678226762359833648190698804070545468650282899908800056541046046644323866025408275983118347064192522257997927377010688;
data[395]<=640'd0;
data[396]<=640'd0;
data[397]<=640'd0;
data[398]<=640'd0;
data[399]<=640'd0;
data[400]<=640'd0;
data[401]<=640'd0;
data[402]<=640'd0;
data[403]<=640'd0;
data[404]<=640'd0;
data[405]<=640'd0;
data[406]<=640'd0;
data[407]<=640'd0;
data[408]<=640'd0;
data[409]<=640'd0;
data[410]<=640'd0;
data[411]<=640'd0;
data[412]<=640'd0;
data[413]<=640'd0;
data[414]<=640'd0;
data[415]<=640'd0;
data[416]<=640'd0;
data[417]<=640'd0;
data[418]<=640'd0;
data[419]<=640'd0;
data[420]<=640'd0;
data[421]<=640'd0;
data[422]<=640'd0;
data[423]<=640'd0;
data[424]<=640'd0;
data[425]<=640'd0;
data[426]<=640'd0;
data[427]<=640'd0;
data[428]<=640'd0;
data[429]<=640'd0;
data[430]<=640'd0;
data[431]<=640'd0;
data[432]<=640'd0;
data[433]<=640'd0;
data[434]<=640'd0;
data[435]<=640'd0;
data[436]<=640'd0;
data[437]<=640'd0;
data[438]<=640'd0;
data[439]<=640'd0;
data[440]<=640'd0;
data[441]<=640'd0;
data[442]<=640'd0;
data[443]<=640'd0;
data[444]<=640'd0;
data[445]<=640'd0;
data[446]<=640'd0;
data[447]<=640'd0;
data[448]<=640'd0;
data[449]<=640'd0;
data[450]<=640'd0;
data[451]<=640'd0;
data[452]<=640'd0;
data[453]<=640'd0;
data[454]<=640'd0;
data[455]<=640'd0;
data[456]<=640'd0;
data[457]<=640'd0;
data[458]<=640'd0;
data[459]<=640'd0;
data[460]<=640'd0;
data[461]<=640'd0;
data[462]<=640'd0;
data[463]<=640'd0;
data[464]<=640'd0;
data[465]<=640'd0;
data[466]<=640'd0;
data[467]<=640'd0;
data[468]<=640'd0;
data[469]<=640'd0;
data[470]<=640'd0;
data[471]<=640'd0;
data[472]<=640'd0;
data[473]<=640'd0;
data[474]<=640'd0;
data[475]<=640'd0;
data[476]<=640'd0;
data[477]<=640'd0;
data[478]<=640'd0;
data[479]<=640'd0;
end


// stuff for drawing game area:
always @(posedge pxl_clk) begin
	if(HorizontalCounter>=144 && HorizontalCounter<784 && VerticalCounter>=35 && VerticalCounter<515
		&& data[VerticalCounter-35][HorizontalCounter-144]==1'b1)begin
			if(HorizontalCounter<444) RGB <= `YELLOW;
			else RGB <= `WHITE;
	end
	else begin
	// Draw top margin
	if (VerticalCounter < TMARGIN_END)
		RGB <= `BLACK;
	
	// Draw top border
	else if (VerticalCounter < TBORDER_END) begin
		if (HorizontalCounter >= LMARGIN_END && HorizontalCounter < RBORDER_END)
			RGB <= `WHITE;
		else
			RGB <= `BLACK;
	end
	
	// Draw game
	else if (VerticalCounter < BGAME_END) begin
		if (HorizontalCounter < LMARGIN_END)
			RGB <= `BLACK;
		else if (HorizontalCounter < LBORDER_END)
			RGB <= `WHITE;
		else if (HorizontalCounter < RGAME_END) begin
			// draw game board
			case (ShiftedHorizontalCounter)
				SHIFTED_HGAME_START:     RGB <= (a[9] & b[9]) ? `RED : (a[9]) ? `BLUE : (b[9]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 1: RGB <= (a[8] & b[8]) ? `RED : (a[8]) ? `BLUE : (b[8]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 2: RGB <= (a[7] & b[7]) ? `RED : (a[7]) ? `BLUE : (b[7]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 3: RGB <= (a[6] & b[6]) ? `RED : (a[6]) ? `BLUE : (b[6]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 4: RGB <= (a[5] & b[5]) ? `RED : (a[5]) ? `BLUE : (b[5]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 5: RGB <= (a[4] & b[4]) ? `RED : (a[4]) ? `BLUE : (b[4]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 6: RGB <= (a[3] & b[3]) ? `RED : (a[3]) ? `BLUE : (b[3]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 7: RGB <= (a[2] & b[2]) ? `RED : (a[2]) ? `BLUE : (b[2]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 8: RGB <= (a[1] & b[1]) ? `RED : (a[1]) ? `BLUE : (b[1]) ? `GREEN : `BLACK;
				SHIFTED_HGAME_START + 9: RGB <= (a[0] & b[0]) ? `RED : (a[0]) ? `BLUE : (b[0]) ? `GREEN : `BLACK;
				default:		         RGB <= `BLACK;
			endcase
		end
		else if (HorizontalCounter < RBORDER_END)
			RGB <= `WHITE;
		else
			RGB <= `BLACK;
	end
	
	// Draw bottom border
	else if (VerticalCounter < BBORDER_END) begin
		if (HorizontalCounter >= LMARGIN_END && HorizontalCounter < RBORDER_END)
			RGB <= `WHITE;
		else
			RGB <= `BLACK;
	end
	
	// Draw bottom margin
	else
		RGB <= `BLACK;
end
end

always @(negedge HSync) begin
	if (VerticalCounter == 0) begin
		// load new grid
		GridA_Buff <= GridA;
		GridB_Buff <= GridB;
	end
	else if (VerticalCounter > TBORDER_END 
			&& VerticalCounter[3:0] == TBORDER_END % 16) begin // is 16 lines after TBORDER_END
		// shift grids by 10 (move to next row)
		GridA_Buff <= GridA_Buff << 10;
		GridB_Buff <= GridB_Buff << 10;
	end
end

endmodule
