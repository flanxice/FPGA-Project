`timescale 1ns / 1ps


// VGA Driver
module vga_driver(
    input vga_clk,      // VGA驱动时钟
    input sys_rst_n,    // 复位信号
    //VGA
    output vga_hs,      // 行同步
    output vga_vs,      // 场同步
    output [11:0] vga_rgb, //4+4+4
    
    input [11:0] pixel_data,    //像素点RGB data
    output [9:0] pixel_x,       //像素点横坐标
    output [9:0] pixel_y        //像素点纵坐标
);

// some parameters for sure in the reference Table 
parameter H_SYNC = 10'd96;
parameter H_BACK = 10'd48;
parameter H_DISP = 10'd640;
parameter H_FRONT = 10'd16;
parameter H_TOTAL = 10'd800;

parameter V_SYNC = 10'd2;
parameter V_BACK = 10'd33;
parameter V_DISP = 10'd480;
parameter V_FRONT = 10'd10;
parameter V_TOTAL = 10'd525;

// counters for H and V
reg [9:0] cnt_h;
reg [9:0] cnt_v;

wire vga_en; // 使能控制rgb数据输出
wire data_req;

//*******************************Main Code************************************
//VGA 行场同步信号
assign vga_hs = (cnt_h <= H_SYNC - 1'b1) ? 1'b0 : 1'b1;
assign vga_vs = (cnt_v <= V_SYNC - 1'b1) ? 1'b0 : 1'b1;

// 使能使RGB输出 // 范围内输出
assign vga_en = (((cnt_h >= H_SYNC + H_BACK) && (cnt_h < H_SYNC + H_BACK +H_DISP))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;

//在范围内RGB赋值
assign vga_rgb = vga_en ? pixel_data : 12'b0;

// 请求像素点颜色数据输入
assign data_req = (((cnt_h >= H_SYNC + H_BACK -1'b1) && (cnt_h < H_SYNC + H_BACK +H_DISP -1'b1))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;
// 像素点坐标
assign pixel_x = data_req ? (cnt_h - (H_SYNC + H_BACK -1'b1)) : 10'd0;
assign pixel_y = data_req ? (cnt_v - (V_SYNC + V_BACK -1'b1)) : 10'd0;

// H counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_h <= 10'd0;
    else begin
        if(cnt_h < H_TOTAL - 1'b1)  cnt_h <= cnt_h + 1'b1;
        else cnt_h <= 10'd0;
    end
end
// V counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_v <= 10'd0;
    else if(cnt_h == H_TOTAL - 1'b1) begin
        if(cnt_v < V_TOTAL - 1'b1)  cnt_v <= cnt_v + 1'b1;
        else cnt_v <= 10'd0;
    end
end
endmodule 


module vga_display(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    output reg [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;

// some frequently-used colors define
localparam WHITE = 12'b1111_1111_1111;
localparam BLACK = 12'b0000_0000_0000;
localparam RED = 12'b1111_0000_0000;
localparam GREEN = 12'b0000_1111_0000;
localparam BLUE = 12'b0000_00000_1111;

reg [0:639] data [479:0];
always @(posedge vga_clk) begin
    data[0]<=640'd0;
    data[1]<=640'd0;
    data[2]<=640'd0;
    data[3]<=640'd0;
    data[4]<=640'd0;
    data[5]<=640'd0;
    data[6]<=640'd0;
    data[7]<=640'd0;
    data[8]<=640'd0;
    data[9]<=640'd0;
    data[10]<=640'd0;
    data[11]<=640'd0;
    data[12]<=640'd0;
    data[13]<=640'd0;
    data[14]<=640'd0;
    data[15]<=640'd0;
    data[16]<=640'd0;
    data[17]<=640'd0;
    data[18]<=640'd0;
    data[19]<=640'd0;
    data[20]<=640'd0;
    data[21]<=640'd0;
    data[22]<=640'd0;
    data[23]<=640'd0;
    data[24]<=640'd0;
    data[25]<=640'd0;
    data[26]<=640'd0;
    data[27]<=640'd0;
    data[28]<=640'd0;
    data[29]<=640'd0;
    data[30]<=640'd0;
    data[31]<=640'd0;
    data[32]<=640'd0;
    data[33]<=640'd0;
    data[34]<=640'd0;
    data[35]<=640'd0;
    data[36]<=640'd0;
    data[37]<=640'd0;
    data[38]<=640'd0;
    data[39]<=640'd0;
    data[40]<=640'd0;
    data[41]<=640'd0;
    data[42]<=640'd0;
    data[43]<=640'd0;
    data[44]<=640'd0;
    data[45]<=640'd0;
    data[46]<=640'd0;
    data[47]<=640'd0;
    data[48]<=640'd0;
    data[49]<=640'd0;
    data[50]<=640'd0;
    data[51]<=640'd1560874275157996115690798615527015252016628656686887639465560760232206245291554929911303623195956733836676545678301012813445685112496363354980352;
    data[52]<=640'd13093574138141631181704007353419280485298290262935203042305711783195886614290246628086407957498762430697434539832898781346963605374783349011933294493696;
    data[53]<=640'd206223657464996605650950506530967900251416997185860835787625428998971656469301686322905969241617367928390027621641172541077128312433945847919444695711744;
    data[54]<=640'd417357383282006296454263527395298650038881148200462971092985776759271921083233894391555047973787675836783211610947451134870273424428901971012099403415552;
    data[55]<=640'd1563044213891670921046949369590907308477552891693234968333152183022115983139618976111748433997495092162708107186601385411900585343253590414381396776714240;
    data[56]<=640'd1674339594846312164874949793042181788187459685356403902341983168254552881218860880736088794059131335169369925855699137636858342001722734698470852328947712;
    data[57]<=640'd6702267866701781564524906989445949134072110749627488689492387126765454385639944315993077056392238363770953764833592173383292561635886201629182623989366784;
    data[58]<=640'd12568184387040289899858392861048392677154947848950001670488114716277554806386272708403614576630282811618577970783329328942322929554136226120957906114314240;
    data[59]<=640'd24745199255125922972992974388594524219876016766833408538195217781039731843551752613493750783513365950073799613291285466803702260311658345292683851295883264;
    data[60]<=640'd52816158465948640949110517055596563516136498956612759404175220668096999330883242151651716567952075059108864940029372847183510880302734226594067914847944704;
    data[61]<=640'd38565456853016490619685454491226599059741948021176906213338976448415625380495554357452988651939786204267013804906126511287835085925860523707452395616206848;
    data[62]<=640'd50287475608707131256170343317573522574427779602618137424396190362604982222026835727096262786674314065325967568588934395125005266952638020896081880778014720;
    data[63]<=640'd207843953441811946752441544746760321479754358068521398687276820751178032132921565041711216301683182447683285970276004039052215955467708879996397239610114048;
    data[64]<=640'd281586897854102976474440453302534394437777855996322629328997427200684478220781420769680459266168107343617739163804765483588229231919291975451710866774294528;
    data[65]<=640'd362033775809932917235589452156667120505681476750361562950688639123151573394305915527236354162842021508989410596782523303821220710488540845697132048383213568;
    data[66]<=640'd831333291635758742242014795100733225645314355755988439291240912841170845462366392790231749299997162597147550923970579194926065748256485384624996257946927104;
    data[67]<=640'd1662614157850088671263851545174688367346325975022342040070821065130160204636645381849399682226046017092721118579741678558832153867809550592830226768374792192;
    data[68]<=640'd1662607630248896115023875694367923919933316808886578781355046512484291412326468330638384108731937358612545379499486873218869053046002661958680472823879696384;
    data[69]<=640'd2788922583621883304436004494798184232638358306674113490421324597927091172945566041787178868067226860644007176807348826402058781315592732129841532325712625664;
    data[70]<=640'd6757608004080583052627868522301533693951437227890790728846686427712585575224167047449156286754665892558720147163065028636578963885093424234546202931051364352;
    data[71]<=640'd6650358557502112026778378789618056703783585209049149155279966860071348110749765125166233276502581179979198124760798074318796409144430456784216483650282192896;
    data[72]<=640'd13300638655863777844430170039640040645014385064310812338877137856313543148026826556497217936666519485202236706312657056789007947174795911584983861204415938560;
    data[73]<=640'd12442645333554695226299039783515406591292812514707948360298123032888027142801104970007169822328340076814882727496418981056308634028824299616499754320468639744;
    data[74]<=640'd26601291632861412376945179998197305586415064659739660342098020058780361420033041244505716050620043522473389315541707276512600208922248773768306228544296452096;
    data[75]<=640'd19736502360794236275900592615804755955703646396901316648241854682316007183478375555812799863684044951162022858617491467403795148225782617756701592852379992064;
    data[76]<=640'd49769876736821750398987454571902764606525705730396284443982756144262809655705736825827703011071307679152860468611761272414186828454972791344844881392633380864;
    data[77]<=640'd53202375814499397116083445032278691755521080221463037344070346709447112301717070635436893212990525491954036532080687106005215040926764947752838973010657411072;
    data[78]<=640'd51486399808325785427957717570429735135383491431818756877901466745020216625986047793217690684279782587407616394229991562656079969261958297759095201970891259904;
    data[79]<=640'd106404777816098683393547968021327994759242854796898843547402907044261812523807219539222329405842250358958849406241899713777065214211649217594803769800556281856;
    data[80]<=640'd212809562178841222451680895880945465005697826227023705321034451003222789112867805222381929892358062735528830627094321620598394527036980401357003916783160131584;
    data[81]<=640'd185350368264928178363121170205988136365190316771674930338992212948351368633541514245865703587643551529197154380029411349718121264404263388064821469627912552448;
    data[82]<=640'd418753377414088240394218627495780104425166249073415823978210337593900434035412352487465926462313536306611948115330941319723076520135949664451724649392569843712;
    data[83]<=640'd151026294856119323916913814378267157557491958587996507459317566722600079653267373174071591439196317358992647783631868512756553059486080597364562619431305347072;
    data[84]<=640'd755128344918626030171610897558341787850507578505111342691994470807135517582066470482910602790139719618601300162159359615939706788266180050393884815899012104192;
    data[85]<=640'd631562510778460143067461551222270237254183504562376425773411688871073900367353472597863287139797710451911027827131794377890056969079187240148350247530940858368;
    data[86]<=640'd741399666147722534286140224918785827770768974850875942870044782154784779378842814168434071218925052615733670678353074725606139016377228075921621804523859214336;
    data[87]<=640'd1675013928649976150262848114806491073731402845680113199794707089565412689469090753577207368972766196426486290438330309467659561457385042766659031614379784142848;
    data[88]<=640'd1647554580887079155171184979595546075145563219533269012114648043275482251384127149077579899249210327491074152636671161873332196497669170856091024537653465841664;
    data[89]<=640'd604105441295301372609018263991595790035404120759839646474821775833338234445399284314722197283191195566519875404403933823204435069955628398789629422197236826112;
    data[90]<=640'd1208207530638720128076557745979800702912230386522580170337042143877027515707330843279785459190360566083910040985715982147616393889310122910463016908173770489856;
    data[91]<=640'd3404942781879965798424541740254495352677622127437073917981332446479635152749142546759351264300749230091394093158971612639668431328567119932955346074430376771584;
    data[92]<=640'd3404941734394871386355569613016362811268948524023303489695002516646187321579694027453491549468005499153222254185675312047263206468076546518013531908956787572736;
    data[93]<=640'd3295105809820677348703244438945479736786752119570644348904123479267051022766805679198867059493496206216618867768362956386111758817487918583688680186966496509952;
    data[94]<=640'd2196737765205781978175647510906545622900039025763215802653288228673121063112443107697620397183617150899508435358418918883469977397074888039828110248756333510656;
    data[95]<=640'd1318041150745077065276524953955980078986928030671079363718134815020968012430342271532824840978910539806079010076181252043342268902095010193502455132878444429312;
    data[96]<=640'd0;
    data[97]<=640'd0;
    data[98]<=640'd0;
    data[99]<=640'd0;
    data[100]<=640'd0;
    data[101]<=640'd0;
    data[102]<=640'd0;
    data[103]<=640'd0;
    data[104]<=640'd0;
    data[105]<=640'd0;
    data[106]<=640'd0;
    data[107]<=640'd0;
    data[108]<=640'd0;
    data[109]<=640'd0;
    data[110]<=640'd0;
    data[111]<=640'd0;
    data[112]<=640'd0;
    data[113]<=640'd0;
    data[114]<=640'd0;
    data[115]<=640'd0;
    data[116]<=640'd0;
    data[117]<=640'd0;
    data[118]<=640'd0;
    data[119]<=640'd0;
    data[120]<=640'd0;
    data[121]<=640'd0;
    data[122]<=640'd0;
    data[123]<=640'd0;
    data[124]<=640'd0;
    data[125]<=640'd0;
    data[126]<=640'd0;
    data[127]<=640'd0;
    data[128]<=640'd0;
    data[129]<=640'd0;
    data[130]<=640'd0;
    data[131]<=640'd0;
    data[132]<=640'd0;
    data[133]<=640'd0;
    data[134]<=640'd0;
    data[135]<=640'd0;
    data[136]<=640'd0;
    data[137]<=640'd0;
    data[138]<=640'd0;
    data[139]<=640'd0;
    data[140]<=640'd0;
    data[141]<=640'd0;
    data[142]<=640'd0;
    data[143]<=640'd0;
    data[144]<=640'd0;
    data[145]<=640'd133499189745056885244540783077509605799792373029558743665569425777073550597423730724612834590720;
    data[146]<=640'd467247164107699090250446494159149940649304354995302053100594063624917944328952176982225846272000;
    data[147]<=640'd12608641982846233347929693329615191588380599801463792761525286286257585952358148115887717036126291614596243987330236416;
    data[148]<=640'd69347530905654283413611511073821995467906860705881375337859773964318495465209171570881070618079355551389817531443183616;
    data[149]<=640'd322150802661721262039593832356343421641802395037548481241899405372716856126112705826979870644120693708407580657444716544;
    data[150]<=640'd607106111474046135702795716861392291624088917448351038442872475653016367778894527258940068893681317757389778614866673664;
    data[151]<=640'd2421489692805619114469821489389564400348158492328928492559875100713188127784809157634669337313757959880538356552493432832;
    data[152]<=640'd4518937286652090031897859352000409250423957448354473526683029238359403486573994562124111969606202207115995234891244503040;
    data[153]<=640'd3873374817130362884483879025002897301621598951751997860267323887506997950551353740056231394726160724591157371294921523200;
    data[154]<=640'd18075749146608360127591435005016221590660604273478089534684741230367592942293524698581150340340558713054910993622928195584;
    data[155]<=640'd15493499268521451537935516634008348186687356479502519343809290875226192913492644585645909621024169132520734114127888252928;
    data[156]<=640'd30986998537042903075871031666026419432650414135767947994808815572584297080737998591448638589958999639843114061018616037376;
    data[157]<=640'd61976518860200157912661398632217220127121706099206988296209503185600154124273563513079016638792378406246342112377701400576;
    data[158]<=640'd82649652194515260118886635676608788779303912058663610140895306929917145003987389196141625913557220658030547435813332844544;
    data[159]<=640'd124267627527239871678891840804649687882769951686632598038723971608628918962446209350271372025099339623779758330106028752896;
    data[160]<=640'd83905163280176801464012698019748121716720079466359176019143954778143538017239804233030443734262617003489531235793257889792;
    data[161]<=640'd248785534760584653829688623609967533851115756283619978231422899164086156723362482793588001679810877897340761800704067108864;
    data[162]<=640'd331177968508717496025908651935120961056692808154220651851004904720080380783725440468588847857072075199627487004929936064512;
    data[163]<=640'd165265260449864111829202825648925674293649232615041886122956696078624808668973085763024810676371654190889504500713967845376;
    data[164]<=640'd165267779715684320620961849185177811961334566688885920530937850621598995701852315270803719875713339180682117787409732075520;
    data[165]<=640'd330545653733327795944282081865537304573994668389092076074639336040380473355487794842089930097357047428012127295467415404544;
    data[166]<=640'd495817208653531770068616519070605095398150325729412143847154655381398412673715979410714740495043248482513984734191849308160;
    data[167]<=640'd495867643221237691760492610798506576553438520994205361642203099489650897001502841281568289543367211468310948088416571490304;
    data[168]<=640'd578444161295294245496271641010504244283599178486672007018932580082024435758079946554061904553009889095322418030048828194816;
    data[169]<=640'd83237220765511686684021423737006202602597947375105159168295141516972863607240618121946062636588045421255064872251077689344;
    data[170]<=640'd159373254365344073560690679311151216189196216325241750827408215498597240214806707974611944243819788144477602656871658815488;
    data[171]<=640'd75853619720828376931961896625639622706042950583308679420399059379970735302554522121496000481012886606018049061380924899328;
    data[172]<=640'd5164509606816279191259417406678059472741344017281339160212186800288490087028236722802972806320673153093413220686388789248;
    data[173]<=640'd162962878106758886901475655072750252884117471493274900050891235948350503981066936494671790080;
    data[174]<=640'd195555453728110664281770786087300303460940965791929880061069483138020604777280323793606148096;
    data[175]<=640'd912592117397849766648263668407401416151057840362339440284990921310762822293974844370162024448;
    data[176]<=640'd1825184234795699533296527336814802832302115680724678880569981842621525644587949688740324048896;
    data[177]<=640'd7822218149124426571270831443492012138437638631677195202442779325520824191091212951744245923840;
    data[178]<=640'd47976271314629816303794432853417674449084183607620130574982379863194388372026106104031374999552;
    data[179]<=640'd12515549038599082514033330309587219421500221810683512323908446920833318705745940722790793478144;
    data[180]<=640'd50062196154396330056133321238348877686000887242734049295633787683333274822983762891163173912576;
    data[181]<=640'd0;
    data[182]<=640'd0;
    data[183]<=640'd0;
    data[184]<=640'd0;
    data[185]<=640'd0;
    data[186]<=640'd0;
    data[187]<=640'd0;
    data[188]<=640'd0;
    data[189]<=640'd0;
    data[190]<=640'd0;
    data[191]<=640'd0;
    data[192]<=640'd0;
    data[193]<=640'd0;
    data[194]<=640'd0;
    data[195]<=640'd0;
    data[196]<=640'd0;
    data[197]<=640'd0;
    data[198]<=640'd0;
    data[199]<=640'd0;
    data[200]<=640'd0;
    data[201]<=640'd0;
    data[202]<=640'd0;
    data[203]<=640'd0;
    data[204]<=640'd0;
    data[205]<=640'd0;
    data[206]<=640'd0;
    data[207]<=640'd0;
    data[208]<=640'd0;
    data[209]<=640'd0;
    data[210]<=640'd0;
    data[211]<=640'd0;
    data[212]<=640'd0;
    data[213]<=640'd0;
    data[214]<=640'd38929182122037745461731691618941890439418782399219861307932913883394773110239244084077295059826296653116948454423134208;
    data[215]<=640'd1291046135031061505869535027921305649937242736936070825521993781683515319564877602893599848107559145886669972730393133056;
    data[216]<=640'd18055496515423413365276322777409609302812129563819545350227290072974751053127338796153250540105953973411947597022214750208;
    data[217]<=640'd82470605481400643082138652619252170501310444386267222967735874661305549943708397866742310911633401211388186946350901886976;
    data[218]<=640'd320521766117565711202037534099695697186222762332596553152740522223202713393153438447615719706717471778846933715319200415744;
    data[219]<=640'd620869705062549266536390539167933624313234481109932054178173912046121343322769067012673139883613903609773809648810881712128;
    data[220]<=640'd331496328099416284367409719038798207289463138502561071189831528175388467640298117196681180661111548906577608776813587202048;
    data[221]<=640'd968343704310773232114255688235803220035111716639467007898397097151230349914701956287492308801616074769080913926163529728;
    data[222]<=640'd322781234779651914369180562323492329065527920322658399495098978533239280524362821529622536707726820916566046120848916480;
    data[223]<=640'd2259468643382410037935503141960639355157758753026579853258726891236498714652682765565097131205509436528130994440746565632;
    data[224]<=640'd645562469578312638678630707527707197054692427151329177704128070431882678859673650421951288316925091034804421409397276672;
    data[225]<=640'd1291125554720277624250720490875906185734967586205234298597207637887123217880031044420265358444843380936398971101991927808;
    data[226]<=640'd1936691873100890181891786366878820693166437522068143884602055924500428013704979488431495800346306596007785888864303841280;
    data[227]<=640'd1291144563648463385934397400398349929479801175090126216652584759082937432949726088499138960317748332431584824920918458368;
    data[228]<=640'd3873404600069790959497017545873283413496196929998486181617205052868255985879219182150823057994973991156093560971459559424;
    data[229]<=640'd3873493562111293306954949428757348114837916349282627642841425092676757948939344976130417937565660655682777545220223401984;
    data[230]<=640'd3873494100773019948643845191273251309093454797732732613176471150891358655704895668513368610949626828856049034731121016832;
    data[231]<=640'd5164814356792502464542594995814879384466715788399621512445380166691299729923511197506107277483257261807910793314954117120;
    data[232]<=640'd7747378835122329812820232278881847819485358454558461870741794453524254432321433128291939334324473316578322118972339650560;
    data[233]<=640'd7747360365807836843252042804847180442991450006983807322397597471707256612921682641374532203785690257015193491148281741312;
    data[234]<=640'd12911406998985697352737087159319754249501051872512942600988306685465602467376585074631082912533798477266550779396331929600;
    data[235]<=640'd15493972093122469519352737048157710448476529073414391041002890325200132401637242330785958755960323614970397508796330016768;
    data[236]<=640'd15494051050748336135686709486344915052536481668757253615893672797995649252143868374270699002933005239754666328793884393472;
    data[237]<=640'd15494129547005949764558829156897985642550533467367048220294200067817381029761949091533218335362178377656638240139362959360;
    data[238]<=640'd10329314420679417046764065083613375060987939733154228023493064440869482740160581754105585510392638046160452338642942164992;
    data[239]<=640'd68953576604029475691364307617098708583009663372846376398801639479363309003783685511018146551155855975014191631171584;
    data[240]<=640'd0;
    data[241]<=640'd0;
    data[242]<=640'd0;
    data[243]<=640'd0;
    data[244]<=640'd0;
    data[245]<=640'd0;
    data[246]<=640'd0;
    data[247]<=640'd0;
    data[248]<=640'd0;
    data[249]<=640'd0;
    data[250]<=640'd0;
    data[251]<=640'd0;
    data[252]<=640'd0;
    data[253]<=640'd0;
    data[254]<=640'd0;
    data[255]<=640'd0;
    data[256]<=640'd0;
    data[257]<=640'd0;
    data[258]<=640'd0;
    data[259]<=640'd0;
    data[260]<=640'd0;
    data[261]<=640'd0;
    data[262]<=640'd0;
    data[263]<=640'd0;
    data[264]<=640'd0;
    data[265]<=640'd0;
    data[266]<=640'd0;
    data[267]<=640'd0;
    data[268]<=640'd0;
    data[269]<=640'd0;
    data[270]<=640'd0;
    data[271]<=640'd0;
    data[272]<=640'd0;
    data[273]<=640'd0;
    data[274]<=640'd0;
    data[275]<=640'd0;
    data[276]<=640'd0;
    data[277]<=640'd0;
    data[278]<=640'd0;
    data[279]<=640'd1291124939043454294827959586001505937164852896414611756415329678270323811008420597314822676640068915717951585986373746688;
    data[280]<=640'd1936687408565181442241939379002258905747279344621917634622994517405485716512630895972234014960103373576927378979560620032;
    data[281]<=640'd5124152101828709232598464606943476688123009932645490408273339660635347624939669245593202497915273509255620356883420807168;
    data[282]<=640'd20574781987608484723900328046728343134568703981807649853419349652956337736883622574110535172194329306882394355034272825344;
    data[283]<=640'd15157478959678599992587853388093769736564193573930876516267103034997204975517413888555734817241785578504697407694744584192;
    data[284]<=640'd40025818758495797753917149887304828068324539539897874698572171523313236931281710570433604284015140020298365305441667252224;
    data[285]<=640'd9038348936519407857828186687846879454953441463533967114265174084449029585800997627482992342587753145491613171705314279424;
    data[286]<=640'd5164740477805426717081199863110190561373947107147187512742294347125637432742843686351660306230421085417864677310303567872;
    data[287]<=640'd2582487521436782887357284228427715698872565510041432819650456648013121093622275588730252125432575876705660290597677694976;
    data[288]<=640'd7746986046297906429341647238841117623736199150373736422927498811379487281412015186361187343043875344578840689145670533120;
    data[289]<=640'd15493499268521454978183439067285312543682442508467148020355783875455751444528333731847836437447241201330844406279311458304;
    data[290]<=640'd15493972092595815152181910400873781683491925828556049131665873477967409858033762242984434910378206270753997707391835045888;
    data[291]<=640'd36153704807987421171937199945844226972962883089087499146583833387831364111004768864466794496898333526620075931821775257600;
    data[292]<=640'd20667455513693044865468130597792877856431817174040845482214734574646873839872593312129034401442615240299639370762611064832;
    data[293]<=640'd31022310130279954549178333705624203479322036579500479168616778254029562647171738011817964225772267173657640017588880670720;
    data[294]<=640'd62528784728162303758479010243345818990683938601787262303179721967070057938660837397010106127513002260163467972233773711360;
    data[295]<=640'd19810713073044998196207609079285314220380035954309401747865219652534955913557813824861450205417380192736573696776104574976;
    data[296]<=640'd60682882002392362654582655090742823889179229976520581340556202358644981804332384862256414810852773021141569904621188546560;
    data[297]<=640'd103290009923287154666797239698334318115860538374021682697862458384158711946500782191872882782413240194543178751936896696320;
    data[298]<=640'd123948018803298499685126822693698306850088276792921228583958908017810997750045547436703638693231164330720116193625020301312;
    data[299]<=640'd123948023767032470051823616631088274869677888524990405430018008758599289544360491390058812744411195890712618240555068948480;
    data[300]<=640'd123948023757422252155634139255458759186626489157144101022547248693418335289637904212517790084249830171929056759174792216576;
    data[301]<=640'd247896017905631432011243208295929967200084047885466124501071684549170169987967118880087218708037459702493772169166146502656;
    data[302]<=640'd165264051435265113634664211828211824418415542895467217787434873587059232038872106691058493334226444463748974916394844946432;
    data[303]<=640'd247896047514844504544205559518633753862412823429894946140450796406789702988959046215618614441820408612489589421078439002112;
    data[304]<=640'd247896027813878964931067788810478057099034557805151197150407690301773559261072909016444827565784426556202092503548513222656;
    data[305]<=640'd578423992507943841682373266476432151034268918217644568645547330810477906213192869371646209431673883803108054410845113810944;
    data[306]<=640'd495792094914253479680401459309330820914516270728544093745822009315876347208539271511276287250365244564367615103603105071104;
    data[307]<=640'd330528023874162772857870292793393649649750878062688640624799166853527395779130449388073160852019119334936810419867858501632;
    data[308]<=640'd36695977855841144185773134324833391052745039826692497979801421430190766017415756929120296849762010984873984;
    data[309]<=640'd0;
    data[310]<=640'd0;
    data[311]<=640'd0;
    data[312]<=640'd0;
    data[313]<=640'd0;
    data[314]<=640'd0;
    data[315]<=640'd0;
    data[316]<=640'd0;
    data[317]<=640'd0;
    data[318]<=640'd0;
    data[319]<=640'd0;
    data[320]<=640'd0;
    data[321]<=640'd0;
    data[322]<=640'd0;
    data[323]<=640'd0;
    data[324]<=640'd0;
    data[325]<=640'd0;
    data[326]<=640'd0;
    data[327]<=640'd0;
    data[328]<=640'd0;
    data[329]<=640'd0;
    data[330]<=640'd0;
    data[331]<=640'd0;
    data[332]<=640'd0;
    data[333]<=640'd0;
    data[334]<=640'd0;
    data[335]<=640'd0;
    data[336]<=640'd0;
    data[337]<=640'd0;
    data[338]<=640'd0;
    data[339]<=640'd0;
    data[340]<=640'd0;
    data[341]<=640'd0;
    data[342]<=640'd0;
    data[343]<=640'd0;
    data[344]<=640'd0;
    data[345]<=640'd0;
    data[346]<=640'd0;
    data[347]<=640'd0;
    data[348]<=640'd10487868401331496898807585777695826548180904680055410732287804945168509238250041531703803734660247305607345011947907055616;
    data[349]<=640'd33567987550931527042192156306755949770644412755123250772505197289639483223122247619445824336121635491366235423550027595776;
    data[350]<=640'd40983129901043396874109373421282176739849979047910684111839722521971294094743850678829097931160937535640916358301847912448;
    data[351]<=640'd81986433629390866106210768371857437923388361795860884755112300482925170293440511634897658039478343291999472757504521273344;
    data[352]<=640'd80049746220957313136537731177049547250464259824945163578347651955773232275597975016629894344622994423222641711927703633920;
    data[353]<=640'd154934992685289778829937480506905733158282580854802590846524107705795430036363792938880440914269895614993052202894826143744;
    data[354]<=640'd123947994148171722391417687779577127287228852555975886850991129191445025261072667914521029204717403269813901540724834304000;
    data[355]<=640'd123947994148171722391417687779577127287228852555975886850991129191445025261072667914521029204717403269813901540724834304000;
    data[356]<=640'd123947994148171685695439831938432941514094527722584834105951302498947045459651237723755011788960474149517051778713849430016;
    data[357]<=640'd289211986345733982217330082311202444563732997797219349907272808087540412474414794943116384061917011842602253833013628502016;
    data[358]<=640'd247956569111891838650295335541858530628361743745492990496389085217804157541446560019561630232560037188043109329361566695424;
    data[359]<=640'd83176758848144294367017695660088990569278193067569090928196085937231065631900623246928107461653286883669468811055398387712;
    data[360]<=640'd500472334356507408425562582227736496116680348192492945195435436356947296161180102701029571510891115323328124417597671211008;
    data[361]<=640'd430590203495621805269960966579735577804583963311167696788670382008770148828792621239591563550127246237623151308576395362304;
    data[362]<=640'd645562486144450419708749214420470671033498413561655625677346140185743135094288540927629970629788348393985766583054270201856;
    data[363]<=640'd640397988236146309065922354194940267787939609839108531212258974703154339261855668738433879671340131994724939699532209324032;
    data[364]<=640'd495791991370543947719500080388867750595105731106027018332806792160519617963986357545232994253646082407213921367433265807360;
    data[365]<=640'd991583985200706267504236064826016513730073177633111601526145511013350726015654773678510534934883972139678172057136267264000;
    data[366]<=640'd991584029528564465349215279946276333424416778626826455532293542342081872280804012123301812537460215828794768752568931713024;
    data[367]<=640'd1983168146478526792386308508944325132031922298929950050371695150365790655111435119597610508213920198832616049554534491488256;
    data[368]<=640'd1322596664758873968128922443211502164112682381381292908348498814146758016159272295362547325660303008699594837256716068847616;
    data[369]<=640'd1984944149426938944743395867703134735197302288756059192831604483222748189105654609089201513879210901651763231281881186041856;
    data[370]<=640'd3314965174448771204626570810911707569255032041584737201036514885496795692659864257600143081630544960229759741999092588347392;
    data[371]<=640'd4190999117939507208313675146282384572004464906097833945061690727723027305355123634325855550704666441367683355882898585550848;
    data[372]<=640'd3956006814157438689272146538789421847143643777361946025677446416539872098366788152826251960241793666700552011039081993601024;
    data[373]<=640'd1322111937582902362380436012178910208199861920878332506714658496943901707037421685027457901835835901311606375536028312141824;
    data[374]<=640'd0;
    data[375]<=640'd0;
    data[376]<=640'd0;
    data[377]<=640'd0;
    data[378]<=640'd0;
    data[379]<=640'd0;
    data[380]<=640'd0;
    data[381]<=640'd0;
    data[382]<=640'd0;
    data[383]<=640'd0;
    data[384]<=640'd0;
    data[385]<=640'd0;
    data[386]<=640'd0;
    data[387]<=640'd0;
    data[388]<=640'd0;
    data[389]<=640'd0;
    data[390]<=640'd0;
    data[391]<=640'd0;
    data[392]<=640'd0;
    data[393]<=640'd0;
    data[394]<=640'd0;
    data[395]<=640'd0;
    data[396]<=640'd0;
    data[397]<=640'd0;
    data[398]<=640'd0;
    data[399]<=640'd0;
    data[400]<=640'd0;
    data[401]<=640'd0;
    data[402]<=640'd0;
    data[403]<=640'd0;
    data[404]<=640'd0;
    data[405]<=640'd22835963083295692796307572051946513295317401600;
    data[406]<=640'd45672100391163898150213262013115221110251585536;
    data[407]<=640'd45674887984313715745755515285502472364555763712;
    data[408]<=640'd12141579755374989211971784270440595481417482240;
    data[409]<=640'd92102251995525334173434820194839742216740536320;
    data[410]<=640'd92105050472393346222340006026735071894232367104;
    data[411]<=640'd40724134896108405176044034151206948129852096512;
    data[412]<=640'd5753778746591798124127606355191857860434722816;
    data[413]<=640'd188444269634341370752959454699504880840286928896;
    data[414]<=640'd182866110978867964976108728753656975618518024192;
    data[415]<=640'd154742504910672534362390528;
    data[416]<=640'd0;
    data[417]<=640'd0;
    data[418]<=640'd0;
    data[419]<=640'd0;
    data[420]<=640'd0;
    data[421]<=640'd0;
    data[422]<=640'd0;
    data[423]<=640'd0;
    data[424]<=640'd0;
    data[425]<=640'd0;
    data[426]<=640'd0;
    data[427]<=640'd0;
    data[428]<=640'd0;
    data[429]<=640'd0;
    data[430]<=640'd0;
    data[431]<=640'd0;
    data[432]<=640'd0;
    data[433]<=640'd0;
    data[434]<=640'd0;
    data[435]<=640'd0;
    data[436]<=640'd0;
    data[437]<=640'd0;
    data[438]<=640'd0;
    data[439]<=640'd0;
    data[440]<=640'd0;
    data[441]<=640'd0;
    data[442]<=640'd0;
    data[443]<=640'd0;
    data[444]<=640'd0;
    data[445]<=640'd0;
    data[446]<=640'd0;
    data[447]<=640'd0;
    data[448]<=640'd0;
    data[449]<=640'd0;
    data[450]<=640'd0;
    data[451]<=640'd0;
    data[452]<=640'd0;
    data[453]<=640'd0;
    data[454]<=640'd0;
    data[455]<=640'd0;
    data[456]<=640'd0;
    data[457]<=640'd0;
    data[458]<=640'd0;
    data[459]<=640'd0;
    data[460]<=640'd0;
    data[461]<=640'd0;
    data[462]<=640'd0;
    data[463]<=640'd0;
    data[464]<=640'd0;
    data[465]<=640'd0;
    data[466]<=640'd0;
    data[467]<=640'd0;
    data[468]<=640'd0;
    data[469]<=640'd0;
    data[470]<=640'd0;
    data[471]<=640'd0;
    data[472]<=640'd0;
    data[473]<=640'd0;
    data[474]<=640'd0;
    data[475]<=640'd0;
    data[476]<=640'd0;
    data[477]<=640'd0;
    data[478]<=640'd0;
    data[479]<=640'd0;
end 

//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)   pixel_data <= 12'd0;
    else begin
        if(data[pixel_y][pixel_x] == 1'b1)  pixel_data <= WHITE;
        else pixel_data <= BLACK;
    end
    
end  
endmodule


// The whole VGA 
module VGA_out(
    input sys_clk,
    input sys_rst_n,
    //VGA
    output vga_hs,
    output vga_vs,
    output [11:0] vga_rgb);

//Wire define
wire vga_clk_w;
wire [11:0] pixel_data;
wire [9:0] pixel_x;
wire [9:0] pixel_y;

//****************************Main Code**************************

clockDiv clkdiv1(
     .sys_clk(sys_clk),         
     .sys_rst_n(sys_rst_n),
     .clk25MHz(vga_clk_w));

vga_driver VGAdriver1(
    .vga_clk(vga_clk_w),   
    .sys_rst_n(sys_rst_n),
  
    .vga_hs(vga_hs),      // 行同步
    .vga_vs(vga_vs),      // 场同步
    .vga_rgb(vga_rgb),      //4+4+4
    
    .pixel_data(pixel_data),    //像素点RGB data
    .pixel_x(pixel_x),       //像素点横坐标
    .pixel_y(pixel_y)        //像素点纵坐标
);
 
vga_display vgadisplay1(
    .vga_clk(vga_clk_w),
    .sys_rst_n(sys_rst_n),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .pixel_data(pixel_data));

endmodule