`timescale 1ns / 1ps


// VGA Driver
module vga_driver(
    input vga_clk,      // VGA驱动时钟
    input sys_rst_n,    // 复位信号
    //VGA
    output vga_hs,      // 行同步
    output vga_vs,      // 场同步
    output [11:0] vga_rgb, //4+4+4
    
    input [11:0] pixel_data,    //像素点RGB data
    output [9:0] pixel_x,       //像素点横坐标
    output [9:0] pixel_y        //像素点纵坐标
);

// some parameters for sure in the reference Table 
parameter H_SYNC = 10'd96;
parameter H_BACK = 10'd48;
parameter H_DISP = 10'd640;
parameter H_FRONT = 10'd16;
parameter H_TOTAL = 10'd800;

parameter V_SYNC = 10'd2;
parameter V_BACK = 10'd33;
parameter V_DISP = 10'd480;
parameter V_FRONT = 10'd10;
parameter V_TOTAL = 10'd525;

// counters for H and V
reg [9:0] cnt_h;
reg [9:0] cnt_v;

wire vga_en; // 使能控制rgb数据输出
wire data_req;

//*******************************Main Code************************************
//VGA 行场同步信号
assign vga_hs = (cnt_h <= H_SYNC - 1'b1) ? 1'b0 : 1'b1;
assign vga_vs = (cnt_v <= V_SYNC - 1'b1) ? 1'b0 : 1'b1;

// 使能使RGB输出 // 范围内输出
assign vga_en = (((cnt_h >= H_SYNC + H_BACK) && (cnt_h < H_SYNC + H_BACK +H_DISP))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;

//在范围内RGB赋值
assign vga_rgb = vga_en ? pixel_data : 12'b0;

// 请求像素点颜色数据输入
assign data_req = (((cnt_h >= H_SYNC + H_BACK -1'b1) && (cnt_h < H_SYNC + H_BACK +H_DISP -1'b1))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;
// 像素点坐标
assign pixel_x = data_req ? (cnt_h - (H_SYNC + H_BACK -1'b1)) : 10'd0;
assign pixel_y = data_req ? (cnt_v - (V_SYNC + V_BACK -1'b1)) : 10'd0;

// H counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_h <= 10'd0;
    else begin
        if(cnt_h < H_TOTAL - 1'b1)  cnt_h <= cnt_h + 1'b1;
        else cnt_h <= 10'd0;
    end
end
// V counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_v <= 10'd0;
    else if(cnt_h == H_TOTAL - 1'b1) begin
        if(cnt_v < V_TOTAL - 1'b1)  cnt_v <= cnt_v + 1'b1;
        else cnt_v <= 10'd0;
    end
end
endmodule 


module vga_display(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input [1:0] choise,
    output reg [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;

// some frequently-used colors define
localparam WHITE = 12'b1111_1111_1111;
localparam BLACK = 12'b0000_0000_0000;
localparam RED = 12'b1111_0000_0000;
localparam GREEN = 12'b0000_1111_0000;
localparam BLUE = 12'b0000_00000_1111;

reg [0:639] data [479:0];
always @(posedge vga_clk) begin
    if(choise == 0) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd0;
        data[47]<=640'd0;
        data[48]<=640'd0;
        data[49]<=640'd0;
        data[50]<=640'd0;
        data[51]<=640'd0;
        data[52]<=640'd2293498615990071511610820895302086940796564989168281123737588839386922876088484808070018553110125686554624;
        data[53]<=640'd1675976290930685468645128323187019804819274807935478584355997288644324119240316295174021690532034581474959799140168891292198173855926923755850975816974336;
        data[54]<=640'd4608938271443963528941588642716363415553844460538933171124528709463054170393956612499412155428494782625729343881662003406464265768870265575791175453900800;
        data[55]<=640'd32262541127990939173762083020509032968594440138823179507501159485634574000849247021006776338229579036834994698149052345903902864697637648985753025844871168;
        data[56]<=640'd58240171439706361472169453622740139551676880264982424390591317149858243932624905087835037248725775054926940671759288438860704227669296539774404515090923520;
        data[57]<=640'd42318407564523126557606423241263499508701606765135631683196970909087290531237324837141462551277584976845020334793376876887606858787731732121488036166893568;
        data[58]<=640'd395530370495227042665516596148738352043683483543209051664862984962215722154818246074688097346266051782000026180473705838717361763032412721084388760520491008;
        data[59]<=640'd875906954421202713545704567525854790768358994252243776699793848151799154343056753832682919968808972452753249328458824810904489328815372625029041313741275136;
        data[60]<=640'd1074300936946527189448081477115531402820708126955742360356077044371693182696136319406376230962391213472250986774014381769145217585253263421021236472190074880;
        data[61]<=640'd2723731004535675457407407214648210750903770826922016861520642014671865412833960365204224421091120348781355315742556081222814866948425965607358914138996736;
        data[62]<=640'd5363542192147591106665945431975488483211153355654328491357949574079026346254569789205797302263463966091837288140978704750469707812894644221288083022638219264;
        data[63]<=640'd2148392389880624983854794822778637342357380469688204162829970252499582343647074513421659901813271610738497426696471688412865232369391466669779185154318663680;
        data[64]<=640'd11157393520650594033816653652288795059042270346749989081083521077635666177081536011080883761299459976071350897937465882988689764126215296351421545708670418944;
        data[65]<=640'd46340318392186936871323099658801396008038326033905033280090403424319477039293533746461577656164197176237198767912607413258782486604516713763506551490862907392;
        data[66]<=640'd6866894267813936637844109936851291657023550013168452068701946928148428461883378977066012880698571175098621288248210288500459301797733256446001671825596088320;
        data[67]<=640'd6866055871643455633919549855401627155405683307443407615500233076853761656628263449134380842739204401454157064456222742542119398180196937364232137528850776064;
        data[68]<=640'd82380932058025304369882760701860083250682292991484941806457284014125123379755651628509720405156100616276445336341233578718530541909729839781497329850521747456;
        data[69]<=640'd123568046953902601885489631601050712319174756009461312869005805972744294597349989309378349784223221026846516048020819811265697562604659577532981444669203283968;
        data[70]<=640'd288324856952856638938360058898595805306574222331048332226622281617419903733234488006034233947574894938995849281914303336068168613552865455582601091901248503808;
        data[71]<=640'd604109837461759778168159595812366405561914221390916897199734931180272979632225765748065127120840811121811655347422247737108184549641653972618942044609571717120;
        data[72]<=640'd604113173047588395015331192328821260737655662434528286280150192127775494254945644991600158879780428058664007014154694790222100112847793335065517706788783259648;
        data[73]<=640'd219675266569980855101283472340255299678830543246909919602823875385570340106129550504925267063655400482168152660230457948423843364412407532088987667975607681024;
        data[74]<=640'd878716280995473004337282926076232960710252933604169513785718377197055657451630564829885256010195180777820288365803555872444941845579307383195420644215244193792;
        data[75]<=640'd1867228394076075483794978113422141474529413092464248978844049179274668247592540852714362839805123260305110545725523235818229294611325658936654682330078214356992;
        data[76]<=640'd2196759186277915900926322250153514691466961015354738301595353246150210141478551945047509799424682666003850921931081454547645667767808867014961711369790485954560;
        data[77]<=640'd5491840118327575789266050286268835412211319625532502477095620565199695451401293084153438916689517108918215411578931448829559414360696935030298648443765439594496;
        data[78]<=640'd3295140691075790202280104419051183345307264370081109106149563130065548234442196278888186533097198155681390201425625669533083696367444166288535752857087247384576;
        data[79]<=640'd12301738147164137008516192307349284430213059126345595918172653360353590957845406813189173483570374230403960158616455187826875596110565138928530713386938705903616;
        data[80]<=640'd10983694272968463208017411114256965826893096936854354198107273535794206413204309036433666244710318396426212727686533691447454945851282655205826496843257263161344;
        data[81]<=640'd16695249082583700151819180632048177262635343246267534392840559284858924655228845405174144134607644664658356352874643028256124293023562727569268576201652675018752;
        data[82]<=640'd15816562523961361330229573309826634226434290288366856178771999537978267005376446045370118187440417277347052876463276094705521338392416505356020586531298431991808;
        data[83]<=640'd36026489125927671166289176420646080071866189211135292775156866507934099707732327272359078617095675212156124947774533078691482697388957364701881514429016937857024;
        data[84]<=640'd5272240021943069727947564190292979055793729966361248715538640052077095891112436303112593429210693090570943905958303872941466164741451264206416949289102920908800;
        data[85]<=640'd29875653048126526639798045377648067050180185090282107520280915163244183757325856740083861989077872004946784096482024153935771661077851379083361887904318372184064;
        data[86]<=640'd63266116017769340614370302764131239925710436011546193109013856643390801955703664349384433193504743177508980454909012615578815823764973452731200254228423507968000;
        data[87]<=640'd31633061360863825370210645136310830404209726733791878434705385420389778471631909814652699262398831417058366293186418192618503535676488482274630290480730283704320;
        data[88]<=640'd63266263503656570665825684773802091766755078915378435853240554166128374162234725728383526188788462984391661037890014737274341293996581484529175727360672803061760;
        data[89]<=640'd70295581671023508211478452617564891644709630344406242109297818921681604012213781017281502757906308516323092188893825690710699206741894451723342734933425752375296;
        data[90]<=640'd140591176749765437835789265421574959863756815093899739696031636517167324564256131031003711274920578246666233112393967661926318979829304773066559488652826841710592;
        data[91]<=640'd56236690588038060701510754154057083807847535199944312387298568698492464460505779782646578450388672046384196427450360965925681982269874295247584323200251139719168;
        data[92]<=640'd337418775931314434710666121368382058581550402986087022736596132649012604514048986252565250960473903116455606423577632442273831910856563706269486414050219291312128;
        data[93]<=640'd84354740910148374275949364164703432233673625957957103591082717251868282624564948702530145342028491063265353316901573768218354216004237376400809978444917485076480;
        data[94]<=640'd112473113019738508644751981776265581042538941086922546215314451586728435496034081217546402872535840442426955979921003800584349379723459316631560600633045759819776;
        data[95]<=640'd309300537899771631082660610980791466418600909513341640781873249643700485657286888528662428914250860760547729443177382375785407577796792937338398326762111705808896;
        data[96]<=640'd56236422431789954785131731391502193504346644638376045558492893439990743552035552631576808305257788610793059377749037847322670386405301057230994913620053708505088;
        data[97]<=640'd0;
        data[98]<=640'd0;
        data[99]<=640'd0;
        data[100]<=640'd0;
        data[101]<=640'd0;
        data[102]<=640'd0;
        data[103]<=640'd0;
        data[104]<=640'd0;
        data[105]<=640'd0;
        data[106]<=640'd0;
        data[107]<=640'd0;
        data[108]<=640'd0;
        data[109]<=640'd0;
        data[110]<=640'd0;
        data[111]<=640'd0;
        data[112]<=640'd0;
        data[113]<=640'd0;
        data[114]<=640'd0;
        data[115]<=640'd0;
        data[116]<=640'd0;
        data[117]<=640'd0;
        data[118]<=640'd0;
        data[119]<=640'd0;
        data[120]<=640'd0;
        data[121]<=640'd0;
        data[122]<=640'd0;
        data[123]<=640'd0;
        data[124]<=640'd0;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd24084754561361768648102764881807084833480156810453237320207177473645930965106688;
        data[156]<=640'd74106937111882365071085430405560261026092790186009960985252853765064402969559040;
        data[157]<=640'd70608395103938906748405107852975316393858956036050582890626880237652602651358048951934797737936631459539297024459407360;
        data[158]<=640'd45391111138246440052546522188883403559323054846082361826329892174494524730641999395236457398525145100652968239135981568;
        data[159]<=640'd1636695303852802729735721062056598689171227159782417379487311097989030145039228099523491731237091973850787271799481790412816552786667439353248692043776;
        data[160]<=640'd1636695303852802729735721062055885040034998062974924581513017296855793489370356461447734507695151320981908907938792924355968481261496945489806448656384;
        data[161]<=640'd818347651926401364867860531031735199525939178478519424977370246509580297618296351778466869166585272986773102139318925346653358677398298558795786223616;
        data[162]<=640'd1432108391049830273401644278722737849120364334060297247134938174134513807501900800215425895994497321779674193266119508278048795711930628599338634313728;
        data[163]<=640'd1432108391049830273401644278735649098510798877008576842994953233506200279217848201550508752554026776391740998501303430948513796217162926072429574881280;
        data[164]<=640'd1432108391240366683943391851477633537586661023558736994503006139883435319970837805366295150217217232081572022588943456326054179354432327137873574756352;
        data[165]<=640'd1432108391240366683943391851560265533685442098427726409075096037822516832042486378403564082627356928761751483328526138566416523094507341434564099702784;
        data[166]<=640'd1432108391240366683943391851436317539537270486124242286682964431933796048692382457126427995832131793975102676007502805636927351288835714611939024830464;
        data[167]<=640'd1435305037176693300102889726780014576429566470681422420386847245326722576375588288221031848066714907782555811250039509689363615958633158073818902691840;
        data[168]<=640'd1435305037367229710644637299496199212568719915731594059278130643385491741978943949843963127844319033508265347311733950057284828604547490761026662563840;
        data[169]<=640'd1435305037367229710644637299827448417961298273229098846927417863473669561179014619152488000536355792201675587252827406296687614509099521024827229995008;
        data[170]<=640'd1435305037367229710644637299334373618732349678270996364183221587829367760609145726026744782561119957545428387402377148278373136728610751125342621007872;
        data[171]<=640'd1435305037367229710644637299993567271371739555789304069914834457587459522536104288487695019206776728729846866371242131408545259898951552500600571691008;
        data[172]<=640'd1435305037367229710644637299333487199138825454724606894071476206184202028858221877983831414751630822537736703386206619778425774892426268893339512209408;
        data[173]<=640'd1435305037367229710644637300653019438121440510868069007907168480577641826757956539973854350149827416275424392591229598479304825936053175413608078639104;
        data[174]<=640'd1435305037367229710644637300653034558641143412569597725777903431964866886898193444370075328131673110808604221924283288817759997577909217358664431566848;
        data[175]<=640'd1435305037367229710644637299991983623461348028344010791960645046074374778705467357024839583392402874487172079292395303024722442452133379642409980264448;
        data[176]<=640'd1435305037367229710644637299330897443181561344417431113677107966919478585359131666779569300610786589534507938519752671279255654159513994981444495081472;
        data[177]<=640'd1435305037367229710644637300653029495482915038838613054143659807267775516853193537903920654581336503892994637717971373035093841031522860826515937951744;
        data[178]<=640'd1435305037367229710644637299992114802589490987460098161908503990359874513499613344915043052155791646944514578423600700997597789590847215077138546819072;
        data[179]<=640'd1435305037367229710644637299828787438695083915449891531911929626210393274776978887610931890986492201089081971266064718119360062608871443242470722240512;
        data[180]<=640'd1435305037367229710644637299437092528518306659726087176161919758242288498105904759736451027421619171134752812288730275521880220238638370174373946458112;
        data[181]<=640'd1435305037367229710644637299507781500724513233078128733369671170587125172353968989771482801333236989287052402859688069010439927259458017806736643063808;
        data[182]<=640'd1435305037367229710644637299361884422014369541227848242073100429670977541832460348276643557836512441370962158324081713487370893782277483959604217905152;
        data[183]<=640'd1435305037367229710644637299330897384075245286961408227572008944085624655223000009162103830482396664431885916192872312702111210533470150330521170739200;
        data[184]<=640'd1432108391240366683943391851436317539537270486124242286683225172538675800307101737124344943615829196905365418341429752739979471967507308473220046258176;
        data[185]<=640'd2864216782480733367886783702872635079074540972248484573365928863867409972176118752152457086422429217901952357002696653524924222322275202749657142788096;
        data[186]<=640'd1432108391240366683943391851436317539537270486124242286685050356773471499840398264461159746448131312586090097221999734582600997612095258161960370307072;
        data[187]<=640'd1432108391240366683943391851436317539537270486124242286703823680331370123611448259925540575580381645302115365707862404963850975670714169246146560524288;
        data[188]<=640'd1432108391240366683943391851436317539537270486124242286774745124883431591190970465013201485635549568895988602210010270848573115003274500008627723567104;
        data[189]<=640'd1432108391240366683943391851436317539537270486124242286716339229369969206125481590235127795001881867112798878031770851884684294376460109968937354002432;
        data[190]<=640'd716054195620183341971695925718158769768635243062121143341482215966852493044029688038114271605607304475488089250674163381231055580568800687414285697024;
        data[191]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[192]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[193]<=640'd0;
        data[194]<=640'd0;
        data[195]<=640'd0;
        data[196]<=640'd0;
        data[197]<=640'd0;
        data[198]<=640'd0;
        data[199]<=640'd0;
        data[200]<=640'd0;
        data[201]<=640'd0;
        data[202]<=640'd0;
        data[203]<=640'd0;
        data[204]<=640'd0;
        data[205]<=640'd0;
        data[206]<=640'd0;
        data[207]<=640'd0;
        data[208]<=640'd0;
        data[209]<=640'd0;
        data[210]<=640'd0;
        data[211]<=640'd0;
        data[212]<=640'd0;
        data[213]<=640'd0;
        data[214]<=640'd0;
        data[215]<=640'd0;
        data[216]<=640'd0;
        data[217]<=640'd0;
        data[218]<=640'd0;
        data[219]<=640'd0;
        data[220]<=640'd0;
        data[221]<=640'd0;
        data[222]<=640'd0;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[232]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[233]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
        data[234]<=640'd716054195620183341971695925720741019646722151651777062513485227841182198836858911550944930962147952097504930445303808734511193412004703859387033190400;
        data[235]<=640'd716054195620183341971695925733975050271917558173763648270000663697121941025108682054202060164418771160341241567780741170071899798113707615747364093952;
        data[236]<=640'd613760739123428908533783747742740951106836389501670883432644008300727774996090104408282560325565701807498331942556538594674181096568959768677637423104;
        data[237]<=640'd716054195620183341971695925775162440173083066321608092275360877847400583774061544656682464485426853248945059637532466554010146754313959091645976674304;
        data[238]<=640'd716054195620183341971695925800790765867416322518107788925878604051471834800992816686952080507283765768598800843670835018201524272156680838057939697664;
        data[239]<=640'd613760739123428908533783747723284561819669846476611648565846264090512837504587917674511322608938258333246860517141884398558060687551093066887677870080;
        data[240]<=640'd716054195810719752513443498454979356758800439428213205417422927204079958898775110336209128697962308883265212617858920508814207947400500444495681159168;
        data[241]<=640'd716054195810719752513443498434320710063628303715722104264378486736449078009609937506835143563140728989218382396221405478484941207118017931440805642240;
        data[242]<=640'd716054195810719752513443498506624652298210471454580631817978684638221256651682055343100676463891433662762449512291550250352994498084041687198964121600;
        data[243]<=640'd716054195810719752513443498454979339520422719331634086085317577553004449140326088157082167534735801866357466995654626418694858991575285603261409656832;
        data[244]<=640'd716054195810719752513443498475637968977217134947546067972745522638726218803218737963866474074639029707315953979441524666868439552122893476093667311616;
        data[245]<=640'd716054195810719752513443498516953967026682825744689537321206210830870755031356310792626601131510055948434664690725965774794625032834905303444631846912;
        data[246]<=640'd716054195810719752513443498475651838503407857783457612004023740012272049318143742879487223216607915566096410483134765841002218758775178906054867025920;
        data[247]<=640'd716054195810719752513443498516972889851300130421028016039157347335497661769359591841987425384638752091307413007997007491500789825376896002756962156544;
        data[248]<=640'd716054195810719752513443498477129571367123143256409622961880200894187855801381105167642950423942030140195393554408533171113187586288060610244853628928;
        data[249]<=640'd716054195810719752513443498688349581229667683819234323872614482215359658453377902801690390410282977332645815467658880462739171969499039438989399425024;
        data[250]<=640'd716054195810719752513443498467889978237535413865193261722516837795240857176937423000817673609967888972696308019079950730225735760304001403993255313408;
        data[251]<=640'd716054195810719752513443499012744682755095901190603710942458311937664230556259154779137599693269315475229028829709518779086258855941445733184438272000;
        data[252]<=640'd716054195810719752513443498434320749542647963546615847128590290717972407571799454286011043581789429640321044974277537475434800497574688132935473692672;
        data[253]<=640'd716054195810719752513443498764848812664846345737906278997849975982598580447173321169773869957056320881961665510260061692698207071969379802162304909312;
        data[254]<=640'd716054195810719752513443498599584702492099270351629887921327346536436747285995343650763722514606921429714685427165654562488330188806306396538197245952;
        data[255]<=640'd716054195810719752513443498434320828500781206688941497732121774492216533516931710521477415365599104042734973635925821243467354688783545621977073975296;
        data[256]<=640'd613760739123428908533783748022824438419078804462979289892749333281482296153378453386459831809598151032801689536472321311761208179628544868692954972160;
        data[257]<=640'd716054195715451547242569713067823772213345384943196004009009088356959474312158081546613895513026045545123624799960285426309255936814095547164780396544;
        data[258]<=640'd1432108391240366683943391852427901650330668318061077787476657549267738494399362547300808388636322370146902998225507789572748439002763179349185906343936;
        data[259]<=640'd613760739123428908533783748353352344318169347744232209393661628026371781389883644313105808740398310283400397837615645710834553518948867682674392694784;
        data[260]<=640'd716054195620183341971695927040270707349433226429013276887335984651203362723913070456874346558756487460550559558322364016292066238315886925744334438400;
        data[261]<=640'd716054195620183341971695927040270865264985409127194942397394261385077602193564080742068802475296351678528346700460949113592381895506742197185683652608;
        data[262]<=640'd3273390607705605459471442124111437211921649132173375251991851805594240128964229260320230813883475049558263568760263610208291932078864297492040906702848;
        data[263]<=640'd776790931223330254907009681665451926923432634146589683220239250695842456566297925992806072473548014703579287154640580429317990534798152161039138947072;
        data[264]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[265]<=640'd0;
        data[266]<=640'd0;
        data[267]<=640'd0;
        data[268]<=640'd0;
        data[269]<=640'd0;
        data[270]<=640'd0;
        data[271]<=640'd0;
        data[272]<=640'd0;
        data[273]<=640'd0;
        data[274]<=640'd0;
        data[275]<=640'd0;
        data[276]<=640'd0;
        data[277]<=640'd0;
        data[278]<=640'd0;
        data[279]<=640'd0;
        data[280]<=640'd0;
        data[281]<=640'd0;
        data[282]<=640'd0;
        data[283]<=640'd0;
        data[284]<=640'd0;
        data[285]<=640'd0;
        data[286]<=640'd0;
        data[287]<=640'd0;
        data[288]<=640'd0;
        data[289]<=640'd0;
        data[290]<=640'd0;
        data[291]<=640'd0;
        data[292]<=640'd0;
        data[293]<=640'd0;
        data[294]<=640'd0;
        data[295]<=640'd0;
        data[296]<=640'd0;
        data[297]<=640'd0;
        data[298]<=640'd0;
        data[299]<=640'd0;
        data[300]<=640'd0;
        data[301]<=640'd0;
        data[302]<=640'd0;
        data[303]<=640'd0;
        data[304]<=640'd0;
        data[305]<=640'd0;
        data[306]<=640'd0;
        data[307]<=640'd0;
        data[308]<=640'd0;
        data[309]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[310]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[311]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[312]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[313]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[314]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[315]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[316]<=640'd716054195810719752513443498444785882909390677394503417248096665387912638568274816216319923546195994976306584519426322962481530122975535690971336409088;
        data[317]<=640'd716054195810719752513443498455968487483977001750781907060838224134704709211147073704256992800668164780831664868630583039747908261161583167644333244416;
        data[318]<=640'd716054195810719752513443498474537234532114649602277376614592304150941807458703701962780977343526620605754526330208115812089993145710677900868284579840;
        data[319]<=640'd716054195810719752513443498469181083417895511379387966348654761088606061502328738306483090926155365809885569869539490452204505213097378866499214639104;
        data[320]<=640'd716054195810719752513443498460143208844760463077529821080196447904555248326788557900137008901452003884198374928910000939410338251252270873223882604544;
        data[321]<=640'd716054195810719752513443498527281705674757012943335194389606949037152868359891240043216593653491645666403208387701926563269058460469809487764755841024;
        data[322]<=640'd716054195810719752513443498496294707137714219955397731849003363864599373346113716124368161452497813606465404624444234571178191844129520710124740542464;
        data[323]<=640'd716054195810719752513443498434320710063628340411699960038642707334417784651430246326352683510526311075218355571800711260941025649074145058756830953472;
        data[324]<=640'd716054195810719752513443498558268704211799916019206224453643091529109337873841922197184505931979417130605302723257670802630712437700647551437725761536;
        data[325]<=640'd716054195810719752513443498516952706162409451976667229383883273086102694855356451481973609612325014781178703990715379981662365375319896323895735615488;
        data[326]<=640'd716054195810719752513443498682277239580970957473452572422737403252585741964642850032475924422476581956582228806857619203036121907734186946087295647744;
        data[327]<=640'd716054195810719752513443498434421638533521882075411746585902044686871280811745016078464176196770890654219677253771343330134798667677997582164607107072;
        data[328]<=640'd716054195810719752513443498520180528360673233561419094502815395445687106779796414844980695166071443563498360276778173398667954563354747162810074005504;
        data[329]<=640'd716054195810719752513443498996605656726023935176777716230020742777013287689054251465974486966298616100244663611899227079591643839540565529680693690368;
        data[330]<=640'd716054195810719752513443498573762205327292022636158609571585341487229762413136362358988649101210667449267486323672056625660151417107876774568232222720;
        data[331]<=640'd716054195810719752513443498682216713136626426241962318096820975062643994920880194237175984206851725341056316457898984997855816749784111530799062319104;
        data[332]<=640'd716054195810719752513443498599584702262693814274499031200694035285404404923758357194094993893866283716026817139533485184985118062016148369030003032064;
        data[333]<=640'd716054195810719752513443499425904673101307019081430866693741199808277343705677208242846533457381245478574006576665460295014574276902122092042165157888;
        data[334]<=640'd716054195810719752513443498764848716623583836033777364462676998056899305882677914285810678489932238168967027307797086834675354174885748935025999478784;
        data[335]<=640'd716054195810719752513443498434320870134880584172952545574899093982716409234873420460666315864822867744868192177266560455333762829457981149911869030400;
        data[336]<=640'd306880369823702018761794786331113062035674069665774299772575104062103108105134521081509791219496056458965289002349821463520873588929329112371016237056;
        data[337]<=640'd716054195810719752513443500419748086310216764306486793198588391973184409535139144672512889177745951175339461993074786741203682943285782144079475245056;
        data[338]<=640'd716054195810719752513443499756435170914068437240284981015065838044139534165305681635603031488482186828731043419821424621212064279135453754324680704000;
        data[339]<=640'd716054195810719752513443499144439427154387888478587444811613870182252570547413135394933489476212387257905581147685948894516168440858826323333314772992;
        data[340]<=640'd818347651926401364867860535221433105301380051923860736978214468308792128689640578898859583951849017517362481346889435950386937788282291303067668185088;
        data[341]<=640'd1636695303852802729735721063377830543543726744987234358969115182131310361193491873149574770423149332809446318453759619861197221749554275471993841123328;
        data[342]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[343]<=640'd0;
        data[344]<=640'd0;
        data[345]<=640'd0;
        data[346]<=640'd0;
        data[347]<=640'd0;
        data[348]<=640'd0;
        data[349]<=640'd0;
        data[350]<=640'd0;
        data[351]<=640'd0;
        data[352]<=640'd0;
        data[353]<=640'd0;
        data[354]<=640'd0;
        data[355]<=640'd0;
        data[356]<=640'd0;
        data[357]<=640'd0;
        data[358]<=640'd0;
        data[359]<=640'd0;
        data[360]<=640'd0;
        data[361]<=640'd0;
        data[362]<=640'd0;
        data[363]<=640'd0;
        data[364]<=640'd0;
        data[365]<=640'd0;
        data[366]<=640'd0;
        data[367]<=640'd0;
        data[368]<=640'd0;
        data[369]<=640'd0;
        data[370]<=640'd0;
        data[371]<=640'd0;
        data[372]<=640'd0;
        data[373]<=640'd0;
        data[374]<=640'd0;
        data[375]<=640'd0;
        data[376]<=640'd0;
        data[377]<=640'd0;
        data[378]<=640'd0;
        data[379]<=640'd0;
        data[380]<=640'd0;
        data[381]<=640'd0;
        data[382]<=640'd0;
        data[383]<=640'd0;
        data[384]<=640'd0;
        data[385]<=640'd0;
        data[386]<=640'd0;
        data[387]<=640'd0;
        data[388]<=640'd0;
        data[389]<=640'd0;
        data[390]<=640'd0;
        data[391]<=640'd0;
        data[392]<=640'd0;
        data[393]<=640'd0;
        data[394]<=640'd0;
        data[395]<=640'd0;
        data[396]<=640'd0;
        data[397]<=640'd0;
        data[398]<=640'd0;
        data[399]<=640'd0;
        data[400]<=640'd0;
        data[401]<=640'd0;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd22835963083295687686091080188131599678433132544;
        data[406]<=640'd22836137307867241909738992724944393428252229632;
        data[407]<=640'd45671926166590717540745122690701737417425027072;
        data[408]<=640'd11425168305238367630390631743024032890990100480;
        data[409]<=640'd92102251995524685136327182220460836482002714624;
        data[410]<=640'd174235205715414699939639567012653407666176;
        data[411]<=640'd79973270849186984475343595013176781527727472640;
        data[412]<=640'd758237586915271256831821758006986185344286720;
        data[413]<=640'd188399493930006087410775984133357220008931885056;
        data[414]<=640'd10634488215193846815244531305132589056;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
    else if(choise == 1) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd0;
        data[47]<=640'd0;
        data[48]<=640'd0;
        data[49]<=640'd0;
        data[50]<=640'd0;
        data[51]<=640'd0;
        data[52]<=640'd2293498615990071511610820895302086940796564989168281123737588839386922876088484808070018553110125686554624;
        data[53]<=640'd1675976290930685468645128323187019804819274807935478584355997288644324119240316295174021690532034581474959799140168891292198173855926923755850975816974336;
        data[54]<=640'd18016743004716045104939568706166646234830913194566828459917631673408091544086843037861291450401948673299982734405370585939836303642089739931020670818844672;
        data[55]<=640'd42318397475031701438889607385923245877036691254239602651234569147285240898305566161081713485969712312403657740930550414975923248456038202051341749537734656;
        data[56]<=640'd57402183344188992557480846249111134803883445987125003633414363911957637828907724366345008656219299889741061112297913938112867822288523357300753250694201344;
        data[57]<=640'd42318407564523126557606423241263499347310989384703844829702022658899048385630712785314992999361375193054543958740802212534772278779117267377539787870175232;
        data[58]<=640'd395530360905215115021967377632711409942006648779440471063266579816800946473045629048871445053568278627989595852987097636404105016876635012054155033330057216;
        data[59]<=640'd875906954421202713545704567352562934563026676853642611817926797221644961654863567688143481820911674474299584801504605189711145700733634866251699676946366464;
        data[60]<=640'd1074300936946526427302439310125071297515937130994533697009700542908227236054607196059323136753822689742996809766773833370569381539617161493151705275232681984;
        data[61]<=640'd2723730804743768237183904232934132161590198535360849222019756894908502785821633132584250944977698014866267721515232107944067370552804837045185415225540608;
        data[62]<=640'd5363542191748007292225498426358644037797628068518507929096833266769054255422522206636867302888064784899710315832520857566929660082277303334339182503433076736;
        data[63]<=640'd3142916103311877827994774634041287214440824010129971401946070220615944633674407965106679014548230495399058990158957803742790727468293186791713320095186944;
        data[64]<=640'd11157391883955290085745718645693946645242694238428966059551126335989982129014637808743606319664413813119272322494123819208654259517587023408725019044406624256;
        data[65]<=640'd46340318392186936109177457491811105143390564853932790665686560000254254661569666650423555483369856326553091574677262891816660630792352920929528114164621377536;
        data[66]<=640'd2096606884159293981315126535532627615023078102265478175759719763157201612263761929777286175608312879866159756539412255745900722075555602617940478057775104;
        data[67]<=640'd6866055053295803659884082352104202948505894945454718108404934879957895628581040891606397478280400890069828080887171596984391567232311544567374210143564595200;
        data[68]<=640'd82380930421130208514591602192456812614175954239596008503794331118824453286272729634887977963833354862728303274743662591346725013435792896395326352926655381504;
        data[69]<=640'd123566370976313023803090396825458558807077497481013248406508153003950354552629039991956389071662517411689116159875761730931895855458626834206801549764222517248;
        data[70]<=640'd233406472398421153322362982492754957452371837391271051293079320198475871542681979470129447661822803978026991749405005742697438182615596978466919612056934023168;
        data[71]<=640'd604109837461759778168159595812365051719290138961786243677184080065183411059435054900128032160108089138751203381785997749605204012738286105816714796771764600832;
        data[72]<=640'd604113173047588382820268264222886635157617763925308602241732751467439116477112097925475867510607460983621322460590903413775070191378235877211246055920150511616;
        data[73]<=640'd219675266569980855101260213501077829681437464241079911053085166377405662230442034181704214865795090685004559815270726763607027574337217172861509719847012925440;
        data[74]<=640'd878716019124224372645561183594217863774359502483167172018946154157074302914062729473940378033073734968744706476903378722072150697136375429262006661899186339840;
        data[75]<=640'd1867228367888950619673161100430435175904078019780503412171713751340883795768287523978524475459543415189443776886969609436705478006197723396692008709323596234752;
        data[76]<=640'd2196759186277915900926322250153512660702702110476281457737819979581075412135074665551500504044479750609692663029874974417062491293293797985828882601537181843456;
        data[77]<=640'd3734451812585640249554143841281928450105880192824227291225780984914582739891778147297281175169046805351828243620487176111287055629663337589635468384718758608896;
        data[78]<=640'd1537749138130371623117224962205775229342215845254144378050768554988013656470221484966380435991139240104230028220114544953081115824182065800004499654551648862208;
        data[79]<=640'd8786961745176465666816578199949556679295545572633687054749229839962912457951089140447432383293854575979817958002147119417324729918099622086327887568555216994304;
        data[80]<=640'd10983694272968463208017411114256965826898261436610528015286585374138212436952968448019324691735979715139294022930567373836714236557842930868698303187202758148096;
        data[81]<=640'd16695249082580503456914996506659553199402015551421791061288099602174596231441956973274026555710445567353584232040205477320890597725521914834538813215415933599744;
        data[82]<=640'd1757456916010675963431116897263003454217930426518018828788947740877615651905808648266690413449289711337892111023783134693021225513345144367168930891265539571712;
        data[83]<=640'd36026485773975688680639901527139830520404657341293837627058522077043738777291319753972334416627100670430268025266568532069969983950486661715239027820604686336000;
        data[84]<=640'd3514850144973642398087560138975016262599364512174704303161934339965326802369341883727908966006340731650767137022466249985703598557385084030274527494533533401088;
        data[85]<=640'd29875653048126526639798045376228416843826357165641766152489070646843781580116908296303110864128845455995782506093753715415935597082546797563620705583817795043328;
        data[86]<=640'd63266109313865375643071752977118740822787372271863282812817167781610080094821649312610944792567594094057266609893083522335790396888032046757915281011599004925952;
        data[87]<=640'd3514830033244166381687035798056207455250404591228774179863247277137251617984081560625554648336540389400059265172303182244137258777918140076375065009842498306048;
        data[88]<=640'd175739108367236480040979677000488704101778534884202464425131953194331274773152521036697160974466964807039099562106772512003321904383933565984467335724821647458304;
        data[89]<=640'd56236476063076019515195519781046155012777856211980571718136330521586745378286078675400513575088202484271654880263712893850577998137566993457519853062412287606784;
        data[90]<=640'd140591176749765437445189623810992435795624837489163965356149666762333898095672649144284224911363478561203128175860853594687231528725570829239145539523128057659392;
        data[91]<=640'd224945904252176205082262517795428012740351067217645091963793851838006239238882506518049539620670322340683642412762174233918148560550936107459003180443837531160576;
        data[92]<=640'd337418775931314434710666121368382058581550402986087022736596132649012604514048986252565250960473903116455606423577632442273831910856563706269486414050219291312128;
        data[93]<=640'd84354740910148374269756930822096636120398362898369227892939495922741412985713164212095828237142016513974768879467824348471207636164236838640447402853665597292544;
        data[94]<=640'd112473113019738508644751981776265581042538941086614718041905119717882505495251709234694217409485329140333609937700334099244527421821785361515272197189243978645504;
        data[95]<=640'd309300537899771631082660610980791466418600909514572953475510577119084205660416376460071170766452905968921113612060061181144695409403488757803551940537318830505984;
        data[96]<=640'd56236422431789954785131731391502193504346644638376045558492893439990743552035552631576808305257788610793059377749037847322670386405301057230994913620053708505088;
        data[97]<=640'd0;
        data[98]<=640'd0;
        data[99]<=640'd0;
        data[100]<=640'd0;
        data[101]<=640'd0;
        data[102]<=640'd0;
        data[103]<=640'd0;
        data[104]<=640'd0;
        data[105]<=640'd0;
        data[106]<=640'd0;
        data[107]<=640'd0;
        data[108]<=640'd0;
        data[109]<=640'd0;
        data[110]<=640'd0;
        data[111]<=640'd0;
        data[112]<=640'd0;
        data[113]<=640'd0;
        data[114]<=640'd0;
        data[115]<=640'd0;
        data[116]<=640'd0;
        data[117]<=640'd0;
        data[118]<=640'd0;
        data[119]<=640'd0;
        data[120]<=640'd0;
        data[121]<=640'd0;
        data[122]<=640'd0;
        data[123]<=640'd0;
        data[124]<=640'd0;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd24084754561361768648102764881807084833480156810453237320207177473645930965106688;
        data[156]<=640'd59285549689505892056868344324448208820874232148807968788202283012051522375647232;
        data[157]<=640'd70608395103938906748405107852975316393858956036050582890626880237652602651358048951934797737936631459539297024459407360;
        data[158]<=640'd1067993517960455871195206506167264853458172803453249877212770887222672897722282443732794302529536;
        data[159]<=640'd1636695303852802729735721062056679384479917375675844126961436192110104845482844076946813509129002251431657566062242728685107779566956196976088861114368;
        data[160]<=640'd1636695303852802729735721062055885040034998062974924581513017296855793489370356461447734507695151320981908907938792924355968481261496945489806448656384;
        data[161]<=640'd2864216782480733367886783702875219850681024450084810081600478838814399709490334229839490749132373384489572576545400871058621458184536325111467313463296;
        data[162]<=640'd1432108391240366683943391851438899789415357394713898207990954479728944774275910305758624481206918348577983029396480038742001836660139123208670194696192;
        data[163]<=640'd1432108391240366683943391851451811038805791937662177803850969539100631245991857707093707337766447803190049834631663961412466837165371420681761135263744;
        data[164]<=640'd1432108391240366683943391851477633537586661023558736994503006139883435319970837805366295150217217232081572022588943456326054179354432327137873574756352;
        data[165]<=640'd1432108391240366683943391851560265533685442098427726409075096037822516832042486378403564082627356928761751483328526138566416523094507341434564099702784;
        data[166]<=640'd1432108391240366683943391851436317539537270486124242286682964431933796048692382457126427995832131793975102676007502805636927351288835714611939024830464;
        data[167]<=640'd1432108391240366683943391851601596672032670643793191471755713315155913362673624275036988434856167672376313555969574319819233216692908321178052766728192;
        data[168]<=640'd1432108391240366683943391851601619368030742766333927284091709935377258825841755387755023006139996733793087972122933635263791174054830127011530100703232;
        data[169]<=640'd1432108391240366683943391851932787872881544914369532746030153642378346110315479267891213889398277586815048074848824201678868331002210464713621700083712;
        data[170]<=640'd1432108391240366683943391851439793765575186021972537001975082814418431365900148917796436548155402928625066224028133069778591550624334934584063128764416;
        data[171]<=640'd1432108391240366683943391852097696301894721300657310169440440291010802036052354946265695403268860819323901807682606887736049493626825319704900285759488;
        data[172]<=640'd1432108391240366683943391851436325104722463131847189983357910680153990639517166386655697802812652825225351447018382036542098500500671860454687275745280;
        data[173]<=640'd1432108391240366683943391852758439573882462609540164844889184258255521395328665233478876428054350936568592542451206802170221647341217223133501964943360;
        data[174]<=640'd1432108391240366683943391852758454694402165513535183429747091589205869860762080608186200982928488693054363076974248251870455480179949672581674121035776;
        data[175]<=640'd1432108391240366683943391851436347810133124628554912045016995682792950372117323359224234050582462315933974616390479971711216107968677422227345995988992;
        data[176]<=640'd1432108391240366683943391851436398293952276754886694679738749233495776634893562143924461255720267917347978930242223379402132907988712518980241656381440;
        data[177]<=640'd1432108391240366683943391852758449650944940247175441577215031711861624836036121848420102488350309449414175145035366400014318496270684891491090137350144;
        data[178]<=640'd1432108391240366683943391852097534958051516186622932203928043192673568193247427188323179442600676475226127943314644601783706513087399220109464341315584;
        data[179]<=640'd1432108391240366683943391851932916469218065658024399015447463948022914892991142494164425735624336524730464001216137266799473331018338780953464333664256;
        data[180]<=640'd1432108391240366683943391851542512683980294282207596853941880865913209292374330624151226263653084747640685832721066597117359182906917748229587519668224;
        data[181]<=640'd1432108391240366683943391851602872656675393251684714943904496310492013522598519222722702951934295630385870967567779878798513803820407135863865962659840;
        data[182]<=640'd1432108391240366683943391851467304577476394740390682301184707769031484908245125617811059271175132344711277951347270769406224545795318454304192096894976;
        data[183]<=640'd1432108391240366683943391851436317539537270486124242286683616283446132021635665278696519544222751078836949278101551891706255513177061869120807258554368;
        data[184]<=640'd1432108391240366683943391851436317539537270486124242286683225172538675800307101737124344943615829196905365418341429752739979471967507308473220046258176;
        data[185]<=640'd1432108391240366683943391851436317539537270486124242286682964431933704986088059376076228543211214608950976178501348326762462111161137601374828571394048;
        data[186]<=640'd1432108391240366683943391851436317539537270486124242286685050356773471499840398264461159746448131312586090097221999734582600997612095258161960370307072;
        data[187]<=640'd1432108391240366683943391851436317539537270486124242286703823680331370123611448259925540575580381645302115365707862404963850975670714169246146560524288;
        data[188]<=640'd1432108391240366683943391851436317539537270486124242286766401425524365536181614911473476672687882754355532927327404639568017569199443872860100527915008;
        data[189]<=640'd1432108391240366683943391851436317539537270486124242286716339229369969206125481590235127795001881867112798878031770851884684294376460109968937354002432;
        data[190]<=640'd1432108391240366683943391851436317539537270486124242286682964431933704986088059376076228543211214608950976178501348326762462111161137601374828571394048;
        data[191]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[192]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[193]<=640'd0;
        data[194]<=640'd0;
        data[195]<=640'd0;
        data[196]<=640'd0;
        data[197]<=640'd0;
        data[198]<=640'd0;
        data[199]<=640'd0;
        data[200]<=640'd0;
        data[201]<=640'd0;
        data[202]<=640'd0;
        data[203]<=640'd0;
        data[204]<=640'd0;
        data[205]<=640'd0;
        data[206]<=640'd0;
        data[207]<=640'd0;
        data[208]<=640'd0;
        data[209]<=640'd0;
        data[210]<=640'd0;
        data[211]<=640'd0;
        data[212]<=640'd0;
        data[213]<=640'd0;
        data[214]<=640'd0;
        data[215]<=640'd0;
        data[216]<=640'd0;
        data[217]<=640'd0;
        data[218]<=640'd0;
        data[219]<=640'd0;
        data[220]<=640'd0;
        data[221]<=640'd0;
        data[222]<=640'd0;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[232]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[233]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
        data[234]<=640'd716054195620183341971695925720741019646722151651777062513485227841182198836858911550944930962147952097504930445303808734511193412004703859387033190400;
        data[235]<=640'd716054195620183341971695925728810550515743740994451809925994639948462529439450235028540741451337475916307559178521450463511624135241901271801869107200;
        data[236]<=640'd613760739123428908533783747742740951106836394088668115412787031522369565600263986001412538662127949282676010716402290771643797236606065988929010532352;
        data[237]<=640'd716054195620183341971695925775162440173083066321608092275360877847400465202962165644898350748738204352527417889068168938072570349747934988601225379840;
        data[238]<=640'd716054195620183341971695925800790765867416317931110556912360783393565824159396720934922850380054260131598422539402557719009724916797066023697783980032;
        data[239]<=640'd613760739123428908533783747723284561819669846476611648565781078939270133949827327412482222507784611344649550557121527904178720485958666292289809154048;
        data[240]<=640'd717652518874151265864066222402269279027787839846796175861619257523818687142082218814817992679711572310004459761804083586737166733379098454488554405888;
        data[241]<=640'd717652518874151265864066222381610632332615704134305074641825222183666954728432874421828783111629005463041302381036565731968423454677141348080196517888;
        data[242]<=640'd717652518874151265864066222433256575542502603155916248852776122527065707065293418314348292950721787322273339470492072799817557309478448322165157658624;
        data[243]<=640'd717652518874151265864066222381611262764714851032969703153489812878113119591359665287229035812233413687691056484277674090381605018292200832336385802240;
        data[244]<=640'd717652518874151265864066222422927891246204535366129038416941852957986868373829670928928751727755942778123671315338700284483335127892308009649321279488;
        data[245]<=640'd717652518874151265864066222464243889305289847408319664706551807231782615080806708559487265778625417614943554355564108103210552528348846075417647382528;
        data[246]<=640'd717652518874151265864066222422941760753155997363957340645349445284091451629662381206239642585659882684510732393112810272150190683876353548242328223744;
        data[247]<=640'd717652518874151265864066222464262812119968119874359281204074661850797047518956100846188507001715740008955873382393081498081187779401915774669946880000;
        data[248]<=640'd717652518874151265864066222424419493636110543674992046593395335460949492590608146411639578177457561994558275334553558205843422834747255462656196214784;
        data[249]<=640'd717652518874151265864066222635639503498655084237817294316810812535102180971864697945624697763048565361384137290870518038527754274647884562071155638272;
        data[250]<=640'd717652518874151265864066222404850940396143799638307386426094989071733526486589153511271329430645730213427859000577672767480467749415025584543981633536;
        data[251]<=640'd717652518874151265864066222960034605024083301609186681386654642257410547349926520011929742823092108272697347875369729277014107534145586338041394364416;
        data[252]<=640'd717652518874151265864066222381610671811616575624536626906963505192944409669247814058411920152646564110017106347736831105814939583791750588168174305280;
        data[253]<=640'd717652518874151265864066222381610750538709446680531595425660786388142555758700960183774004641841009710024683102583580712716851135856975197608228159488;
        data[254]<=640'd717652518874151265864066222546874624761086670770212858365523676856183064079662707158119253235780059224649630232176024489037295469165907686078732566528;
        data[255]<=640'd717652518874151265864066222381610750615854520402718549706966991657617018741970816461631098917102044983181923321716996129796342907773975464120745459712;
        data[256]<=640'd615359062377396832426154045347332309252271104233890161903574413610289970352565400269832510605519953362670280927196771114792326473639327897189009588224;
        data[257]<=640'd716054195620183341971695926709742802065848854615835587395456484507104630355011217702115843703670360993952987542844175742838034909412690888906495754240;
        data[258]<=640'd716054195620183341971695926048686911771784329263129912737827550379945916191458990394396533085233974919266313840308245764022185255354348966966781280256;
        data[259]<=640'd613760739123428908533783747692296375374006368519828120208772101620735172956313190320227323430369426721036796450286682887675172004075482133507338141696;
        data[260]<=640'd716054195620183341971695927040270707349433226429013276887335984650171319874918151887948382420756493041396780925075914895627040895642094024229067423744;
        data[261]<=640'd613760739123428908533783749014408391758215345188349167726041406132073421055918000901966612090111846767563137821474696894554342628447823664269167165440;
        data[262]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[263]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[264]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[265]<=640'd0;
        data[266]<=640'd0;
        data[267]<=640'd0;
        data[268]<=640'd0;
        data[269]<=640'd0;
        data[270]<=640'd0;
        data[271]<=640'd0;
        data[272]<=640'd0;
        data[273]<=640'd0;
        data[274]<=640'd0;
        data[275]<=640'd0;
        data[276]<=640'd0;
        data[277]<=640'd0;
        data[278]<=640'd0;
        data[279]<=640'd0;
        data[280]<=640'd0;
        data[281]<=640'd0;
        data[282]<=640'd0;
        data[283]<=640'd0;
        data[284]<=640'd0;
        data[285]<=640'd0;
        data[286]<=640'd0;
        data[287]<=640'd0;
        data[288]<=640'd0;
        data[289]<=640'd0;
        data[290]<=640'd0;
        data[291]<=640'd0;
        data[292]<=640'd0;
        data[293]<=640'd0;
        data[294]<=640'd0;
        data[295]<=640'd0;
        data[296]<=640'd0;
        data[297]<=640'd0;
        data[298]<=640'd0;
        data[299]<=640'd0;
        data[300]<=640'd0;
        data[301]<=640'd0;
        data[302]<=640'd0;
        data[303]<=640'd0;
        data[304]<=640'd0;
        data[305]<=640'd0;
        data[306]<=640'd0;
        data[307]<=640'd0;
        data[308]<=640'd0;
        data[309]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[310]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[311]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[312]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[313]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[314]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[315]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[316]<=640'd716054195810719752513443498444785882909390677394503417248096665387912638568274816216319923546195994976306584519426322962481530122975535690971336409088;
        data[317]<=640'd716054195810719752513443498455645706249216138177074917164337847650413495987043420765153160381100583828079559719301877370587891032232095271147739807744;
        data[318]<=640'd716054195810719752513443498453879235507419380885030023238568209156304161116069913860135702491201439629619796773170952985848890494223452525086304632832;
        data[319]<=640'd716054195810719752513443498510497081467286048813882673100702951077881354187596314511773640630805727762155028983613816104686710516071829618063174533120;
        data[320]<=640'd716054195810719752513443498460143208844760463077529821080196447904555248326788557900137008901452003884198374928910000939410338251252270873223882604544;
        data[321]<=640'd716054195810719752513443498527281705674757012943335194389606949037152868359891240043216593653491645666403208387701926563269058460469809487764755841024;
        data[322]<=640'd716054195810719752513443498496294707137714183259419876007859178091465048512722663379328334759999833805043974433678217155421262723832670948113755668480;
        data[323]<=640'd716054195810719752513443498434320710063628340411699960038642707334417784651430246326352683510526311075218355571800711260941025649074145058756830953472;
        data[324]<=640'd716054195810719752513443498558268704211799916019206224453643091529109337873841922197184505931979417130605302723257670802630712437700647551437725761536;
        data[325]<=640'd716054195810719752513443498516952706162409451976667229383883273086102694855356451481973609612325014781178703990715379981662365375319896323895735615488;
        data[326]<=640'd716054195810719752513443498682277239580970957473452572422737403252585741964642850032475924422476581956582228806857619203036121907734186946087295647744;
        data[327]<=640'd716054195810719752513443498434744419768282745649118736482402421171162494035848669017568008616338471606971782403100048999294815896607485478661200543744;
        data[328]<=640'd716054195810719752513443498520180528360672884949629464011945630600911020862581413767102341587340635449994773464501007948977127920534674423705717702656;
        data[329]<=640'd716054195810719752513443498831341654677359009438988984845728250751230595399040954295930091273722750741024138770869931854569551962827351533791681183744;
        data[330]<=640'd716054195810719752513443498568597705571117911889023924498425831553495752160349493373008716848145533793862362408284626593044442791861272334534858244096;
        data[331]<=640'd716054195810719752513443498682216713136025199340772216790481268029865924641872019504655454319950658852344070947469645236329109806197610742822886965248;
        data[332]<=640'd716054195810719752513443498599584702262693814274499031200694035285404404923758357194094993893866283716026817139533485184985118062016148369030003032064;
        data[333]<=640'd716054195810719752513443499425904673101307019081430866693741199808277343705677208242846533457381245478574006576665460295014574276902122092042165157888;
        data[334]<=640'd716054195810719752513443498764848716623583836033777364462676998056899305882677914285810678489932238168967027307797086834675354174885748935025999478784;
        data[335]<=640'd716054195810719752513443498434320870134880584746327199572416971885421633060395155659807563156893148679265402023997279477454964846962619427443290669056;
        data[336]<=640'd716054195620183341971695925718401015768362491668746538908309926512466936160717509631240497434714115793229533898363639637246696652543009422681697157120;
        data[337]<=640'd613760739123428908533783749677723672508453639714040057671219231125749261623483559289212113580140419466065416983728004058212602728018369001831398375424;
        data[338]<=640'd716054195620183341971695927040273230619074789451038326700742560079559370057039332171767219196093483207679324237204615505148157406177362952817362337792;
        data[339]<=640'd716054195620183341971695926428277486859394827824986483955597564587821603773403629851734904263791360459596745017325418430563127492650331714001754390528;
        data[340]<=640'd716054195810719752513443502627894512384596109292216884018894224244649881100013510145154563991506566203014944728624244659254980417640361988814272462848;
        data[341]<=640'd818347651926401364867860532349971240563314498639868401812296416505884653785825610814556893644778550221301856454459734724881167850135050860994599321600;
        data[342]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[343]<=640'd0;
        data[344]<=640'd0;
        data[345]<=640'd0;
        data[346]<=640'd0;
        data[347]<=640'd0;
        data[348]<=640'd0;
        data[349]<=640'd0;
        data[350]<=640'd0;
        data[351]<=640'd0;
        data[352]<=640'd0;
        data[353]<=640'd0;
        data[354]<=640'd0;
        data[355]<=640'd0;
        data[356]<=640'd0;
        data[357]<=640'd0;
        data[358]<=640'd0;
        data[359]<=640'd0;
        data[360]<=640'd0;
        data[361]<=640'd0;
        data[362]<=640'd0;
        data[363]<=640'd0;
        data[364]<=640'd0;
        data[365]<=640'd0;
        data[366]<=640'd0;
        data[367]<=640'd0;
        data[368]<=640'd0;
        data[369]<=640'd0;
        data[370]<=640'd0;
        data[371]<=640'd0;
        data[372]<=640'd0;
        data[373]<=640'd0;
        data[374]<=640'd0;
        data[375]<=640'd0;
        data[376]<=640'd0;
        data[377]<=640'd0;
        data[378]<=640'd0;
        data[379]<=640'd0;
        data[380]<=640'd0;
        data[381]<=640'd0;
        data[382]<=640'd0;
        data[383]<=640'd0;
        data[384]<=640'd0;
        data[385]<=640'd0;
        data[386]<=640'd0;
        data[387]<=640'd0;
        data[388]<=640'd0;
        data[389]<=640'd0;
        data[390]<=640'd0;
        data[391]<=640'd0;
        data[392]<=640'd0;
        data[393]<=640'd0;
        data[394]<=640'd0;
        data[395]<=640'd0;
        data[396]<=640'd0;
        data[397]<=640'd0;
        data[398]<=640'd0;
        data[399]<=640'd0;
        data[400]<=640'd0;
        data[401]<=640'd0;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd22835963083295687686091155745995325592756551680;
        data[406]<=640'd22836137307867241909738992724944393428252229632;
        data[407]<=640'd45671926166592015614959756397608870041507332096;
        data[408]<=640'd11419593118938734974605247813455870800613605376;
        data[409]<=640'd92102251995524685136327182220460836482002714624;
        data[410]<=640'd713798081558695355229084985473875756514803712;
        data[411]<=640'd79973270849186984475343595013176781527727472640;
        data[412]<=640'd758237586915271256831821758006986185344286720;
        data[413]<=640'd188396706326222447116603965185342682481500880896;
        data[414]<=640'd10634488215193846815532761681284300800;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
    else if (choise == 2) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd0;
        data[47]<=640'd0;
        data[48]<=640'd0;
        data[49]<=640'd0;
        data[50]<=640'd0;
        data[51]<=640'd0;
        data[52]<=640'd2293498615990071511610820895302086940796564989168281123737588839386922876088484808070018553110125686554624;
        data[53]<=640'd1675976290930685468645128323187019804819274807935478584355997288644324119240316295174021690532034581474959799140168891292198173855926923755850975816974336;
        data[54]<=640'd18016743004716045104939568706166646234830913194566828459917631673408091544086843037861291450401948673299982734405370585939836303642089739931020670818844672;
        data[55]<=640'd42318397475031701438889607385923245877036691254239602651234569147285240898305566161081713485969712312403657740930550414975923248456038202051341749537734656;
        data[56]<=640'd57402183344188992557480846249111134803883445987125003633414363911957637828907724366345008656219299889741061112297913938112867822288523357300753250694201344;
        data[57]<=640'd42318407564523126557606423241263499347310989384703844829702022658899048385630712785314992999361375193054543958740802212534772278779117267377539787870175232;
        data[58]<=640'd395530360905215115021967377632711409942006648779440471063266579816800946473045629048871445053568278627989595852987097636404105016876635012054155033330057216;
        data[59]<=640'd875906954421202713545704567352562934563026676853642611817926797221644961654863567688143481820911674474299584801504605189711145700733634866251699676946366464;
        data[60]<=640'd1074300936946526427302439310125071297515937130994533697009700542908227236054607196059323136753822689742996809766773833370569381539617161493151705275232681984;
        data[61]<=640'd2723730804743768237183904232934132161590198535360849222019756894908502785821633132584250944977698014866267721515232107944067370552804837045185415225540608;
        data[62]<=640'd5363542191748007292225498426358644037797628068518507929096833266769054255422522206636867302888064784899710315832520857566929660082277303334339182503433076736;
        data[63]<=640'd3142916103311877827994774634041287214440824010129971401946070220615944633674407965106679014548230495399058990158957803742790727468293186791713320095186944;
        data[64]<=640'd11157391883955290085745718645693946645242694238428966059551126335989982129014637808743606319664413813119272322494123819208654259517587023408725019044406624256;
        data[65]<=640'd46340318392186936109177457491811105143390564853932790665686560000254254661569666650423555483369856326553091574677262891816660630792352920929528114164621377536;
        data[66]<=640'd2096606884159293981315126535532627615023078102265478175759719763157201612263761929777286175608312879866159756539412255745900722075555602617940478057775104;
        data[67]<=640'd6866055053295803659884082352104202948505894945454718108404934879957895628581040891606397478280400890069828080887171596984391567232311544567374210143564595200;
        data[68]<=640'd82380930421130208514591602192456812614175954239596008503794331118824453286272729634887977963833354862728303274743662591346725013435792896395326352926655381504;
        data[69]<=640'd123566370976313023803090396825458558807077497481013248406508153003950354552629039991956389071662517411689116159875761730931895855458626834206801549764222517248;
        data[70]<=640'd233406472398421153322362982492754957452371837391271051293079320198475871542681979470129447661822803978026991749405005742697438182615596978466919612056934023168;
        data[71]<=640'd604109837461759778168159595812365051719290138961786243677184080065183411059435054900128032160108089138751203381785997749605204012738286105816714796771764600832;
        data[72]<=640'd604113173047588382820268264222886635157617763925308602241732751467439116477112097925475867510607460983621322460590903413775070191378235877211246055920150511616;
        data[73]<=640'd219675266569980855101260213501077829681437464241079911053085166377405662230442034181704214865795090685004559815270726763607027574337217172861509719847012925440;
        data[74]<=640'd878716019124224372645561183594217863774359502483167172018946154157074302914062729473940378033073734968744706476903378722072150697136375429262006661899186339840;
        data[75]<=640'd1867228367888950619673161100430435175904078019780503412171713751340883795768287523978524475459543415189443776886969609436705478006197723396692008709323596234752;
        data[76]<=640'd2196759186277915900926322250153512660702702110476281457737819979581075412135074665551500504044479750609692663029874974417062491293293797985828882601537181843456;
        data[77]<=640'd3734451812585640249554143841281928450105880192824227291225780984914582739891778147297281175169046805351828243620487176111287055629663337589635468384718758608896;
        data[78]<=640'd1537749138130371623117224962205775229342215845254144378050768554988013656470221484966380435991139240104230028220114544953081115824182065800004499654551648862208;
        data[79]<=640'd8786961745176465666816578199949556679295545572633687054749229839962912457951089140447432383293854575979817958002147119417324729918099622086327887568555216994304;
        data[80]<=640'd10983694272968463208017411114256965826898261436610528015286585374138212436952968448019324691735979715139294022930567373836714236557842930868698303187202758148096;
        data[81]<=640'd16695249082580503456914996506659553199402015551421791061288099602174596231441956973274026555710445567353584232040205477320890597725521914834538813215415933599744;
        data[82]<=640'd1757456916010675963431116897263003454217930426518018828788947740877615651905808648266690413449289711337892111023783134693021225513345144367168930891265539571712;
        data[83]<=640'd36026485773975688680639901527139830520404657341293837627058522077043738777291319753972334416627100670430268025266568532069969983950486661715239027820604686336000;
        data[84]<=640'd3514850144973642398087560138975016262599364512174704303161934339965326802369341883727908966006340731650767137022466249985703598557385084030274527494533533401088;
        data[85]<=640'd29875653048126526639798045376228416843826357165641766152489070646843781580116908296303110864128845455995782506093753715415935597082546797563620705583817795043328;
        data[86]<=640'd63266109313865375643071752977118740822787372271863282812817167781610080094821649312610944792567594094057266609893083522335790396888032046757915281011599004925952;
        data[87]<=640'd3514830033244166381687035798056207455250404591228774179863247277137251617984081560625554648336540389400059265172303182244137258777918140076375065009842498306048;
        data[88]<=640'd175739108367236480040979677000488704101778534884202464425131953194331274773152521036697160974466964807039099562106772512003321904383933565984467335724821647458304;
        data[89]<=640'd56236476063076019515195519781046155012777856211980571718136330521586745378286078675400513575088202484271654880263712893850577998137566993457519853062412287606784;
        data[90]<=640'd140591176749765437445189623810992435795624837489163965356149666762333898095672649144284224911363478561203128175860853594687231528725570829239145539523128057659392;
        data[91]<=640'd224945904252176205082262517795428012740351067217645091963793851838006239238882506518049539620670322340683642412762174233918148560550936107459003180443837531160576;
        data[92]<=640'd337418775931314434710666121368382058581550402986087022736596132649012604514048986252565250960473903116455606423577632442273831910856563706269486414050219291312128;
        data[93]<=640'd84354740910148374269756930822096636120398362898369227892939495922741412985713164212095828237142016513974768879467824348471207636164236838640447402853665597292544;
        data[94]<=640'd112473113019738508644751981776265581042538941086614718041905119717882505495251709234694217409485329140333609937700334099244527421821785361515272197189243978645504;
        data[95]<=640'd309300537899771631082660610980791466418600909514572953475510577119084205660416376460071170766452905968921113612060061181144695409403488757803551940537318830505984;
        data[96]<=640'd56236422431789954785131731391502193504346644638376045558492893439990743552035552631576808305257788610793059377749037847322670386405301057230994913620053708505088;
        data[97]<=640'd0;
        data[98]<=640'd0;
        data[99]<=640'd0;
        data[100]<=640'd0;
        data[101]<=640'd0;
        data[102]<=640'd0;
        data[103]<=640'd0;
        data[104]<=640'd0;
        data[105]<=640'd0;
        data[106]<=640'd0;
        data[107]<=640'd0;
        data[108]<=640'd0;
        data[109]<=640'd0;
        data[110]<=640'd0;
        data[111]<=640'd0;
        data[112]<=640'd0;
        data[113]<=640'd0;
        data[114]<=640'd0;
        data[115]<=640'd0;
        data[116]<=640'd0;
        data[117]<=640'd0;
        data[118]<=640'd0;
        data[119]<=640'd0;
        data[120]<=640'd0;
        data[121]<=640'd0;
        data[122]<=640'd0;
        data[123]<=640'd0;
        data[124]<=640'd0;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd24084754561361768648102764881807084833480156810453237320207177473645930965106688;
        data[156]<=640'd59285549689505892056868344324448208820874232148807968788202283012051522375647232;
        data[157]<=640'd70608395103938906748405107852975316393858956036050582890626880237652602651358048951934797737936631459539297024459407360;
        data[158]<=640'd1067993517960455871195206506167264853458172803453249877212770887222672897722282443732794302529536;
        data[159]<=640'd1636695303852802729735721062056679384479917375675844126961436192110104845482844076946813509129002251431657566062242728685107779566956196976088861114368;
        data[160]<=640'd1636695303852802729735721062055885040034998062974924581513017296855793489370356461447734507695151320981908907938792924355968481261496945489806448656384;
        data[161]<=640'd1432108391240366683943391851438902311143753963960567794917514406880694723402274853763262205921158775538596398044052544296159347023398723736638742069248;
        data[162]<=640'd1432108391240366683943391851438899789415357394713898207990954479728944774275910305758624481206918348577983029396480038742001836660139123208670194696192;
        data[163]<=640'd1432108391240366683943391851451811038805791937662177803850969539100631245991857707093707337766447803190049834631663961412466837165371420681761135263744;
        data[164]<=640'd1432108391240366683943391851477633537586661023558736994503006139883435319970837805366295150217217232081572022588943456326054179354432327137873574756352;
        data[165]<=640'd1432108391240366683943391851560265533685442098427726409075096037822516832042486378403564082627356928761751483328526138566416523094507341434564099702784;
        data[166]<=640'd1432108391240366683943391851436317539537270486124242286682964431933796048692382457126427995832131793975102676007502805636927351288835714611939024830464;
        data[167]<=640'd1432108391240366683943391851601596672032670643793191471755713315155913362673624275036988434856167672376313555969574319819233216692908321178052766728192;
        data[168]<=640'd1432108391240366683943391851601619368030742766333927284091709935377258825841755387755023006139996733793087972122933635263791174054830127011530100703232;
        data[169]<=640'd1432108391240366683943391851932787872881544914369532746030153642378346110315479267891213889398277586815048074848824201678868331002210464713621700083712;
        data[170]<=640'd1432108391240366683943391851439793765575186021972537001975082814418431365900148917796436548155402928625066224028133069778591550624334934584063128764416;
        data[171]<=640'd1432108391240366683943391852097696301894721300657310169440440291010802036052354946265695403268860819323901807682606887736049493626825319704900285759488;
        data[172]<=640'd1432108391240366683943391851436325104722463131847189983357910680153990639517166386655697802812652825225351447018382036542098500500671860454687275745280;
        data[173]<=640'd1432108391240366683943391852758439573882462609540164844889184258255521395328665233478876428054350936568592542451206802170221647341217223133501964943360;
        data[174]<=640'd1432108391240366683943391852758454694402165513535183429747091589205869860762080608186200982928488693054363076974248251870455480179949672581674121035776;
        data[175]<=640'd1432108391240366683943391851436347810133124628554912045016995682792950372117323359224234050582462315933974616390479971711216107968677422227345995988992;
        data[176]<=640'd1432108391240366683943391851436398293952276754886694679738749233495776634893562143924461255720267917347978930242223379402132907988712518980241656381440;
        data[177]<=640'd1432108391240366683943391852758449650944940247175441577215031711861624836036121848420102488350309449414175145035366400014318496270684891491090137350144;
        data[178]<=640'd1432108391240366683943391852097534958051516186622932203928043192673568193247427188323179442600676475226127943314644601783706513087399220109464341315584;
        data[179]<=640'd1432108391240366683943391851932916469218065658024399015447463948022914892991142494164425735624336524730464001216137266799473331018338780953464333664256;
        data[180]<=640'd1432108391240366683943391851542512683980294282207596853941880865913209292374330624151226263653084747640685832721066597117359182906917748229587519668224;
        data[181]<=640'd1432108391240366683943391851602872656675393251684714943904496310492013522598519222722702951934295630385870967567779878798513803820407135863865962659840;
        data[182]<=640'd1432108391240366683943391851467304577476394740390682301184707769031484908245125617811059271175132344711277951347270769406224545795318454304192096894976;
        data[183]<=640'd1432108391240366683943391851436317539537270486124242286683616283446132021635665278696519544222751078836949278101551891706255513177061869120807258554368;
        data[184]<=640'd1432108391240366683943391851436317539537270486124242286683225172538675800307101737124344943615829196905365418341429752739979471967507308473220046258176;
        data[185]<=640'd1432108391240366683943391851436317539537270486124242286682964431933704986088059376076228543211214608950976178501348326762462111161137601374828571394048;
        data[186]<=640'd1432108391240366683943391851436317539537270486124242286685050356773471499840398264461159746448131312586090097221999734582600997612095258161960370307072;
        data[187]<=640'd1432108391240366683943391851436317539537270486124242286703823680331370123611448259925540575580381645302115365707862404963850975670714169246146560524288;
        data[188]<=640'd1432108391240366683943391851436317539537270486124242286766401425524365536181614911473476672687882754355532927327404639568017569199443872860100527915008;
        data[189]<=640'd1432108391240366683943391851436317539537270486124242286716339229369969206125481590235127795001881867112798878031770851884684294376460109968937354002432;
        data[190]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[191]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[192]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[193]<=640'd0;
        data[194]<=640'd0;
        data[195]<=640'd0;
        data[196]<=640'd0;
        data[197]<=640'd0;
        data[198]<=640'd0;
        data[199]<=640'd0;
        data[200]<=640'd0;
        data[201]<=640'd0;
        data[202]<=640'd0;
        data[203]<=640'd0;
        data[204]<=640'd0;
        data[205]<=640'd0;
        data[206]<=640'd0;
        data[207]<=640'd0;
        data[208]<=640'd0;
        data[209]<=640'd0;
        data[210]<=640'd0;
        data[211]<=640'd0;
        data[212]<=640'd0;
        data[213]<=640'd0;
        data[214]<=640'd0;
        data[215]<=640'd0;
        data[216]<=640'd0;
        data[217]<=640'd0;
        data[218]<=640'd0;
        data[219]<=640'd0;
        data[220]<=640'd0;
        data[221]<=640'd0;
        data[222]<=640'd0;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[232]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[233]<=640'd818347651926401364867860531033023802736586063526677795500824789374085118993324709360679195491452077832178144388559175842876329562291030954944736788480;
        data[234]<=640'd716054195620183341971695925720741019646722151651777062513485227841182198836858911550944930962147952097504930445303808734511193412004703859387033190400;
        data[235]<=640'd716054195620183341971695925728810550515743740994451809925994639948462529439450235028540741451337475916307559178521450463511624135241901271801869107200;
        data[236]<=640'd613760739123428908533783747742740951106836394088668115412787031522369565600263986001412538662127949282676010716402290771643797236606065988929010532352;
        data[237]<=640'd716054195620183341971695925775162440173083066321608092275360877847400465202962165644898350748738204352527417889068168938072570349747934988601225379840;
        data[238]<=640'd613760739123428908533783747774928292360646253992264782241007928140561643021750641094820659994869755220633213660416305499971685649738147490781267492864;
        data[239]<=640'd613760739123428908533783747723284561819669846476611648565781078939270133949827327412482222507784611344649550557121527904178720485958666292289809154048;
        data[240]<=640'd716054195620183341971695925738817416463807378774612244561406621609641403574405348038827264337467752714227304585783342624856277106966463240300037931008;
        data[241]<=640'd716054195620183341971695925718158769768635243062121143341612586269489671160756003645838054769385185867264147205015824770087533828264506133891680043008;
        data[242]<=640'd716054195620183341971695925769804712978522142083732317552563486612888423497616547538357564608477967726496184294471331837936667683065813107976641183744;
        data[243]<=640'd716054195620183341971695925718159400200734389960785771853277176963935836023682794511238307469989594091913901308256933128500715391879565618147869327360;
        data[244]<=640'd716054195620183341971695925759476028682224074293945107116729217043809584806152800152938023385512123182346516139317959322602445501479672795460804804608;
        data[245]<=640'd716054195620183341971695925800792026741309386336135733406339171317605331513129837783496537436381598019166399179543367141329662901936210861229130907648;
        data[246]<=640'd716054195620183341971695925759489898189175536291773409345136809369914168061985510430248914243416063088733577217092069310269301057463718334053811748864;
        data[247]<=640'd716054195620183341971695925800810949555987658802175349903862025936619763951279230070197778659471920413178718206372340536200298152989280560481430405120;
        data[248]<=640'd716054195620183341971695925760967631072130082602808115293182699546772209022931275635648849835213742398781120158532817243962533208334620248467679739904;
        data[249]<=640'd716054195620183341971695925972187640934674623165633363016598176620924897404187827169633969420804745765606982114849777076646864648235249347882639163392;
        data[250]<=640'd716054195620183341971695925741399077832163338566123455125882353157556242918912282735280601088401910617650703824556931805599578123002390370355465158656;
        data[251]<=640'd716054195620183341971695926296582742460102840537002750086442006343233263782249649235939014480848288676920192699348988315133217907732951123852877889536;
        data[252]<=640'd716054195620183341971695925718158809247636114552352695606750869278767126101570943282421191810402744514239951171716090143934049957379115373979657830400;
        data[253]<=640'd716054195620183341971695925718158887974728985608347664125448150473965272191024089407783276299597190114247527926562839750835961509444339983419711684608;
        data[254]<=640'd716054195620183341971695925883422762197106209698028927065311040942005780511985836382128524893536239628872475056155283527156405842753272471890216091648;
        data[255]<=640'd716054195620183341971695925718158888051874059330534618406754355743439735174293945685640370574858225387404768145696255167915453281361340249932228984832;
        data[256]<=640'd613760739123428908533783748683880446688290643161706230603361777696112686784888529493841782263276133766893125751176030152911436847226692683000493113344;
        data[257]<=640'd613760739123428908533783748683880328559078790676989812724103629254100449217365137862013653318485856082987778663857923523799995642353772355989979267072;
        data[258]<=640'd716054195620183341971695926048686911771784329263129912737827550379945916191458990394396533085233974919266313840308245764022185255354348966966781280256;
        data[259]<=640'd613760739123428908533783747692296375374006368519828120208772101620735172956313190320227323430369426721036796450286682887675172004075482133507338141696;
        data[260]<=640'd716054195620183341971695927040270707349433226429013276887335984650171319874918151887948382420756493041396780925075914895627040895642094024229067423744;
        data[261]<=640'd716054195620183341971695927040270865264985409127194942397394261385077602193564080742068802475296351678528346700460949113592381895506742197185683652608;
        data[262]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[263]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[264]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[265]<=640'd0;
        data[266]<=640'd0;
        data[267]<=640'd0;
        data[268]<=640'd0;
        data[269]<=640'd0;
        data[270]<=640'd0;
        data[271]<=640'd0;
        data[272]<=640'd0;
        data[273]<=640'd0;
        data[274]<=640'd0;
        data[275]<=640'd0;
        data[276]<=640'd0;
        data[277]<=640'd0;
        data[278]<=640'd0;
        data[279]<=640'd0;
        data[280]<=640'd0;
        data[281]<=640'd0;
        data[282]<=640'd0;
        data[283]<=640'd0;
        data[284]<=640'd0;
        data[285]<=640'd0;
        data[286]<=640'd0;
        data[287]<=640'd0;
        data[288]<=640'd0;
        data[289]<=640'd0;
        data[290]<=640'd0;
        data[291]<=640'd0;
        data[292]<=640'd0;
        data[293]<=640'd0;
        data[294]<=640'd0;
        data[295]<=640'd0;
        data[296]<=640'd0;
        data[297]<=640'd0;
        data[298]<=640'd0;
        data[299]<=640'd0;
        data[300]<=640'd0;
        data[301]<=640'd0;
        data[302]<=640'd0;
        data[303]<=640'd0;
        data[304]<=640'd0;
        data[305]<=640'd0;
        data[306]<=640'd0;
        data[307]<=640'd0;
        data[308]<=640'd0;
        data[309]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[310]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[311]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[312]<=640'd613760739313965319075531320408458236556858239776876329526145666308279278680393113741210666432843826362831716502048441626146057261718376763829329592320;
        data[313]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[314]<=640'd613760739313965319075531320408458236556858239776876329526145666308279278680393113741210666432843826362831716502048441626146057261718376763829329592320;
        data[315]<=640'd613760739313965319075531320408458236556858239776876329526145666308279278680393113741210666432843826362831716502048441626146057261718376763829329592320;
        data[316]<=640'd716054195810719752513443498444785882909390677394503417248096665387912638568274816216319923546195994976306584519426322962481530122975535690971336409088;
        data[317]<=640'd615359062377396832426154044377073155011433474656812112937181322717155631643064706157843113125738871714582669885975835649477700443377317343088179412992;
        data[318]<=640'd717652518874151265864066222401169157776406781303612993682764539476050477909737279092927845621024232427088115818831163483776739172427593129943260725248;
        data[319]<=640'd615359062377396832426154044431924530229503385293619868873546426144623489843617599904463593375444015648658139150287774383576519927217051690003614138368;
        data[320]<=640'd717652518874151265864066222407433131113747863496112791524392778224301565120455923132929152031274796681666693974570211437338186929456411478080838696960;
        data[321]<=640'd717652518874151265864066222474571627943744413361918164833803279356899185153558605276008736783314438463871527433362137061196907138673950092621711933440;
        data[322]<=640'd717652518874151265864066222443584629406701583678002846452055508411211365306390028612120477889822626602512293479338427653349111402036811552970711760896;
        data[323]<=640'd717652518874151265864066222381610632332615740830282930482839037654164101445097611559144826640349103872686674617460921758868874327278285663613787045888;
        data[324]<=640'd717652518874151265864066222505558626480787316437789194897839421848855654667509287429976649061802209928073621768917881300558561115904788156294681853952;
        data[325]<=640'd717652518874151265864066222464242628431396852395250199828079603405849011649023816714765752742147807578647023036375590479590214053524036928752691707904;
        data[326]<=640'd717652518874151265864066222629567161849958357892035542866933733572332058758310215265268067552299374754050547852517829700963970585938327550944251740160;
        data[327]<=640'd717652518874151265864066222382034342037270146067701706926598751490908810829516034250360151746161264404440101448760259497222664574811626083518156636160;
        data[328]<=640'd717652518874151265864066222467470450629660285368212434456141960920657337656248778999894484717163428247463092510161218446904976598738815028562673795072;
        data[329]<=640'd717652518874151265864066222778631576946346409857571955289924581070976912192708319528722234403545543538492457816530142352497400641031492138648637276160;
        data[330]<=640'd717652518874151265864066222515887627840105312307606894942622161873242068954016858605800859977968326591330681453944837090972291470065412939391814336512;
        data[331]<=640'd615359062377396832426154044603644161898242535820509412563324743096608060297893304897345407064588946738847181114143603515218919217342832814763326570496;
        data[332]<=640'd717652518874151265864066222546874624531681214693082001644890365605150721717425722426887137023689076513495136185193695682912966740220288973886959124480;
        data[333]<=640'd716853363439600646524677188316731723675578660205953099308361143989941438870815068241597331819765499423190922271032540390475808958676019893080575442944;
        data[334]<=640'd716054195810719752513443498764848716623583836033777364462676998056899305882677914285810678489932238168967027307797086834675354174885748935025999478784;
        data[335]<=640'd716054195810719752513443498434320870134880584746327199572416971885421633060395155659807563156893148679265402023997279477454964846962619427443290669056;
        data[336]<=640'd716054195810719752513443498434562956063355552322347499764326232106897902934727015174439082647135142591538370028724170101199737600751504032013257539584;
        data[337]<=640'd716054195810719752513443500419748086310216764306486793198588391973184409535139144672512889177745951175339461993074786741203682943285782144079475245056;
        data[338]<=640'd716054195810719752513443499756435170914067850104639287556758865673990336831048837714965804408514510005988160367565145969101198354385857562148922720256;
        data[339]<=640'd716054195810719752513443499144439427154387888478587444811613870182252570547413135394933489476212387257905581147685948894516168440858826323333314772992;
        data[340]<=640'd818347651926401364867860535221433105301380051923860736978214468308792128689640578898859583951849017517362481346889435950386937788282291303067668185088;
        data[341]<=640'd1636695303852802729735721063377830543543726744987234358969115182131310361193491873149574770423149332809446318453759619861197221749554275471993841123328;
        data[342]<=640'd1636695303852802729735721062055718605960824492694731914313637531250851414815332524670035753556741565176288923998599770272632107798838449221998483603456;
        data[343]<=640'd0;
        data[344]<=640'd0;
        data[345]<=640'd0;
        data[346]<=640'd0;
        data[347]<=640'd0;
        data[348]<=640'd0;
        data[349]<=640'd0;
        data[350]<=640'd0;
        data[351]<=640'd0;
        data[352]<=640'd0;
        data[353]<=640'd0;
        data[354]<=640'd0;
        data[355]<=640'd0;
        data[356]<=640'd0;
        data[357]<=640'd0;
        data[358]<=640'd0;
        data[359]<=640'd0;
        data[360]<=640'd0;
        data[361]<=640'd0;
        data[362]<=640'd0;
        data[363]<=640'd0;
        data[364]<=640'd0;
        data[365]<=640'd0;
        data[366]<=640'd0;
        data[367]<=640'd0;
        data[368]<=640'd0;
        data[369]<=640'd0;
        data[370]<=640'd0;
        data[371]<=640'd0;
        data[372]<=640'd0;
        data[373]<=640'd0;
        data[374]<=640'd0;
        data[375]<=640'd0;
        data[376]<=640'd0;
        data[377]<=640'd0;
        data[378]<=640'd0;
        data[379]<=640'd0;
        data[380]<=640'd0;
        data[381]<=640'd0;
        data[382]<=640'd0;
        data[383]<=640'd0;
        data[384]<=640'd0;
        data[385]<=640'd0;
        data[386]<=640'd0;
        data[387]<=640'd0;
        data[388]<=640'd0;
        data[389]<=640'd0;
        data[390]<=640'd0;
        data[391]<=640'd0;
        data[392]<=640'd0;
        data[393]<=640'd0;
        data[394]<=640'd0;
        data[395]<=640'd0;
        data[396]<=640'd0;
        data[397]<=640'd0;
        data[398]<=640'd0;
        data[399]<=640'd0;
        data[400]<=640'd0;
        data[401]<=640'd0;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd22835963083295687686091155745995325592756551680;
        data[406]<=640'd22836137307867241909738992724944393428252229632;
        data[407]<=640'd45671926166592015614959756397608870041507332096;
        data[408]<=640'd11419593118938734974605247813455870800613605376;
        data[409]<=640'd92102251995524685136327182220460836482002714624;
        data[410]<=640'd713798081558695355229084985473875756514803712;
        data[411]<=640'd79973270849186984475343595013176781527727472640;
        data[412]<=640'd758237586915271256831821758006986185344286720;
        data[413]<=640'd188396706326222447116603965185342682481500880896;
        data[414]<=640'd10634488215193846815532761681284300800;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
    else if(choise == 3) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd431895724276146852830977159046070056467417078723387852467328750087181887064079715333668321043822420951087286941007451361404270074957102972420397963508726311564607488;
        data[47]<=640'd228497919586486263430877312029699219911028689096061489821504387260523976261328252787616651596956943661478685623854851516667697908800149485002736051972102815534821670912;
        data[48]<=640'd3773660090784995245506048679358193937811722789130580324090229290824194936866332802975318672096147353141206667372181560078356365898369527320639908893727530004470120316928;
        data[49]<=640'd7547806062502412955509311931052063658436180718616534579248465686246563531523429294171109087756701207588969498169221879910342223094913524639101725396896223259012240506880;
        data[50]<=640'd105669105129368583765200805132790894110951482840784741636629989946058911401059457603857049857906491500160214585931049581742287987220469106067475412093818047345919583584256;
        data[51]<=640'd241533356631917302690906770287657974446474315656264739503185543366548765200272019911819594284289656929694019574690764758319537106631132137284634939925881957629936204251136;
        data[52]<=640'd966134377139367056742601970207836612350912729461288549725173816585962162113359512199166195621366615918867166138004553222846953810310247277975662400427372215038838501801984;
        data[53]<=640'd3592810253839269060329853827044096611354510445561682323474351637255952848030289787753998887421881375269547898336374926991627263586395381050227324975361281861425225736912896;
        data[54]<=640'd7649820913732204422183487345775079170323264499427987117051315817983495420076536051203043107048824255595630334571926459425407591426698906795308954576219656180896290708652032;
        data[55]<=640'd14492013882938578808340826175769905664467702354322723609858706877540699561609022877596506853084439416827633523896740310854898406783807780709954342704272744107339718699515904;
        data[56]<=640'd29215894239259061193887916129795074451736415815720894414412949946219634118487290491755984718688305207927398346822633353273829670383514238354821614792669603136420308148289536;
        data[57]<=640'd53437420954267644330077737259441538062396207039972045300882505515343843234042718199046995071057399754736395529406121560634332073310071398793146837024928794141927330390474752;
        data[58]<=640'd121729158012618816317388870684855874176710613959469966170525893549682196552955761694758139901475754017952978293215031561539679958120639968110391918380547592531893747347095552;
        data[59]<=640'd118698666185487118611067892135882898410314166492812507845277677840957483040379946689930537446739086773873335251787467418237820707097552450025674088275590776891097391910879232;
        data[60]<=640'd208654834543533378284406841078015218160909833642051580505137921711961107846991481044157714394608698999098644588591417014853589196686802904417552019167720156965257506874982400;
        data[61]<=640'd848205602903491062002232486018965500899495478789979628485906118656341371162268408440616666069843272495741337853937142678774421849146349639218321173181920487901262305298481152;
        data[62]<=640'd958043005315497201517452105720061935001731770549357881767474838964552506860821746704059596022140393134755192998773528916600338066421400280308421417976973221116390909511991296;
        data[63]<=640'd1977918610999270536546640245720557131404918110283328844545414243853225816582046841609763260179927978610694576783729993001589177783102950416020337908700065323115452177999462400;
        data[64]<=640'd3925403989004780163630953576234107919140139392872598245592575974021993352483204386795659637219369769904719371173170347912559877971984612208159146606597801168149298115948576768;
        data[65]<=640'd1479151736934855631441674776313804205993809976005043141803966916015739517100602592165219563684691791107819863694345806604082036278019522465225871186714418441600200934009339904;
        data[66]<=640'd6905928553631840661983160375639174958612744938799899871182102249836751342034532810995435275398715617037410380623948506354084127761813144801921955907919087220795397293505249280;
        data[67]<=640'd3951489617285146657476130401565383827313510164257655629668092529572278260916339177755573602934181827055725256196162672953640933999920685850545039702993779948738223377953587200;
        data[68]<=640'd7416047506670118763493366027547130612271216425796493530416825005331807350133988631017988693884709624974328249077724049807172184563102337929187552350657427625626431642897743872;
        data[69]<=640'd15825281156755672921540638117172662345010730729519976133903577002311254085615950741699313879295846421335214742818419488673686298295338113851749603355218438328529778508220596224;
        data[70]<=640'd7651784295574171522547036743095324974743687666684562912586656018669134170469538057434590120099930567410282378557205632648550565261984016522514842335984316056656534007913119744;
        data[71]<=640'd31155901510565136774953606569028353669882164698110672714742077448413667404270616385693110185335694847602542971962784845748360069375165792342188656650947038735677235561645473792;
        data[72]<=640'd27677817739849604264761715287449800625998820148068332392033276285142366527453396383664157493173501088838999138832619652159062061450890597365106564562376021668577651219190775808;
        data[73]<=640'd31642833238465311326419146327546019627108145368451807038127325214763466635390644732879416060406053953086557721617179952167089377331934575260326378616938572464972032765794975744;
        data[74]<=640'd31642833238465311326419146327546019640423836475974858832416293796129820654321768726153154928511135458798122188617703024411647539510338426892890131038031749603349359600628400128;
        data[75]<=640'd59282005603084743007733934283211363510875399067120394885539873257429223299320411056718993796648627596311573606241394912114998379629234621901641409507445839146657482953841442816;
        data[76]<=640'd63285666476930622652811477039232154039119072846746146287204814275214521403742110673700403122085003548091753712635459483621258166202391551099576848730669839320366984145649270784;
        data[77]<=640'd62791005673984413584663656381332974436287810422295569935568206299122032115431078493421960782961983523059985844011318710819394458408385505433696637697235055750676965534241652736;
        data[78]<=640'd62791005673984413584717287613052744829477424559176606551105300217302326825448214073045959408935046526815650429727445302447421975644432387717050829727116471051599295066237042688;
        data[79]<=640'd62296344871038204516596282571013450452407554954080214895180147103148440397720739658936550450197909687805643698670419135605327993933651443415948137734708554556807773766457229312;
        data[80]<=640'd126602249254045383372434200499561260636873002409056063669366762258373524759171571023429616942634132554603031534766565156522868929900629354827762248134792291893549553467246247936;
        data[81]<=640'd126602249254045383372273306804401949467212416987005384780301806784837730601653266650403154247390182326224649597285794882946953075377593263961600581472220569048216986830612987904;
        data[82]<=640'd126602249254045383372434200499561260635332092956694309942544687944834895655524113487948122135145564486430645020123767406354237472563271036449149645680848137779969622379344166912;
        data[83]<=640'd126478584056533652073931830926171238897674893174786800105671732550485414019318290988073135137506231396128856285554140720395433496595307245899799983636752848682067193593195397120;
        data[84]<=640'd126571332957546754827145848788693665246823609350605921389340569650831134715317250858968384295739554069591134424940416213181573176478403141481088731836253413212298988404799963136;
        data[85]<=640'd126540416657362616980008179866025949835765724888107371395408014035248195668751343014615044314169932339393068281088196884380491780514114789648508336243590585026022912525212844032;
        data[86]<=640'd126571332957431583073245330746213196429465489082187721456207428211896699424965281297427064696054676378709662249881878694390204197958689446813231350308253094396984909773840318464;
        data[87]<=640'd126602249257615721140110156024780193118268196322168524533712204559983171081501491415286839257134734108577275777838226135892538031549875846099019291710457505941208335432944713728;
        data[88]<=640'd126602249257268404995158013456097276948654364889367557556593612402299761092895760172415283505057184266879906044230760052942304271144870345434394093585331184852339857207261659136;
        data[89]<=640'd126540416656425943347711442735024076986627693013555633244848371990972755747694667702453652183223335331768828782603269153583451097234751763537544517954066984109661194971061944320;
        data[90]<=640'd126416751456622465801535372325009733102666032800512861849771616385649780975724159850825512234869049264928879344484476777976501661707980435853102056746626753870103911371653513216;
        data[91]<=640'd126602249257261206733046520918094952295836386278536119744242297966425221032613894207143430669638078654361646169891712025333249012847457352825566964591853059224083062645323726848;
        data[92]<=640'd63285666476931072324544221850550809386978023378066366271925014424145408903196997012712271729221272497858833962919743886006791371129558999636545859647816394320817239470116962304;
        data[93]<=640'd63285666476931072324544221850550809375092750879957068838235239807470238158128827681977147192020087052290421933672252042618874884425132430237783140743011969422341928763695038464;
        data[94]<=640'd63285666476931072324490590618831039010325441062690550238693767940209533855903997361238504943378167746823333318143589097778147299694205406730079784456631448892637529208935940096;
        data[95]<=640'd63301124627023141357896213829379515335131335624147397085171828143257410095823704386495809514062016206146474841378800427786240890670102853090712226029407139142057139950812397568;
        data[96]<=640'd31519168037729208731148455494214736609804481573476891197649410955265077715714401473995960428971984473257069829563434622872270729675060358208287887760280253467026236709812568064;
        data[97]<=640'd44998674918013405837419027273925623272519992049496524780711176907857102831894180904457417898692046729169078143609453909607890095990457628390334937405104768998483696403137691648;
        data[98]<=640'd31395502836992656464051165194055200076899881052553389466458423277717996337024683256855118701153011706602439833352571648645034148768432836422724791467706144117307270285265731584;
        data[99]<=640'd27198615086995913901725407754870572833453566267799342958925485173146129293935855067328488502505244765846444796631760641478518728498293099694556621240360132118853449794141028352;
        data[100]<=640'd31619646013327657448056903411659197939992054542452129589781840297658207566940465428998427596362614407444272268322162778996334867952670114603026624942404676680592359122362433536;
        data[101]<=640'd15798229394095001784874145863746073336883431910119140066127143141187660693123751627630843152888457839422020809304253191434675072353859769438468277311757035448014700760174428160;
        data[102]<=640'd10874808589771014653705451938838836361362170550705333757888238189453049211479931635065136345344705857141882437499900750305185321837458999063203895931666048256762663280744333312;
        data[103]<=640'd5769754521865216380362898637698896871873545256363282738512972082763743225613311263739662508339727690040653828307797938017267117426161092888259372262827217318188642234234044416;
        data[104]<=640'd7769652690026647573742743241256200513038132968862885331335847038594302372591037953856698519134502829734705401049021300427915253371611742820767175443796238981860907695002877952;
        data[105]<=640'd7874961337528867863620506321254066960081023257501424885859449861743464678094133477815848848496456939330418200207230968766567674646348879069289749570467994586884469040147857408;
        data[106]<=640'd2966998683296949765855627058584443967157939169850647300119054777564191360930437226828924358523544188314345311516764693105917656058517330512061872607787782630060539350611918848;
        data[107]<=640'd1976227875833400157731112287454330637030825029794083244997833394528890664901189381461884847573927659455077067303295088856073225171768517546758269718810474084311833160703803392;
        data[108]<=640'd1938790168579170467516772135859127057923884524428214636761214199970207494036936097643775194948157308964066500543821265811757781066917144841677677016187269656120312787596476416;
        data[109]<=640'd1961132026134113992318467596434754249526173344394813507800210508082198174036873398682888933816695358056976779992570434298494108344146716834121085160365274794475927463882915840;
        data[110]<=640'd989261222494070663287455238984222672121013582736623018089736540737356846300182373166424243505308617797634803289080693980388415640431005444094012314438668335800673618783895552;
        data[111]<=640'd366617805797313484829757829024441114258431376416569845995500673404339346531022996004734655986235912394523801362535374162115296964602789352319164306631950813734283144268349440;
        data[112]<=640'd494019229334439077797891110068214099902240231834475355251103587337617530316113364674530295863580538952667893709263193246592685178263104004433665817599049950592467867099201536;
        data[113]<=640'd237357705765963282743521867899250866735100828129793758052614961003313975840699763347526313906691439099217306524113814493465796448486374286930965424471058839165493092512956416;
        data[114]<=640'd119769528023979902675728407366609004777665787500497614308024478563915750091105575718802645279546984625475279053341035689075854751037462751001851043070950415967736919069032448;
        data[115]<=640'd30795327003372146886382952461496954673372391357243188361171041565846513733671961650171624728332181429344103634740328647090679507241346455035560987379483451762077364324925440;
        data[116]<=640'd28433032833023521126034322674569664848413929464020181414594708767492302302573599812484485691771471276409848479283811882698866517325118065980436035960197046481291110902661120;
        data[117]<=640'd11593612453879362220307475021310777717673832905471827687771032501840939053910346491860523655214459956208420838520213833743296652255574059602367796998186049072833919839109120;
        data[118]<=640'd3856753667929747671988133972783950575043030316210607873116383978798874578957560354248322958924866582502398611001229264552479476372206780112683678734613823369773353829138432;
        data[119]<=640'd1807551097000635124452604227822980692803309903755754272045843150551132787369237451409171873697570621390911703659822243592899726602739554744376689780314199485672380098936832;
        data[120]<=640'd482933588832450652885872289239547593210678889708833741568178514263710791452042372209198001912354457299585096204321159691864132439358227953102114004872640732631303173701632;
        data[121]<=640'd120527001888151747069384576324811300420641789837885846323457162580513971964969372133823588886123014259339317412883678691848571564732031817092699540859705618827924329201664;
        data[122]<=640'd11319464145435777483299695034266588835712935291767801343756229713115700839390244132624242621946020889747090827523526725945383644196322512132176324978665043635069914185728;
        data[123]<=640'd941352272478838956829228612731650408937000358393345031289481611054277775067553879797107795145511842378094999342368103878040169316019492455665379934689717719187931004928;
        data[124]<=640'd6795159395278043816784342275027866533519695616054367924460808287983682664866521938369622172405271328050352938991837858742519764757852736816089139692116332862144249856;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd0;
        data[156]<=640'd0;
        data[157]<=640'd0;
        data[158]<=640'd0;
        data[159]<=640'd0;
        data[160]<=640'd0;
        data[161]<=640'd0;
        data[162]<=640'd0;
        data[163]<=640'd0;
        data[164]<=640'd0;
        data[165]<=640'd0;
        data[166]<=640'd2404907604760405225358828131112281116032698930082119547604265954848982041717359046106827774346003151904701415424;
        data[167]<=640'd225966000196679199302367116694592893265725867803609040642871570818141414006515693128818279001101907621668191107533366624180671486377020044585858807471037437053672466939904;
        data[168]<=640'd233749797701388404744170545964817196039464493250426943775204130042126013255833596973025305736092108424206759168945283235326066943996789563483062887518151008876675286958080;
        data[169]<=640'd222427910426923780687445880271616953451946654688046958211095861131545676237587670576040436326739951765773448355932093025124234101847461544073800682614313097394758124306432;
        data[170]<=640'd482005763459180421821310258297570210540068800232038071206407166154550177157033106626446922038581023496705391989992117930938841859872661048742389427527021643153693388832768;
        data[171]<=640'd208865232962721366452827594859695917982739058486193301478069737090979754636560327097379632204909018590485181723438140771027562820836956585082585480465233489063548305801216;
        data[172]<=640'd300855567067746436913715538099334253109316714190688122113675802432638508779745111736786506815949964456156477130050019191842205490052930653685084556541795330863298097709056;
        data[173]<=640'd694114245366728613134011418019667609488335496250869617457894284200595130941349212228783727810149791613467693471655361366132132768788137053348604374707072101221132828409856;
        data[174]<=640'd775490310151943098541719551645524320252412922690017776067063500966114909387262974014165621074406022099779893233530142173927865550274575091592966918519011498276665287507968;
        data[175]<=640'd894370126533821651137328520943796744158169727542393221243297899005725777707576051286859293751919023315188737088962168045529823492091638066674721046381892945249715114475520;
        data[176]<=640'd1919000924872870128270910589688399449589991508785090142993182266482543276251070558587164243705154721956701603660157920890701387724415865765316699923833493507388896230506496;
        data[177]<=640'd1905762572304550815246250761509776537621071996066598098008691595853692639432717375412344483305018624665089328675040739680193539225472186731449663940338362953374872033558528;
        data[178]<=640'd909259587663000388503594029257889725314743063194450806094635784345810604609139915003456009165329215073900514085279304993254393134484803582428583682857324591906586923892736;
        data[179]<=640'd1903344877626149515317471015606330927862828343409768818410542987349595860003824861623343385568601502771991516052754801276251192881198773901076232652089855637643885348388864;
        data[180]<=640'd3805893685039309049516244718747041982496321253652206854350051770736069707885845870042035147901523896362096737568733904804694300801402997975640890585727348634533742818361344;
        data[181]<=640'd3685259565811517358557679714308655246815176072610536026165225277001635817227135304339210642111048471921136359436174812095720825141994293452586494268791592200161347179118592;
        data[182]<=640'd3806026363405806681829409460900279851324517551663862128265891197911721682345412046792081609111580956092035657234511293236504417678616436176705904033348700167097010066817024;
        data[183]<=640'd6703493386082906034585816587240314285038661390750342894509211492702915988179088836301168574105405025853047923932209313306770466737423895439526932493080467841967723064066048;
        data[184]<=640'd5495353664836910109199488927001444706333793259629029588707057977503463613187997297548528271411153582170721866787360326580665432530827264402522893337552689495647960745115648;
        data[185]<=640'd6159924860582828406695775178997347681343783581218932178664071698982813324680761503518299746381415565073788251480791862646724033775004819293767296608772914596609984213024768;
        data[186]<=640'd15096303017052369839942573385856164275755916153892502817789395624331301478631009149703006214269475340313246437181101306077572458561590363835121544294235439741162021166514176;
        data[187]<=640'd14854692026150000907883101126416859643255715746356198663961015507162334475663146251842362767614409241851642098236651323140807703771564959397674207621339961363719224641454080;
        data[188]<=640'd15337851354281670445631940072611995470201196412240349960395597427291191473717551487447710929681899572343003061891258572336783746486555067543930172465538442230615465688825856;
        data[189]<=640'd22946041666396122138583656559303689670887134615101069331168908759921366635491055857782241569695026514453998880600165378899374929766716690643426637474391759412729786325270528;
        data[190]<=640'd30674996933349772909913864393390435727903224561494786881319545254346462599238459890180980900845314732669751989351468000727323570306008548726279699238625697289411972491640832;
        data[191]<=640'd30675000618859953399700341191783581224260494964599621455789046420900018349101769312767244846593145445877099102554203071614132585149170931123074909513783838011170549489729536;
        data[192]<=640'd30433452281630652794010974505027750029816456862280028973620319516976968350758774023511735582612645791476705497074579820710164648750002865205445228893419953564025198481506304;
        data[193]<=640'd22704274041311082390598920368155701443241071830584788016371884909038331324788035981174452942043244744388123211969656376107140881052462333404407696783681047190526935892492288;
        data[194]<=640'd43959229496528458163976736568683345462796131810121076401457149187859916309538850768156638556472848077181441029178100213803428187047330746916781469454970013301062867219382272;
        data[195]<=640'd28984109739734777180417480007390439540074389456297513402492803014577231713526894494987650559294555932782914831472740751026036625039547870733627717697004542385685306865090560;
        data[196]<=640'd45408429685593612359567564728385411155774602514027053915650564293145340492214460701166134108468391470978576710881794643877132728845830595892140500516396889641809103609135104;
        data[197]<=640'd91782817308127644169541681846885785849303172578708199914872552880247683226192793794117155597277285929770142034840653938089911443413430195407719628192149584279417094414532608;
        data[198]<=640'd114003915436497240631112908816531004071733617591470078440873514568067676416637855274877581594413704728664083336617201312108470926430928476357032411518464521092305266380111872;
        data[199]<=640'd245398191449428410631366527908118145371421015033361174462125805120803256466685809388919250862026673831238923030905172523667883049975157112397069389940664854907343629228965888;
        data[200]<=640'd243465834235675449704141772105912711715784591359178863364245292853678744150330764206201796300058301349312867892150315732322045322216403084700975037990067921568058136793710592;
        data[201]<=640'd245396243657297527513775463772225479566498583813984082702982926551656229634401830869331771829662447489038396566503749960018761411980589742452611931313416710928774564537171968;
        data[202]<=640'd247330396635885547660793708972650965406251516481582259437098175711026110748381206182023331231019549107432614576981811555567732731183226827048754519906570647933434157181435904;
        data[203]<=640'd475338105771844695021001399508166746951712566226662315140642134208987968178862713734560014135485679574280037065825762095031814767661850234893329278450206236461689061460934656;
        data[204]<=640'd432827258050787260695101400310594009075198930868246578456379435753757686716863800336919312244542316950788039733951656460357965712874694467438890024083763793034257829554290688;
        data[205]<=640'd475337982537591060259342519368045300393401399118896885015580863761088150753271594963400771407921351719046990382815924988770824121170030020837170971598674713831559630931623936;
        data[206]<=640'd923624480324554627641147324259754822990905754121402592531473652196979824240829005484202651824837504325292961788194573239526844736605974592851340706026323731804229963154980864;
        data[207]<=640'd950676245346703638042081619063858359797061953532652650423278163643629977624253351173765329545405464433701389493288553724440956842284766577634758534665237454635808496071737344;
        data[208]<=640'd981592545242913006796286229907701221992173353718515729090576393285866110190662173262596191092479881747058307658371887082777551435868708008482696100819419303153758226331205632;
        data[209]<=640'd966134388096545111593663040393617335814319051707339975146348867681306584904452414304686054109862390149152728147459776914943725493794896190567409332617538776190542730460397568;
        data[210]<=640'd1654022067136031027838475551964561481971852941082864693977713595490422251086691806264321704799898205150303818348802479733184302664058482154501905534102707981049084472778031104;
        data[211]<=640'd1468524263986896020567956634818988990631932974514848260098844124630762856229237495246879390186734233902215385069253969247371133372408820180792517620805694562307632567106404352;
        data[212]<=640'd3941828276688031868962948585298059899614110009971923683200270096036074299560402643959205103452110998910351419697504972851788650435563012977990497596893684392447596889452314624;
        data[213]<=640'd3941828277148718911595215143755415166685274649790375468151899561906429661350938131537295718039504975054402881355256351576396063539224565241466677587589410173705310384024453120;
        data[214]<=640'd3679039723222515367617770714950693859453497729607487866758367498627116454775505729122529076177424340862623094929044649119271323785623646848346122346773083151127142997222752256;
        data[215]<=640'd3926370124292516377027223870811214739943391363328226086574400460698976872736624284732244237520835337697659143700045646834187391274275242048312386078632653755537751173297602560;
        data[216]<=640'd7821823947832230485107772844466623648658076415990473764618482211629579674832647595089617560937891463846163930489615088441258326493135742646235708533431529592322962178025979904;
        data[217]<=640'd7852740247534084920895958298494964654665023735492684947948599372382928783407663691217699056847669866114600022754787380540710878361511004805755923142495862115800477873161109504;
        data[218]<=640'd6863418641720847591361786959088801716467857481216726821215433858971295039643816238953671902433494135642460218518299299344199296817261690348779144748386261178783571518517411840;
        data[219]<=640'd15705480494459916367902446344685852485222684299285647318159416183798587050560457214224021708462601823676899052096775359397354311416370729094407709723539148227654423752071970816;
        data[220]<=640'd7852740247688847380750965743195226151595691549775510732354320583556651197947712483424712060669188438819728309056601574735956970620839137183467658674986099925264700241755504640;
        data[221]<=640'd14716158888042025062916046561317603685393196866660281933040495604438295351818067986427938510762060495042486247808952842184108230136898552930291497206101409975761101316222353408;
        data[222]<=640'd93854655509598179697018174987440922892355575173592382206496282259021134884201525033806700579885609619425952101197652660130553820650272065643946971251081216;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd0;
        data[232]<=640'd0;
        data[233]<=640'd0;
        data[234]<=640'd0;
        data[235]<=640'd0;
        data[236]<=640'd0;
        data[237]<=640'd0;
        data[238]<=640'd0;
        data[239]<=640'd0;
        data[240]<=640'd0;
        data[241]<=640'd0;
        data[242]<=640'd0;
        data[243]<=640'd0;
        data[244]<=640'd0;
        data[245]<=640'd0;
        data[246]<=640'd0;
        data[247]<=640'd0;
        data[248]<=640'd0;
        data[249]<=640'd0;
        data[250]<=640'd0;
        data[251]<=640'd3705346855594118253554271520278013051314167415574284326239617177261309658398720;
        data[252]<=640'd164623458708069902826763918936602400973957899765456654442779638821494976910087624533689314208145162854249457221829694160387289016147615338725376;
        data[253]<=640'd192060701826081553298033274691018164526740861612476000147422249484490386182957668616305158675980335865396083913076447197304859801507254551707648;
        data[254]<=640'd94506059628706796067293808795622139611225776053683426000002277139147550810939422802808558026185885401857996706584489842552429981969057730002944;
        data[255]<=640'd143283380727394174682713898137671243355728278842792338214452976100056139799093304612049411417469644825613666698426104229106313278075185347428352;
        data[256]<=640'd196403436665829214026906207144036736742836253773428709490825908515258677382937727425042762854556254459545538771050837237065739446554171051264656428498944;
        data[257]<=640'd15543139489988962886039220272454040723786316440354806750644898456047873993786582466577304127667876675148152912640609313604228727069695912120619870673624472221756815827250708480;
        data[258]<=640'd15334467436756201055356679699057297338400910639793062948269762357086887995518720997673490945720005262418314655070682661943706890124640402089377630997493914805006979732936327168;
        data[259]<=640'd5935868013586485969676431769578398743956532775065080083104261624653786540737451075944104911451019682027212874344047831557271408939133412948760589204606584787907585685384593408;
        data[260]<=640'd15809821694606651611518164894341938485915791831027129498710067868017649602947283677004373007861458869227385893646044620121729025003737171447599056979118994376757791455348523008;
        data[261]<=640'd7904880751430341934676228642282300039405029034900361528428602183135401572980689812464679287311486621277184271774049577619898329176909503328846782318042584515661795989884239872;
        data[262]<=640'd3597057936158031624687504841778568097443127304978134725066768482266162956930763193235607067385097350721974330469001738886036586862028346731445827688647878437766160187392;
        data[263]<=640'd3420153447494521856215723258303488029184593377099887487855540181255803221919505547647464107026424072858292617386618820975885157073428275179404685223651733693155879419904;
        data[264]<=640'd2712535492840482848585086855529010909031311784634550809655487494585330683882973093590633729146793933965561349716098452922098950511493967049160152994878461080719285288960;
        data[265]<=640'd6958243220764716868216943784677056088386383170300241258974841015714800261535410212887731300845629823139557344164431082584677778946992277784968074828901556371042869444608;
        data[266]<=640'd7312052198091736369992786197160439202507029841241849359951771203628243815242975838742553510798227098788619273046600721276568816281181896864495690918363986493981987962880;
        data[267]<=640'd6132688940335004697417300390601581915256314500549668642602004479421935553196013827009557544792662341337201307264880241380984188138375589572714276654026284229633964507136;
        data[268]<=640'd8963160758951160711598466326342806842283185233888879630728006320208288506989175586914771035176237797402932432432065532284947349586668695641173814928656937029291596578816;
        data[269]<=640'd14624104396183472739959999030482133900459954401158064282378254403910310111285601204647329313066233958617724090717793439936318691122917291434274380407638944902658184445952;
        data[270]<=640'd29248208792366945479872048014615243666100802353438663178986756922828243762405801837633228465531533314572583469911635485140158143380389071728315004359607445880169769730048;
        data[271]<=640'd29248208792366945479872048782691331611202986070084726810199629833903529924035548425072953627269936716961542475079320812528409464538020576258903073401403069443848806596608;
        data[272]<=640'd57552926978528505621683907095543817712652000378320229118097601465280456945736465368500337885155043745016943767747374109770338407526448824488767371366809894418393769967616;
        data[273]<=640'd20756793336518479532298935316979051788112338150429941420753824096026635401633449590027841758916222226784411874891051276218976409208874209982844983103671945750295735173120;
        data[274]<=640'd58496417584733897244654256702132301814733691883396197237370679471881439820502318248456684912034503620395875816504830821947598636398860114336897662934240996598548860502016;
        data[275]<=640'd98123023045360077619870524609922614701149675648317561737653857224162827667113698765556414216327625032204010032691485124606872713519082649852831091482367540387019380228096;
        data[276]<=640'd237759632763757117747944647640704587626916665356715351656885452729244882792367310614610872699583963181040920695942200839073863134615396252995819962961658453127515382743040;
        data[277]<=640'd105670947895003160785901703241758055523143694558778271357118931532074483150715605355298852911016295245648429987716370800911169687449762982240873859054898268413789944676352;
        data[278]<=640'd445327566128941881237206166061486237344746508191208537394006274564524339818139666286222302174591405281017038517562092067659156727138081064516559439331105263655478718627840;
        data[279]<=640'd951009046959525397267737210539688935906763583335898658327935727610790619640264338171416345253209243718811626142695715628832376933103986846050196113013853947458948232642560;
        data[280]<=640'd966134380747285033468066333718559864939913188542701536870826196240865767539677334687209799877073836893787148807727799866139084081705726242944505249680598308222076176039936;
        data[281]<=640'd1902077045850701205951566793581498974711071234846556832357727607583536750383582482982884102713210142417510656511147292551230198601693157847037954983010597620946584381423616;
        data[282]<=640'd3860763556958158003688684804927972752010406622719783254147994157397082966473100591685665459220633996587651861605481960746203055097027953018623464981442496725881586913902592;
        data[283]<=640'd7706431264280295817204166831552134258069581463722124716736489623813985502134484946064897446044192267253278440700009718074178068238321790371307763072641532795822737511677952;
        data[284]<=640'd5736422886157545576449561761678234181588449265214775904466424693359812090655869142874517657775466515508355158881319625893296304740354948457894501244229565372664805081481216;
        data[285]<=640'd30886108484957410563668069152698294164879844886259003419536774310787138105739591439229723794261152213150918103783685625483341103631512558272904831877342179272146251478466560;
        data[286]<=640'd44411989815679494484593196890967122245618901888626146373206603561851389242393732265477967606142173305617672336533886498852293987825361276421362307414803395196913042046582784;
        data[287]<=640'd123514242240002267202811944607615273542644071778736040147455287070970134454629954332783732838494729156109768818157580552904893049868409417657092343848404307513380815771795456;
        data[288]<=640'd244401806631885879797813420945831026315468537940322192747941680002124803380662253385755048061353051502792002091406730708325296751316359074417570652008994149298308073482354688;
        data[289]<=640'd321692557092231046691720458514730603371551904493412026246890099167897018637708499768333316713077046477063200047040131386493496926974235873966321262589616548279819897640321024;
        data[290]<=640'd851134197745595439914990214603369307995166526089591500489105080925895690993635211455923765214491479853195945271122521217208911346980220007657020034288215011802387606579183616;
        data[291]<=640'd1956391929328531326497896862706604546025229891634347742097154550205665775849881125232699134932136528903781635127794734913527125546180571507655256231564948105804455560270053376;
        data[292]<=640'd7389931686690796559139570623181150085426843169973208395487222121929592857716135244811133292475626542479179660319456007150315059347370706008013769005760962831502662572523388928;
        data[293]<=640'd14809843730883932580954645435173173452079010429014037370207083980314183749564254088369454841547492473804434558826789962261475185905708888081925034519152859928279180221899341824;
        data[294]<=640'd55341113272288938100119492794114502189109331988785336741306812721409487906389560954191813205951496077439947900095689013486686997681722278246746649317887533938537629986425143296;
        data[295]<=640'd63070188318323454789510244142061136940183373161906455985133862809251306503586932528632083070096584385402826073386060973907864653418866678612671831592884839446761163594152280064;
        data[296]<=640'd29185802549710539333898127007043270756357001211448329405185814202034311210132491302464230546414734172130796933175653336869438473983147563305230363712263917675856648530691096576;
        data[297]<=640'd10883232073903209524097672007823408766361209557116791465048070494246777089234708769312024928432970622954228324011417942500599992101198657011290704780106621156872814171831402496;
        data[298]<=640'd5936865578036307421534269808306551067629773177144961009696962701441966691846106451015053561451444276553348679663358847998243171938417131795105566304251431892479747018389979136;
        data[299]<=640'd301916994428585134967254959400106686836127964354457047255756799850900859641364869438044355074315946557277479482109971754884793418126809315981308272409240370759903425331200;
        data[300]<=640'd875559283001459420671538492648635819084427819612145138129483761989064372763221517108478088574671074700946563161213297381219960502046021055573406173329047087117347843997696;
        data[301]<=640'd452875491421446789272858629304287973221965778460874879992075950664060083910248044568852584510337634154113570712164816550223823059272230506310484075578751984997100924436480;
        data[302]<=640'd815175884204314759127328556373915489190148491982784350942791460040156780973693834860284142948669919703315621257466286054434668432744867869294140954123950474876041971105792;
        data[303]<=640'd905750981950140372336303233185430272116362837396349719828432806253878474493560355172245056758200390539107896013347908294253021788961150858375101722340580307437116553428992;
        data[304]<=640'd966134380747285033762671123184798965629396803793072558565141631376106418515872252176393036711536721023369399257591031598245314229568148410160464436616147718581359657091072;
        data[305]<=640'd935942665082327514863739788269748081109806627806827196503059998147092750431445514893631502878362524812508253993840162772404032386554416688396782322797955759082608248487936;
        data[306]<=640'd962360414610859612043228204026510758805787562538244356491925841926871077517706771881358756988148543002830503997847300848503315610731022924963578783854944913632556048449536;
        data[307]<=640'd943490599000093716867884794839060564593033576668329409800922932548482239208056367960833201166794542928301895742996403145126374852208806979830760348056790609320068046127104;
        data[308]<=640'd905750982400031754278400420252256458523715964520965990077174196527850845608807796106621005011361830806444339823937701730703138605646518960911344222390677082986817175683072;
        data[309]<=640'd935942681559599292851308649202732842235933694300473677494394635923578301221402122995956028053541940962616073141229007263035031584798126213223899137904760054478186748051456;
        data[310]<=640'd935942681798604087557928244402924203344189430559580271812309238987925727625058154989342914624747996082503629001907865870767296260964138565660463555574486679755834248921088;
        data[311]<=640'd815175884204314765333689835731114889931913009833965115189232046046134998078346634832225181242045332623851601060042036886653361699658282966225000890105055531895204196909056;
        data[312]<=640'd875559282987400321257049821837219397592491360891848331856658835491406608914280247541482911460415793116295936888695287357088737564778060747194304634019493048531414144778240;
        data[313]<=640'd905750982364883988635030758255729715149636366668079651206071836952746257269279358673675615898014740444565011769453764588249725424152224651041434748205030046543397190107136;
        data[314]<=640'd875559282558597594139133757385966052017877111266055960945722787554933034603654081467795531711576533825793557892134599995665407144039450367592436258314572945925253153947648;
        data[315]<=640'd209522572269477268289203618641472811360241783462740857970598485771965814021899524208253650791021279314388387741873250872481220818430250952347753895690240;
        data[316]<=640'd332306998946228968225951765070086144;
        data[317]<=640'd0;
        data[318]<=640'd0;
        data[319]<=640'd0;
        data[320]<=640'd0;
        data[321]<=640'd0;
        data[322]<=640'd0;
        data[323]<=640'd0;
        data[324]<=640'd0;
        data[325]<=640'd0;
        data[326]<=640'd0;
        data[327]<=640'd0;
        data[328]<=640'd0;
        data[329]<=640'd0;
        data[330]<=640'd0;
        data[331]<=640'd0;
        data[332]<=640'd0;
        data[333]<=640'd0;
        data[334]<=640'd0;
        data[335]<=640'd0;
        data[336]<=640'd12486994201263968925526388919172665222994392570659884603436627838501486955279062480481224412253967884639307724485626491581791902717153141225160704;
        data[337]<=640'd24583769833738438822130078184621184657770210373486647813015861057049802443205654258447410561624999272883637082581077155301652808474395246787035136;
        data[338]<=640'd73710203609795729535980154794843995995132182625350912709051664406859090245628165197835687502347750630673527905100418845335086049594509144682366339127532042225920770048;
        data[339]<=640'd914006524761467046246024132760086162962619374649522666703079140677271422870192279002566100199070676064695244297010329003454097210310540913714464355592530913139808534528;
        data[340]<=640'd906635504400487473292440613900432293252030634679123427448206294289210514305411264692913791768848045288226325177966388209761662051662485031251298458216838403892107542528;
        data[341]<=640'd700246934293059797211539556217256941605769491274685356528253766731566331990665604672151628558151963794144959888746829434551697116598293395637289397281380933363593904128;
        data[342]<=640'd468059792922204322845463195675771758673244899744315740138820751504407273701288452892034988941864058094584743081503395996587333659063419074226067306546309264954567426048;
        data[343]<=640'd350123467146530422348554193568727120562088948061059760410582316077260771100403352014607004222133271320986773732743865132659861144199593188580291273165213030884971642880;
        data[344]<=640'd200860304836693651044160633614355453821548499759881780875650398766710729725308937582298415985339602891446742722882529188463019915584719165236820938567154145722198130688;
        data[345]<=640'd57125407797592305789182949068661305430805344439209744049078438151108419045905241628086835498606421911039482145234236295696362427748299601630334658598715874392271749120;
        data[346]<=640'd232187141370856849191583292938373363928899308817598367467960663055349044903157134042334901271758996848109119851868205047589080602959485137471134567175712856548954865664;
        data[347]<=640'd103194285053714401069958974629347846307315328371942953292563506771234944593908165881225203106270921879235788320894177559987274628533968420321100955078821733736174845952;
        data[348]<=640'd399365441891571393644527267105591720604747075309397362525110850105198274777740392563040167561403871829432700929312119461866805484812825432718036663533568;
        data[349]<=640'd196427011930252683206627629994905142977083611746243442837034590664318407638846979753891751787749349487693021566835657562367094120747895111052266840260608;
        data[350]<=640'd41049116595478066567115869541267401395421280016614577384780797799853230699299159425533040433044965139284870137927809310130313987724697039250033865077815273149131438555916140544;
        data[351]<=640'd63281801703534896714194131352350132913073291751457238518593586904355540097919071624418017772599811157851312416478799034879039224974381310200655802881674553650069104564753137664;
        data[352]<=640'd31163147371000386653876555548836746070757282811897280245353393547627612047638380167072267160376436720396908006842184591930946420677971472300647020108765113618059187637142421504;
        data[353]<=640'd31588419953383419766670077407225298662131860247833161116448794359865822518953646314063880527288106641257681913620453535746913792217978547926730083808882525129971986864996876288;
        data[354]<=640'd54396626340002956752453103485447140033557716898792472927265237561870967564623596792896362902035215687220700992698249113668949634472902536854495623745830431481182804639081299968;
        data[355]<=640'd55402023610589205635099157229291333918844106404197230491095604789876855464941294716104191117986498521603637105170519064965140370042525366785313628680557944724100432171431362560;
        data[356]<=640'd14152359093080780070912023416844838623004737610235925387814604171925522952327163751812881291118383636675005525871682431674472680615699397521886574802230821632792770641920;
        data[357]<=640'd10850141971361931387700663158479359060602132019627895837600315229636946625625699473468268046124152248436320637160756844393945841530374056207450697306098356793382522585088;
        data[358]<=640'd7076179546540390035459108479937192255164175604855442561723594885246911413979290881967801619108636603275330171241152003549946276500493051948840013132433448585272190042112;
        data[359]<=640'd14624104396183472739942217739466883668664074806039600686275409300764165258615630053306875035675678406256527300869218561050436719803815423569445362920168961829127736786944;
        data[360]<=640'd14624104396183472739942217739468372234367273248866278380288814592290611355771015453541482732088756633040293090058271622529676552720902057917401815236643744018340524326912;
        data[361]<=640'd22172029245826555444425127060759996552589634651789331615946836882801172242336503443945108028955892026517705730465284909207792069895275866692079877057715779010137683918848;
        data[362]<=640'd10850141971361937963942394415730094355483532642569506341387987779548158796841695919641683601197521946624041948930365358897312616579456027701611424020697422447727205154816;
        data[363]<=640'd29719954095469644378170563097872206209636821663486252301016242082621457072741146207194820907043052769717173373410470403986065493411977066332029157134819923714132108378112;
        data[364]<=640'd29248208792366955322963799635719010146929056849849289767877404671352400105537570381145056957055990385415548182294119927021499718708015899892077753990196008213023557681152;
        data[365]<=640'd29926342623399762719926962959264344205607505960692048416663204564111927924710982767636134826164983933137750100139570935540190328724761449741802589621644121018169850593280;
        data[366]<=640'd29572533674190952810447759335134422747194641997826938546723565158691513358690842383482224676500626311141189163176048819879518914133636563578929320789573371741417628499968;
        data[367]<=640'd21626573725054961539386984052205187214348054517630109966605246800052995743888502357199944206239121948168494099495706537937510129934102463524222942047660225052815789129728;
        data[368]<=640'd30191698934621845857146711765317732067513819720552513437630265373781508736555188649409094966426245198899589164482967606016601335681013866808165549792125971369890020327424;
        data[369]<=640'd29719945983365702464682367537860167856402110576067729699083700944898974980121347323792220745008268118372542771548312678408805464845163665122005356051955245247658922606592;
        data[370]<=640'd28304718565757411657874357749156455513032593500155055328509865227147302300687552785493833425771738929944187939655948540794386140065623631872955891005869699464246025256960;
        data[371]<=640'd25474247028323367802643764711593507074480487991739795089598877602597445783187212953881584395407941919544664771096185384190982864998880550874475849596602794081102298349568;
        data[372]<=640'd50005002550658591257100368565477051547809869846266997710678743511276990087840785421841568406792518220935985405687893439681173210772028436247459317306096404502481125507072;
        data[373]<=640'd20756794222242130839495447454818256376935415453726070706028280432657290911509079456815503669407226231793283790772000173497223507585741148774989642607616615036545727987712;
        data[374]<=640'd39626606332290731992755731772476891916247156466691704338378844848882506486259346724149359122633252639494063629359892234345733990081978680693763247903558311629460231684096;
        data[375]<=640'd88688117854970769571895942104212672458659812447729999083085007254771470327891593219409766605282963115305040910511941121543554192777420234426974342763779321886087067992064;
        data[376]<=640'd86801136642559998895775166424895914119923064852417202162931301544462458060395505181386857761213806308877349029874655614004543277310071570966178266891068481366970588987392;
        data[377]<=640'd118879816803651720935508745203976385724465938981741327387685419386119275791181087136823365291869747299076799681496945300659107677246992036865980624952265599041323927601152;
        data[378]<=640'd177376234585213090406517682859696877491865861775292827838295056597904523000356777472217597091704562238794291092143036260792962067902311577258082718822339837486694517440512;
        data[379]<=640'd203793971812027780815263365947216626167743138942968956853483052468478237191917846816290681873438086469890719393665275565854846946658583488854510613362750746124830730354688;
        data[380]<=640'd109444912091272005917863791252048944274983073672931972623408889997440039475528779130545250857357323576014340618608701006275021480066094176368742624588673994854599437058048;
        data[381]<=640'd415135868473698644233534758722865578184495121258408402377873845774707164541773981672326209864773023609703004676172476178472721568382675496940829478417839360089258673045504;
        data[382]<=640'd460423417599675351676328391867727825571660923958374328559903333674202714352128848619344279873110989069664153024100073592734092772114363594907292008485786992442074015465472;
        data[383]<=640'd951038532826475727467730632557510394343342085153981974196769944048774682863452322921689930187362102068374014072975875143459661860223801111861271523881893404618823842136064;
        data[384]<=640'd1902077063881504148232602986342275838783753835424930948017767706782791473363754244219729491425821803511869746208824397962869395795941573458434075871166008202573374468128768;
        data[385]<=640'd1886981214182217982823638360110083511596770897338905996183105817351388338757208501062262966840356455196321500358142266979404789540612380639365432888224489693356367137472512;
        data[386]<=640'd3834345824912123729841328688811742301757377495543392572999311606213709228428122520991093643198406332340794059052113029209750047777544848892846176410822675476643281184489472;
        data[387]<=640'd7668691648980701123241828089231509703625921067859072977355561010977687103105542672416551910371556616318247216874754651792697262060372285282107755472460978190289868972621824;
        data[388]<=640'd7668691650724030218594569894912585083232661710248398967244830146489555107584793280323248720430310281876772217489259791487198895099450231908461997766895506902768493021626368;
        data[389]<=640'd15337383297792692979086766252066416153913901374861734197620209447583678935289533019688532560274548009267471136083933326407248526607531791695545730480189606363774112283754496;
        data[390]<=640'd11352078975156634103522867597124629349672312482333323000288670855536907526180599801054578507965230737953580587076357732018793455713089569992542685512558447168809141998190592;
        data[391]<=640'd61349533181216925145826927403922152788750142596053093026902406941033056397998201122800004557445714220405422188049047084250177053569982104643386739060055673734207531621810176;
        data[392]<=640'd242982796766852144072382264246337268396123000035492248016376329492360013556958658350421354670940663230552453547196263371261501253128791063130769381017409036816494038655959040;
        data[393]<=640'd422200724400151685156063816464896652024050580658998389294879485516429634790026887685381920548889268223276095349311154974990691315974182856362607379318044419912297265603018752;
        data[394]<=640'd399979637316784163568254169987457467207391649784612566359964041239148178256502500607489478232744469609290079855812819052998826949389723037608883654551589959659040834808971264;
        data[395]<=640'd3686768797872081379679583549345711108734042488578653648062649742641941522671147230275672794379605616426112580968254925132075399204148848884373890951514622701000218494120230912;
        data[396]<=640'd2898403143529612937380598190062666877450871181688698397183040658071051676032206233868690960495638718906301920316957453924837185160660273639128459666471003587822805946141245440;
        data[397]<=640'd942947156306569357884604356991914998457455870655810946954233899076145591219726172436225346246586251938946937732646354010217269541705316456433389861444613974504523358435016704;
        data[398]<=640'd463744503668152239587374942775385286911239319470527305795976392986616314360551353884500371890389155862350726119278085220527983074461155598935564728527315772228066083839410176;
        data[399]<=640'd185497801561918042071803632046051116565557144322562822081622334762447885000685572288931699776412054937452378593423790705918891687219517177831964030084138634924947863574151168;
        data[400]<=640'd403102675991070395912308099894871150966600018704155306478322071258333704875452073665852315093489527436270657083873535864707968448300283104640742697878673465303629824;
        data[401]<=640'd38491662245232981164558545157669895751727176974360612988132016033434028615688539057448151047332054549841431657218767323136;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd0;
        data[406]<=640'd0;
        data[407]<=640'd0;
        data[408]<=640'd0;
        data[409]<=640'd0;
        data[410]<=640'd0;
        data[411]<=640'd0;
        data[412]<=640'd0;
        data[413]<=640'd0;
        data[414]<=640'd0;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
end

//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)   pixel_data <= 12'd0;
    else begin
        if(data[pixel_y][pixel_x] == 1'b1)  pixel_data <= WHITE;
        else pixel_data <= BLACK;
    end
    
end  
endmodule


// The whole VGA 
module VGA_out(
    input sys_clk,
    input sys_rst_n,
    input [1:0] choise,
    //VGA
    output vga_hs,
    output vga_vs,
    output [11:0] vga_rgb);

//Wire define
wire vga_clk_w;
wire [11:0] pixel_data;
wire [9:0] pixel_x;
wire [9:0] pixel_y;

//****************************Main Code**************************
// 这样的话每个VGA输出都有个时钟分频
//优化的时候可以将时钟分频拿出来
clockDiv clkdiv1(
     .sys_clk(sys_clk),         
     .sys_rst_n(sys_rst_n),
     .clk_25M(vga_clk_w));

vga_driver VGAdriver1(
    .vga_clk(vga_clk_w),   
    .sys_rst_n(sys_rst_n),
  
    .vga_hs(vga_hs),      // 行同步
    .vga_vs(vga_vs),      // 场同步
    .vga_rgb(vga_rgb),      //4+4+4
    
    .pixel_data(pixel_data),    //像素点RGB data
    .pixel_x(pixel_x),       //像素点横坐标
    .pixel_y(pixel_y)        //像素点纵坐标
);
 
vga_display vgadisplay1(
    .vga_clk(vga_clk_w),
    .sys_rst_n(sys_rst_n),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .choise(choise),
    .pixel_data(pixel_data));

endmodule