<<<<<<< HEAD
`timescale 1ns / 1ps


// VGA Driver
module vga_driver_color(
    input vga_clk,      // VGA驱动时钟
    input sys_rst_n,    // 复位信号
    //VGA
    output vga_hs,      // 行同步
    output vga_vs,      // 场同步
    output [11:0] vga_rgb, //4+4+4
    
    input [11:0] pixel_data,    //像素点RGB data
    output [9:0] pixel_x,       //像素点横坐标
    output [9:0] pixel_y        //像素点纵坐标
);

// some parameters for sure in the reference Table 
parameter H_SYNC = 10'd96;
parameter H_BACK = 10'd48;
parameter H_DISP = 10'd640;
parameter H_FRONT = 10'd16;
parameter H_TOTAL = 10'd800;

parameter V_SYNC = 10'd2;
parameter V_BACK = 10'd33;
parameter V_DISP = 10'd480;
parameter V_FRONT = 10'd10;
parameter V_TOTAL = 10'd525;

// counters for H and V
reg [9:0] cnt_h;
reg [9:0] cnt_v;

wire vga_en; // 使能控制rgb数据输出
wire data_req;

//*******************************Main Code************************************
//VGA 行场同步信号
assign vga_hs = (cnt_h <= H_SYNC - 1'b1) ? 1'b0 : 1'b1;
assign vga_vs = (cnt_v <= V_SYNC - 1'b1) ? 1'b0 : 1'b1;

// 使能使RGB输出 // 范围内输出
assign vga_en = (((cnt_h >= H_SYNC + H_BACK) && (cnt_h < H_SYNC + H_BACK +H_DISP))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;

//在范围内RGB赋值
assign vga_rgb = vga_en ? pixel_data : 12'b0;

// 请求像素点颜色数据输入
assign data_req = (((cnt_h >= H_SYNC + H_BACK -1'b1) && (cnt_h < H_SYNC + H_BACK +H_DISP -1'b1))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;
// 像素点坐标
assign pixel_x = data_req ? (cnt_h - (H_SYNC + H_BACK -1'b1)) : 10'd0;
assign pixel_y = data_req ? (cnt_v - (V_SYNC + V_BACK -1'b1)) : 10'd0;

// H counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_h <= 10'd0;
    else begin
        if(cnt_h < H_TOTAL - 1'b1)  cnt_h <= cnt_h + 1'b1;
        else cnt_h <= 10'd0;
    end
end
// V counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_v <= 10'd0;
    else if(cnt_h == H_TOTAL - 1'b1) begin
        if(cnt_v < V_TOTAL - 1'b1)  cnt_v <= cnt_v + 1'b1;
        else cnt_v <= 10'd0;
    end
end
endmodule 


module vga_display_color(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input [1:0] choise,
    output reg [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;

// some frequently-used colors define
localparam WHITE = 12'b1111_1111_1111;
localparam BLACK = 12'b0000_0000_0000;
localparam RED = 12'b1111_0000_0000;
localparam GREEN = 12'b0000_1111_0000;
localparam BLUE = 12'b0000_00000_1111;

reg [0:2559] R [479:0];
reg [0:2559] G [479:0];
reg [0:2559] B [479:0];

always @(posedge vga_clk) begin
R[0]<=2560'd57773361369990237240164763066017403883580237145113726174237184464633430536881379704668765882949592769943095726393019195080462436110363548445401715084698459841028804720554902658797917499672002546284335684299428851956696145193687051064533984917986117588265178082279972299963448370517262940711401196393493785948946391031390212656556196078529908776626520098456552924873713331570781743344007272375654812391946626983038622980391777307398228455721912090214557028816033489281662535282256277936157945663097328812396618759730569418434161833682606279052447384793699421351145666432457118783159884422467460781508768303013775325807625349073694943406561017475943324878474682604333835662100419831213315705742077550981914250740031789378960689210356679965010245019266395543649263974228514;
R[1]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216088429764176574501715678693841121967005747024074171202276246624088493021737110524699468503125261701810236879024817040830069340769061379279873840948439722211629580351034406346611401581758567459769282064012343433941323293442646943430773547195416564914482697354782658914282337598440339692087669623842130433660382000798614631721697639771750262520310434245839077123876327820676950438156811783014032158960479487655080012756721387039865005655949661088204289626259320903591019200966799666230500896552365794627077346660489231099739086310161685650431601195469583812466059903344102030012484897204042957444661445739434209243740219843250908962234992368789134055372950217250;
R[2]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713664168093303524910524452971021490350172490437450354317788664934684426241290213337230996453027222904174072909745368027041822195712787735534177734524762104051879940128748202768596837656022460235736229405418116829153124227614529894034675531120700559133009090840853794077967124796479662784386085477138356734953639084599901164502212000999199846592724083100949017437838690984147965532103752764267723902025581347968441414756199250378304553269598740910085392756620186487139974671238414387642749608856059769244395355471496258406201497544120169880374351761307784896490999979584268371927157158174870201941787391115795171051840526176990938310207469184241502619672376242281259554;
R[3]<=2560'd30692098227807313533837530378821745813072426625859374633279472014017725084571737912433901425251006783517886740174884802759395351739350849896827899861749878862779748577022881944868651600722661676566575011048452230221223228844741781002165358656764311248043797008065665858311197977789489852738981996677925463363453940761485231938941581650736137272199444992429990747765471568206604260816335895789745552689506320230048975817128513437214414776577473685708320464001876218499491098968630421386375051054742019730145178180257970951194389867072233349762934500677328186609196933530102595878836502922044829061080386537378917832637661044580598062213217988030162663890992245289257188925808648386371026818194078477172116958315263694159359436283603367320975536096054597340533817602089506;
R[4]<=2560'd30692098227807313533837530378821745813152011305451294277942221797086083963356503086880359007406440266948310936451834750739615634148023284954389064762283809336935828302565986918637568481961293298878944554309717815161532424378801406979614257263258798831516965528472238966316825136661402276463515125837102873914220503442617255076920930442584298492242984955486846082067547086784124487679610934875542805536768030560710315650163080083461474184200593123880912778369792713999373398053029104786826781095602620284752208541092792176921609261161114292920884755459921480922980927002138087533411607297392310147211593559239205847617391138605626605928180818276444493830926783147991457738316715814963357266900926984976635612346160073896314496476167480011607541185787931013158618452337186;
R[5]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478987703174675699725083475815399968900807590842845489558260995171488520159947707181790279877926310771254769280586542744827918100057703622466556989012755670758340944933631687589444024697178887451180323965527020605167072868767723894035475864108315467691297843489672465763936698519735085163285856945144331545828622621777740111855337044153921297390757054460163872846432058011989492667139067022033017353005124665027437016174598347659906551917911560368158440784344930682542765505644831421369201536609652847972933745355670831166946410418786978254126395062603036834161847977811626873970108985727738539551587450510526002491181247768256560180969668604819134280760369087320496029771419378792931874;
R[6]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661228337411958397705942183078003852262345519021338547303876438626762374586278906266824968170714550572011111305369817014004157502333022222607221998803717511837111783557950693373286481509525038020478427842498146332318119171025486380203349924186038585457182968459033775049674037702434105617821638910627835641685827602148171788449442362428890673440353893563812044794362130233262138235007927854794113972556379034947381089143541543805462535957630439727825340610556401528040532275390090830587842418637833881285476050649429224126877366278382281162988194683867341786438576625680766379289859282365444275588431927226466832105114736677033880745576727320351568919027414277956130;
R[7]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661227616718640421333015426271627208581362591230083995801291952254796521672200830716457480355152468402572808827371221927929572757393964327899000909086975306328409277648164047024307714445545726697245131823913066439449876077387349488603925008172744089187704093106423790873414702623815711455863643304688464036543229931113422718259615122764882864979858234361285355909374605204681309062399152433320483141046017484670371885637837570269843827337473987875512296330493698309207467782443639509492324690524985884373850041758092182843604416140145733961997958277958773189341270714818600787555705801468788889920955964564172251657635190035917785655805118394890747196693227436646946;
R[8]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516479804513887292444896417371762181161000709713768085153373143030196806614527170808845080655822930521734703617094073296796865624609980420913154456523598113580409695633353262931999136865180691564256507186550180304715173916042630109830757232897751070177884065717851106558278445780183648676823415547724570008698754571357211806859109698424524692351651367547387800704839390803636878102474107209364163087812580379650339215798907736690761696259600484244999417137391231866947225687083452469729851008573714391118704579974940816577136067046700934830983617597654623159020452385950089813909939350777243145338270055953855353172229571096182291491554342109087294073640886854261114098134671229727805678114;
R[9]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516479804513887292444896417371762181163685458001673307052009043586791471421229999582145415440846807209742169854505089433349763973193160174993690785591753820243093829099554795717491278318997651658106869117839056449644986885454270737246423721194871969778106910540325695144915095665951793550566480752875693022406731307098456823636855505930734402512387565602136962719148921181747382410581673058060694213752620539997364907859384069633938709796926570609461141918080885098258138206452652718514573131239079954553768598280380553422279833153474939490268775554038894838486824230852434102975586602593692199796148893462965752114802632518037446214703997677023006105555046774465938746066927213394364867106;
R[10]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770577146841253006716859050671651194216427324151852519691032985088607556505151543216944595795796979507321307972496371515043736824526805521145902840578101662905565657470123075981047119535954824270350569510972958522006594592222195373586524650066147204783218845089299672610460152208032041871122995529937091173067542373540673959967865756150032833391312788244701752289126137237638430800910743368506691210016277400415940304687529495463097575203297658615017949538388928247493943257052513890208321150256066847624732058430599422385503308274431138014274193886272307171673208271690921344539156057306499691298763787755824024714903894453408818784455871254467523827946217188991864018641519215515812201898530;
R[11]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770577146841253006716859050671651242074967803215427862052218139313921459498489560711432190865931790826813053658749787612410757884306883841178783355085511103376449297413748602098600411371519896577503220114810835088571494690897939653762930109632858014598857622557149784458348534935596538082151858552199925907223007751013012981232062603836861534584740159494518015086093586279610426092064029854509524665974274754758656922506475143339887801310058934563030724831914680347189571212567168207120819070090014898934447950187115967003881234269910936618066013263902880470495055655726960496384256125746307520984938133514767885993152796504772239334252063845824004526655018718621351876771242234487150362108450;
R[12]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770577146844656387931809647169194031097842564863688708668282928215194353203274973249964507359616765307549012600366109823313748675153935594579397233076546247526379596538838003404866853941540927543791411120123524808649632201748086011755784882819343511078009050146836430117020445385192449178734307384452633554383340237951677272739100538625402455777060963823640647463073417310081771555590587377451329641713390103791308009783742779070333077069458785379145697910107378052184344616623554202065766936622649727707703150278031651793553886997997672440171139457678770859268868472922342328548896565508129339296319190084827224737920422202416459396626145062901560977657367719256641665552020970233124586922530;
R[13]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460436004455500951133535289977962086482813396623742845387405627396667627003888389847663839254612124751246866695494814846981868481839718103862091948852888606926691384013541689660301117565871615654878948164851830808092541324006725202275170220713405020212330671269703161745525937500469247311008172458273578169433120538402635389024425591338120000138715847955772368627691804238130967992038202739210609685841959804981690817054523159044664121652644044215815940327583419251959509941577781087052215558617912831229603838868339930848565842369950274061978184713725617839794651710865306928161851241961154578863894436302034546224437698091167810031881631285408211131541908407896000822989320668976031407429445100066;
R[14]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460439761126785901079117762509515395512153994510474385781356158826256150431744019643121246522469170410910627958098096812201302437120632600791487210392633164134602897344129868363444960065932787245547945334676577570590262895484015118414978887810483373385213284787914905134344366798113499369369693190735999125908436080316067719474820596628910659937389028824068100756319597500781586365356840820399189967539269821050050769394965562515812600162604518743692809269804807738144443041516172845690189395686383179417198160593659498625064028092001169722132214537890043497402675179831982526826730462897848617750745139825135338137370029748087669192794888966875647539543589213119514758348256687828882569215093121570;
R[15]<=2560'd57773774597272069865343387443957577157171419115330751726028671677111126571881120180076725499374404477624141084618576618988030561947118405339958765121562973059445710653955943953211226048191052124449808868339360095192249762676527520569677744213363790990162129253519361892866462809135601927043196658611136009619674116096322052327748488824140232475572928196407914842093951897404685369893814664667825221211016523699444492249710401582879724456311794026059032845368918437794556567726287496242011783715291691427174666100556735107936946864320723887784987310607180173296643042917919733827940469031872400732466204883710281366993742979328998463584949517348025201300038563553787909474198250214033598292147213024894888214018348547848691931031742993876569773166584526005545580833677858;
R[16]<=2560'd57773361470875804093833019566451488029810786959545174181716649553466660748833806846972465752516924522999249499874769953927742992076926484267667269471714596692472904002995130036422065131958356176079700514940058214216446728287604318129842854162236295841569953770603035943831572650067133483090163059169929234435271583524343118399160877208007233855965807616970759880682253600515360444611985278515424027616781969039011346954994249708163359862180560651569728049427401239565906715211967880191437940073362885434949951952773504927124322674959759113817614447998967517975541079655512684016067965977845366843036928104618889221032177165512605885870779147713545713597779217845684787190500292725937475449713921996811347103256897184569036317885085838824176500855424621159851289047343650;
R[17]<=2560'd57773361470875804093833019566109674433775464096976142774271424736635792587648861165766805244872608383672477961986805567690923346316645683479232565245606614909389537636457227536738052372524964957608537348177332123493937917282757528339935225431899093034495498560421107396587460745175077183417201728689551322645898607490413446198925652343968175150787639707364078961049466034735249016343639346282227403752287081025271628692030483033795325387793733932908505562006775552856639552758811248536801175876579055938824502275674635125668738374113882171615325879277508011817871972576953256611874614160316403033380995203926213531526204462163939872628959872772830129405947845172299906385375671964859558635406933816238879513613790243207710119154800825233971682898364502157228529720369698;
R[18]<=2560'd57773361369990237240164763066017403884853611448456386255867676658629671397973046024396669717504161779406207433729881804632830388313982112693717344690234112952941704705490473167642925897211836657356168768383279665773847924181611295628614152549340470985191458181115937155024939639275459054007112529367370630635550795826391349507536951238852005848112609170450200589531548069513773231551949686680256985184540808808675484340654693335310425185700011362497442488260733650780454295487466917809308488386891788862786710633625638210361143245910833584062733809301443081269173907082378449633299252001601164058226799463248232030278372762326658420503666360035434943332370449850043493079148391725980814098981652768716440863558012319479466877925739699053421983004807204435176967060464162;
R[19]<=2560'd59571728114694891677698238079748136556057732165180109097654362621880363465268737487360071908961733131164504939192006519823980234891618468029637517931610246730999394990191015120853075450684283843740434658679518057653530228806846836558952237115222639352060483755624671920051920477941884392700064774772255352155450249419754165628463633608862375751395375611644648179659999779039325722497569628997648221886473257622174964710047760446494064604419562100120119276738798257878639216781704934790801796897608292386967630475473192575720453409603653375592246468097255808774559887711900680111132881020770595623469842189686112151659816639268966762871319380123136302717123961260580995683697796195638483651311451102858930104152141504234595323277749127820328946656571294513889609137660450;
R[20]<=2560'd59571753941400006216771902103370816045601972028715787622899576152871784209580395884329639732451681690721204826241716275175276250307392354816321749849389963033638190747429773512875017746615015998028068028973099971845587919751251637660724245741474581988878169270579084774328333318471646743172606864845169022726530830940804808894476511773295499433129154661786035652938976446796270403752673192709301151171653331211659146286483348704835874677797659661436896973964627512297735572123933752333716997198612023827309549802726240861311139322249659007172962260623117036869938192887566273514916699477005804863368367411138578252362682697176909822849972138790004963833524897901326993848610302012006459197142577399356703267532261928150088212478912069378498583626128760472653992678269474;
R[21]<=2560'd57773387196695351780706505306281763924849086410639552313078743576200123017318038823444762673309893740702224549084415660829651178305720719879453644204068600437603116522976601359088293716169880283844329931389804165030773303512590463094051021114826609191183966786829887669850421303369613317080545649717477252735635427662987752532993244140406124893933609911112789673912076938952629598182435710733446588859774301267485833166052078658337297832532490630063200297076878284418742688818655008220831313186393135708429478948905494594174771769722516875272934865527103440169958934313280197494052930541998492868385971945112146561623600840632331772963449252070457666304477218990909911036801708391516619165531233857366789266779092989235653367305753228407773578530318045873449076946772514;
R[22]<=2560'd84855037739454993571676354812050085287620902975521785313648051914687671805555741680075379630184645753606064501268542625670688398569170826904819160369167033581690368634141524232846007690201067183835210862156533647333092486565685604348315718141873669855847825215196623125840228899250310809978044100481125232733424617155914057548455742114858709247379782104309649923967170154452137245294154399769130932711423197697044379939513608507370033880134493682561741162699764779822767829358514893790560310186314284651543783811841425208319755084398727483063751820118055457075008353219109122796308694250193435939324840645802251828763838103325594559365970977718459750683785967146476490662920872517491006987095230907818159640744049733519748277950897712257543576497006446736256324696416802;
R[23]<=2560'd84861649375964315574534703276604848906599343724610112110207857906947313895283423044253936180758442554400416019252901221443715454146489678242932970178078625063688789813374140501473168536885747187172449956087535917152426626059934542303685565884628235870424999475060697094511227702764069292123761917808363076897232550698739546972055242379422498728026497984325439997061605980135048705175467175388344528034510091427070149444538732741170395334615657171930010458608884619431744777237056401943825027465547296924129238512125094104360319462851844596100627443207692591363773757975638976643957015807339679234902817388390619986385563428699513292088636997384125836205330879424183176014210926836172100418551659552887770620749017964850644822342104861299940093626832065245436954634494498;
R[24]<=2560'd57773800423977286631199288167698527425283551472069132515992267034625772758056592628731792675974686172113055831683685587774018553159458732493094908281600846620034756432176949005122154059497817673958975918720683860322946254953703997935441407175043329138400457506631271083418840576970037424985967255116393613351892478351682228223285393639873422626412127685581945262287199940436041096935925477859887686102365272739176599785921608585519187781364394304951755167512585694166330563402125335118914360719196681938222226622886784686685398574786188453559404132217012229120318156560941479976776659956047868907528884816397743774923355449185663341893307650004712280096539471137225344042955237756424188018740342974628325423784776236655561866706258783679791095404379028049162181577679394;
R[25]<=2560'd86660014513199332527338525956260624693852715527042283708600032213176010953371552011717489775079219120796266846697707884762927750683352752182511547733394917588183677217844803845682068743843616621303916913975141258559610146501285186272014604299418773168730938210191341330988390895648904522360187009963925445061218318876709719320931449359948747999285685461742413446120894580288098663719170092192512836768230165079025728312889661182968313546483816946188244649267047924962930276129476569706430741900991413788656825941306582278735878946625565725643594724730068437497830119381134260595467865487712671162357134162070605251203382088183327784201576019656910643433882922222014790354693698915843055834084067178326181765277591804611848613557768124263464470971822435674288525162979874;
R[26]<=2560'd86660040339904447089907176126339298658372385550005500412844907312321895809690773594729787991810126860132749379633350250610523899379677833044574233793795125174668865424858048496836108325384418940790253154761309240566234132550675206618642041830308171867430389161944971336735593916210132022131503530537889276640071219741698132106585619083033078011939152519957903070068979415213717612557968256672928519252437178561013139846494255541335085634657490650874728186597025938793318471802674701438713479970922766770069316053977301031567503364609443192865008274147269627258508942448598478158278572359056728706631591557240080030986537164228163400683759323271928779255009644467443410983305858645561780584692941748688759453146918036906572334709173412634328070033088993272005854515831602;
R[27]<=2560'd86547644233906525683987586255959996178780177997147997872238240032073269924095194978006632401899283121123159986973669782514802806617610392338429356188969010571405452728691543893886078557031259378784701744497890552644424698074255220202923599241055182339369292742282041704193838968282107348722417470510026363729128538109701390388070213211521405608743445275431893536783715770969424151178325263197093878177645772979283183799834511316411771335680431246572852585309424200902827184539073956062131391100994881389148516651124884593556520806061092836269099951461061547986220524484233583170111118780297363967311441660837166650709627727135236239650196250340110051823069280071009638244155378367711833864098072735636665017152485211566547812428152915839720452697845936937640251913020210;
R[28]<=2560'd84854652053934553616298397146624536070538405817058795791924372022941743820520470230941590271712037180602919722013743340454328164096577216058187903529732050798498586634277863102569602142576291516451026515288934382451154787808809327755103774427980792576872258156047822403159640862882035327291064441941101412182420772980914398086519994979424008127860473672084879593065895871789924935146406586154777994941426366353735256351612948067531739489928591117718907137891727967351293934361974090100438830448416227896771334931776106721073589421338727550823563227038486511103420906199040018121767714967660437023136383361959210309570147128873153967453498893275832288057580110472253007465240434725688514733755877197293623892297599257557389657279158212075623668066763231393243529114427938;
R[29]<=2560'd86547203465285291722482633879994214875815498975382692729280487970860287460701414385200255970318623556746334272869381669311096238224468381210547890770423106354435688581003206258407953893488933786378791751915781472531612365244017597544249648277442070230123583307952948019214605531007597840715936387558279604095131424961528662324132312998631503135389959116820519422192572640471630263442010329949258207701526306317463390685335565874054041007597969956740717950506839656760509799215976725775922632727885979057554479034001955848623026512638874018429794958727338960576419281895324545614036925602851291897515804428447176454222114615066182882099044737877142010984915940204950536035299599612153072355618412392530042050399408658175791155816902537636026998207822435892485463037129506;
R[30]<=2560'd86660040339930616723341394790270152571184390368878512106172621765721761786334940882317348557350115981369538283328281307380971933914934572412019315683515460323602683126835711739208266027009483980063056403761789137044299932557788435826725385959496673747324612807970047750311784421496086925726238433309531533625184308966626480117925629871939538614258984676207805307644116444641756444329058617013468027523616568601192605257497789952848450230756953643323492745599653218312302393190581004587989248981335753017744959379788285806784946726533178761221137690711679957573770373013219357439161499594901346473285352103974364907452831783993862459954507223018131790959681413478751892490149539995229508689724957635794938511251978717343928600180224075707355994505089151502967251521450786;
R[31]<=2560'd86660042054983714243434959341365726246495501958022391305058741483538812193193512051140921299861090788630797271441700407132062652736259783848185445206712890924420752261136589925011526371798819243587942597496120514131354469309368529728818924387321812522608260999913810195140623009015812785977759473158622388249885673805556821446548211834368271576699838533418920514493519830693722143502965448998635824699131719201738384309681366426356354838822652438158917655932935060919757430635569367099944752511663786231191592030186867506931887112961013482100795520886875360160209863299745370046711447841909152093770400346771215625321707800411605177606495687822059067536051707443892351518632099274447971843916585869092640814524572477509810661777545549210451381612593390039786637906621218;
R[32]<=2560'd86660042054985349471078990978866873383091253928810700187133553067155743843200631518745500737262686373512211606600663811041295368135079097879957475673853053530199190497913877777104499248986550134855620124242746994467879621536033113987131746722757912166507160203623231330756025300266536996397491376234064128643431893500187293052189737704638924212782143797859339400465394492457790930067517994976831619134652290051505460921375358806983168229107537861536530742276403770391883848554804535534693160013240732440632153859148089486517665037450505671347659432791099686377303995985548588682448883339361870345335605661918560385387843864809000146831847049702609616071925845801506719456126904210381434281977166952342923476996665132398827404022965848883340509063816712299970021253395234;
R[33]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190657397828370163498723164913685864674604617611832076045901993997060241425768530503295962087441676672526096593656057675529032768822325345317787245001546690868033476231727400250427677543031936970352614325898729171163338123081017573164312718840866067197200331696042156170747968491170799849874707365393818741831059505494822523773896582561035147031496004120688104659795679187778441920133657501682062924203244353197531261743320598589302545276603401799649678068001091681851430885058924638923118150984079006652750602731440828566189645072263058271840641485688748303943623249718046003044544140568077720876050658336538857831623516903268377480886996635707503599997644554141416005752978621187735647620856754978;
R[34]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190657397828369292234014971812035646943822631590102383456438229367811963837047098782979556255159641393552570655490129934526296865439669799244866722657119836841084276889479123542952554282470385022152274795495621957013480389299800462920665170810699985243856780458223868360843374778163127160565177397070711106698505592927449940797414710756915765368760968703584625403297349013717095289817551422575089049273787086692426910765102735892019283623395926173089909278744886942519602601434478719990081749655260981101645184836029094194050228683761617612029284741559524076190765264426240417536067503343686247937430731350027266912223302643804182428842464628197365534632658852519579838334407258754467459055035298611;
R[35]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655778510202194070040161637417840900771471126594280959895654037703205549443451705331734426120302890038027626411650512251466303380351849959568248800570872694192159108235665223117982692034753284865807005281431807393147686334592744165370486019114791506275256411762253343999288511676827592420567772128568766785968295406151420415790795729285100265489881441019662675831910331779263387009743619300066762956453000221421940406872330379884283866249880684697352142141649249313444657200737042199370064025123557634707548023007465950754730725955012173166315959801014856087170437732410772188639969214737505676321789356282994820385685133205978391940304285333464365761427757983256176804850455244240309057696563;
R[36]<=2560'd86660042054985355860247144599026105825370384862450713255366273309420535690531809473154932743249057817960235194511538639483657108702584117594483549706751669993070060604135443235778016595193572530866041647824603335615946624991648011946306688776333337586893825044884325836406083916308991286584354641722301564662847016434433334374352514722325555239091441758688041587303661435674280792999912751013003971620549902391436174574767265090172318172955380343109096374320803588016649193108722850005635171263569617912065571393519190174976399184967855484254137357704749615382996489953129488088395423301599118179602198627141036077497085833835722511209144738720831045174562152776435381936900858090572942256301072510553897862018364809863945259366808264623663376585822018502469380100797235;
R[37]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653889656877323188571555612547409708236825627004531490970559363074718354930358376364126985645716118612110964145874307956049559112198443894452957986659319575107696609302942473597942669599872016311265148867229023005173142254772751930569000003825840204532248012810675726609370890294128222379096465142468906017735078404235596041513610336176403120317186255558238468077373612703401185314589231420607657466201681264232437405144331537838648832357875437908038388363570647727130423233122483543469278939969751277342360697257895316307984859161079954388547057487937484074020261551183868504359662321516224398030541164744774538941282045048615640224802838567082354516877311311343561195861857178935981929449861939;
R[38]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531206999195592058631515169666085870834112215180850712390801272940727870457721771369136713814219035557895172422339617333997389407243558208709928066636020987871570716482981243002303478933367314551356367101769105652767502163755149642053652315807525023245392905916975246841618000391795168654740183356848483491110660055349977867276867265485211830769984595523755878866113883992969540578929834217104591833860336645959151897799803041712681738528943294636731407835904570705479361248817178876443015977666559901284481937915382242958028520070787908597641591323338589686182499710885422517499770322137144442249643539449574790018369186665038480849875047590012558038448088104105999938940218063493060079969658482144051;
R[39]<=2560'd86660042054985355860247144599026105825449969542042632900029023092504966583652700713258564343580945446434503036217230676100177214570808110423548599902692897236229713371170339198121667546392903080238522631668676183078894976247648345234481740751658215289813668522080149862384027219361491548816237799294768246870093499258909754380271744639050254643749180999996873876795430651270530153152125106786698856905484544072267301506091070179026141025424573837248111327709615233682349410074304490502489993043075809560734034023659792066176487668779371481291609180005771713020838670742115618772734180585023102026930464068158579812052234981384414556401660094492808766172282087665252745720022154211553524721713288312055839787382764257214440802956844999141290532693954263320443993017496371;
R[40]<=2560'd86660042054985355860247145999094595491657999583195198385710377805869607512396466731678987761437164972739107030858391033238520402439539630334889622473537769223704632270839317187942177018404210977727094424850787920253479721927428136085572251020596373980629949971442245146379685705449409672537304522564597712924107208958314208419091156163789979313585724578363181082249707468828388402274707269788218623638066568898142327029629448327660211516401922854060996102493235449118519130297447045948581186117849278097339921048144617437041912330332475395504008331440676802824937174923867845712331137281204425048898848456099691225611922418826310914538946403218352038094748234235621365429995829856841135583715497922842648762513492360395868381273425084582397999893444004480391874140648243;
R[41]<=2560'd86660042054985355860247144599026105825370384862450713255366273379364933412339842983667055047579406082263711460100440995334376837721761848840631372329508764203044248349919802125093496978063216703683188686996590615444302333877479206426108392116004896307220607487467785168437029651672268191249678499342200570378707334526834768521380778250803137546874274698295843841074750359029668018132410204531675088437274707169953899582139330462851165060769364792714018188986665353698532431930660166289366972965911796335904748989053243367277052308974685592458146172124511779449724931157260177656609321916834440369489465644343841424174051710438391100523786656589450857221135900635791397372221889590987958326028960106638809298239411399053972428134495899663596034637604737731530175510950707;
R[42]<=2560'd86660042054985355860247144599026105825370384862450713255366273313808258124961949203538259139998459702056690386339957481819378899749425672159066314793457451577240781638063008135621124236601545533106135810918564561510481750284939662457173114619262226107534778546517588708549864344255077008336752270680402330667102514093759456736893536255318470465215786095801727285610237541274840831226346291160890977179416461971452103978732218562674825598002331744350861507771502234248922500679685876761707952789841735843590356453424711021690306577722269957306366667617521910324448240289929818976416294594792544912317039349286350001951742033091445988279211328987374403734985852959453466087757380391244541222510046771399578014182344042589037074529554947025534796527809710348910537888445235;
R[43]<=2560'd86660042054985355860247144599026105825370384862470473498900560383790969233441429082679984810915182786798554000589142097913456665368701439641228964520369299944441966372142316836296012441426454755047847902133710679288449747723865415630375009040572882694667339045376782776900775377336546142151578099265244474344423257483945124601322886754020219466213606640849796661959172891400980485054038055082569629271221272748396409731256653140007087843266726902800804163647533299589847174360138852882496309338560180578725218191789624918481747782649190529603761616806285352943683587575505893915895564067541362571991386245377393385684093230353337641840168283962559436056695275959262571679457013796970412981947011218633499309393101149130729914652462691915708444771501502375625706475565875;
R[44]<=2560'd86660042054985355860247144599026105825370384862470478022761271364532961295257704729221021131612876770568028465369627106275238964448085990526283000209666828557148346999043649916562142048044789654538224907986114647718881169296998646297860381251367123775011475464341201410632095235216534223447957421663158619323567892975855817761605800733923137795239453552729717742211564987090535939419737951382539239862305893331275251186747432609265153679532732664258623524602518288937567862975673841714290405361197961318294155092667997432251158662727655910938819925580958746769581351758008426699217326433714124105112264325629694703848473695649774549596203759666456702441016969602176716288397897292071638156591009685350146744363269211632687510518315374964705984813915055130378960215683891;
R[45]<=2560'd86660042054985355860247144599026105825370384862450713274211128025582489645378578319359534944713072904378179078903205061258955086550259735056424359365807955694828947394988227746318288296013831340056171385161032690446591086833733016052598612922586478096519079627263377138180034100981624266389374193185674290954278371436418280041886491533662734669332332843602156578019197760209213695048587015404418379889032054199514946501514280483504547551688657794996230414894643074193333402105889151886121777962929599874127795621299076530964881475722283225284633189595220600366941235274718933372591375418800286316537973432950665001100806337831008952117972188780043702087134290044747031669105036035860861870819030368366053525311671557114886335727124301323014007162950885173638800361075507;
R[46]<=2560'd86660042054985355860247144599026105825370384867490805865641025949292390543496542608523677042732505848431334203470616109546754390498819825304410010157883509087011339056074816876439722622183531849093964254660698277164375661648826159886665179276365371593709108878499840102591708420057386504341744840850245188437196951956872157149438257289537378380712632380707195147273599421874549154142470815487018034175937668226408235301960324270534547946968069076394385630547675872100999215476757991762832086186350851553094119266118993156366870451846785516175551707000139511575659382588108648804839694878211496723776144920421227951543153507797380487212783117439520767903005458152049019287194550619050955583143923030579993844353335724763722253481270980688773063561467073665335192823477043;
R[47]<=2560'd86660042054985355860247144599026105825370384943408430996629323382492495282544801194201851668714806843852744017366940954206200390443704160354779651618464754910635216163852899837414858143995145742208850515986112831337224936263793528561737911572920611443483107843901638810984096480072664422267815555037890594797856123363715088247129490780720765788864730026535740616607630693950827787237217014825359952846254007398458708863063677847574531545788037542670095583546841426566795013229422231390425547814050846531832256637360966494161967215896236077316683277200747917986919914283282408846602797433286434172155988982326018770133863073202957289477562819910090832348621666833300117729944133716148863683519822875662727759964116161129879766580796007493815022778056171230519273022763827;
R[48]<=2560'd86660042054985355860247144599027524485315178286342881503313359107810210882286758420859735697677702715371224890610223535319203454168840169112673762386350707273111350432092416304987347201827089904471491364658274077861817454089395882524183094291436050836282680183711760696597995966985593914721487986095937378218087337733653572617363580878920207084070009259039877067514778625774367786200657459040548434018303378217066407130043588814946903441909503802525058005524626821660779172415231756529639535750313109758197850846896479395580784424784713625376513136954627422151127676269690724852166141113423351662884680657114737890860980501209577442373198134926068421224862036953346833978796160049354664362283794907694010061503455531824797591035990127798363773683552556536385966336848691;
R[49]<=2560'd86660042054985355860247144599027524506962230641077776001648326611426741685203825183219895866240491356579364002356310457530253206754002034201795084953760802861847321973770594245467025372329167061525642166234772030790923171770597914075954245251283042568345438630306915012870076946752784034073795315032882164432373955049482305821989331497146609125064748101258209444389814720368290319437971840993039842318424156272479663736966056321906409465694773634595308531499880158292938803971613789213477994804496055463425468192591475648377098696470188963804053865660514586640093550548203411518030347482601235432633149441912027233402039771011016136615960318880495174580731092324094465408519040656680315091298000873121178135433015039256990662494407219162694537064275278374643008760132403;
R[50]<=2560'd86660042054985355860247144599026105847101997153654925205710892427117570098319315596922880966436658556203602568488338170605979333380608179451700721505915991930054063847787019275281673606709554753470797273430339037216304662475378842362780203642370176966883101149800876162682929584475535753010433387703693358721346321035763267034940356925387000284263852583348623457456026286321765281183052856146302354936692736184072173933610663857115382750266188826627324985550079944329002456042464968755635736407285281646715129608085335038708070275193893804650032321334641530685827152357605974854374646979487930198873827595953867897952437942068739996765475422648470884018171574772717425157514903854447332351540395119680025262722675448350930966917020537781433578795032738975825158611350323;
R[51]<=2560'd86660042054985355860247144604495123384860933153382920155216575593502789486967465264227853012545893953269379804173428824746731646092879389397345441214307147369601249388898420866646979295832034206543994916270041296030163502357390706978124357888729507742824898009660153076811353570442906386252642132363704161150990411839345736769691335259632661407369119069733095904493859186660373639578276272661163412799110609197763778548570988250243956641048463053518528351283031585666048644938172751595020307631735558838704044023863121331103493391343487128623761335493384284380236015442734635786430243668498849295435071838711638336800105877490922097339489918282868315729922358719226896978518719485605035331404210504104529273789977424105193141238498647336174109196122448174399984416011059;
R[52]<=2560'd86660042054986991463805219899333553356456294087975538600474899124939883873852140346898673950175484734079463223189413310560910822457714413521657952037128645427440649915636808286721332995644758388077729815813113589675846957328274038199215589030792138397033995072804616843467602630128790390802193732825610428263833916415447683995523705308066239206226999073244731865848394332097612273973313519668736175493304099779801208710704096063921661834108172807280758731072338396611544248795578697631218887496928827811482497101076342881260008470924937979355467653601834332803826008580338515874911443543031784814507444436728334860296965371920481832422506841410554375371111575557131789861513575463441223075141977388832547188933489794763776361427705968815552073106618400083705955089593139;
R[53]<=2560'd86660042054986991463805219893864535818617753983843458711239995000166463410691050226424640965390937583620509999166887975386495656051557951067473704689088700790425229100032446501941656230427710592509771301369924363378125024648905597026395882523611836979513978352029282219226912677707927958154458689806896236220049042154549908614898478393267381741628623672631667399262893511034890040314930328049640529410515007244328798690970184573107682285322088446856844648762309041650930132398087020475850387101119967344844681436563728623247868885576716287782633429805590421808804993549269743024809139209312231417397414810890443137748042645626721579992907423733366837283923276772470335799340962712143880758818951006041834086288958174774794024735270057469042290345621081466780966655832883;
R[54]<=2560'd86660042054985355860247144599026111387384492907707816508030576582809955086093770473639743009215524073147139389162198128531331119567814373080521468347892160076526446537214356146979136778415577692839761748384987107825904465224524085871578225816709697912033426558106741762816332083837644462597280168705880488600075718067639077817912973437930030548867433537337033799966744512189604075349853968188374392900595145268188272855616970093546179583569361216741486711476729841546911592578882293200115566397109995447951432096322613839536586831820687622558547122075673933926602077743939834559815783789862825371785120486070110491353156011248671307594540491744249915162375342339296018194387121746917033812099203655543845194742978772465202081374464788743159640659153893502093655746491187;
R[55]<=2560'd86660042061290703812090662096206953526977180103761846843533160057564913533641316529548496579156688830755124329601510661902801047760447210681665988247260777465487606824949932595372924642149443518627106578998788849605093181469876554280374573284784700299416528530079985264839193049590472130274831951577290772998277167072280606438764559573910660447587892763065222571527421308907956040737989018421734665043409995365839191289769661585241994752983683066727102788997129001486073355093758404534685433402527420169979543007055044889312203965162915823327398837670992921749413665310253174612373087666885865062057109561537193768845469546789032153782322884708444665494402461071138206028322096155904012922279269289564443437046260008441564542008038837432609017077848413277335270869644083;
R[56]<=2560'd86660042054985356259661909176670921900115671537150718549270095808602670518788928195169449956380894487600080751486788342617758245904200992557493550791932161484308035803435780493991116927045874698677603486310549199463769060127472676929857317176612893656063014768373840337324383339618783424429594887890233992884772378946005328782081878853296665804478423301641872293730868576259170384555757057537839257819690251970432187068951483597327585514916505539831366587965148552850577021937415947968680466418474225834801640513670757040475024349442711756535462211883383994090760076400791901077856248753668439177350641282271085223195398786206816599079760612456305843168192105475398161264527086678505806462632499217700732930082085318372277054637730683392438148624777202709706891502760755;
R[57]<=2560'd86660042054985355860252879279559778961087294531968257063724679241628012323114888132273903295990674863046123341897961833080183342937132613171031102060768080241827386971198245589566576123129483677216594685414317703711532600789893343737014630818446589617919513375000112390020437295901385048634061802198815177529635876109444704902548996381388321640935511219127909470443392651278349485780206812366966945686557360670887503147811313877634767086162804086027575158774564167259667568720575416103226998746804926358167376219354288828678060705500316287378994075039513296937605029108578423838500439226964685175153356965693134495516538805021541726489637879351885808211500055129422641272967894666858597989158210420909386179098055717663291544007946404210124201081239883368011905776169779;
R[58]<=2560'd86660042155872558317473476393956806370006731699731253985208197846010288411345225679579996108018080512303140477682782058501029414276750142769240773319352283307532336251034764920748548727983268531417850737167659011810345720266418825328787953469248244737426423747497510714248573991834117154992341832256583937645825481032132361139168968619215193172805289827615271606713750247327720680683147849334858061898232072953145071514886973513541726206369765042542031712209836605854604784077389073871556150287037640114001242313642722430433731938148171270876078792327541646904091733744988891997001743160383150450796248638961927430879221377780893503367409198723691454358956715284061884594079762731951380485463231996473959243293848677835950508036992344012393661873842403658677160101753651;
R[59]<=2560'd86660042055011525518644808357159509687291433515085964417039928896126589523036157030202254624748351347726032316177712983415544815224926344480181451280092230480513733731852473090894348689112160045452570364983360406450457174953985408887907607321656775588617371753084710375378877178011321580925218561517507530380449443033441978121556865986133151210082691428903715907926746646488983199534555706911776629436604729625426845641605609387902608117295416122796081883574681407109470063003396778576422726980178113391364287138922140614816627127566105128471889545984170149177091707221802971952211709231557873960703944370540445142069041198299026618222883561103774516458185755624837808775179378085704302382847864104624506194896261342230005710652863813058352810289416753129021733491389235;
R[60]<=2560'd86660042061709418700254420070364753889614508357520476624721847807459521337465306055389381869949376590007380915637880869426450037489117619135789536092530397393851945932863022784825021387527396467559900916438545666252329053036781639038463359581704323711559190413038180880636256561073128020105037350598327671619805554752651591679236676555929692944556941839183913375307598826956062552907148929684487485586095053206010103874629023429709003614237620274158062630924146955184024662835353185610528585105702830476895914802121256876289461022881976696866118527709748142146797670490009332908599397334193689830455001318338486271207303318949634446854851412072834764067280890678919137492267658627226670678203799482992627192653923657606018274089623855056897318758379734360346225072616243;
R[61]<=2560'd86660042061684788434908905394581954282049706344425075286964609985642652802841224492871943418896032920217549067834880581168342327028364026700841481509562565424444504679750194453926303611173663643870951586117099927157088254226142055044924940080892482010876829113501699527993612513785354736727224336428738218836522903515473845347614013102648912334529848578521941485655230499593292233105051707831003364176168518680666868929309106955468830138409697890405768926037839380741507899051255828496564543604864800534136155758708991589921175442987352028988051086685076336849536761795789670665990635151958961997599890768867165253672411716233320894599462567959509898835662237083481420850656800581906291520653850831730768528997330294445394728776131916381729126748890625332872406681989939;
R[62]<=2560'd86660043776739430959049564356418068482798466267026363645601927613655931042305459210632621960045613066769626593953648692947322220930649655467775417323791225067833944398209637963838618216928797479491032369568743993350634981293284067391937476790979468979978962684723201343643735098506263324123787609210878912941327632287396887860931845872967156706196488095078673188039453156455307014089082197659108601219198261739905764833834663395952373891932466972639002788457767609981403853284278662892499114008624106716597183104282282056465016295469538830356531480417950311075682933737402319863163268435928323948760288777599869566816077748920891144742944538657102139917151964715192950054777411601410011529147713326102333381581204182035410436375916063186697780663278715230165802041946931;
R[63]<=2560'd113741306912222916102515745629827062024192846773927718299790363274151204559617680307635052003802028957875899325639540199376878760337092314724543667534944988169781894723172922937953579341649351582081891973233548183540508808131879053295095116121399567394249309717907159171800997128998960298614170432743606107529604609252205846070857375295591077590224406238376339356905491272859010413650985127707959827791231728202206490056528592517276373696812171830955169620102624587275029547663361542814339649378827065888128641680066336429917062427401531388847564651748485690726477909204471635618757351730018378467634390693169402235337565915335390789898219718563461991448867360983494256492174345159061931083291053766698616648565237509751676533037825122619104559483733742666533982811927347;
R[64]<=2560'd86660042054985356259662291307887107396128118975143391241736401332616567217132706008379085197971092225091794459131020786618339251093417034592598131674106841641838066241666930693489942136868867164452742704985300188312826851427890339833782054782468361844056237456371254762593063893246375696235840959523580585718604936108734862445531279209409324722263224928230836226165077729707834824289407046228829047869907569866137238683554422711910436635649786615326669203664097441724607625170472070983221933721735247090656505859367163473587248713567777977045979324762921016886829477407717417150343450162779919193827212598676872341666921873070558490445669464604127110581560391151121248341915635229773655737033433064079576328307468212566400469204734422694491056853570533748968307201094451;
R[65]<=2560'd86660042054985355885302346157210501844775657980102160230944711620244891574782170445457337435667824447536769870527047746072772298950173304770324538343618175406629605672691825396395552723433292116446955230933563664624532058050881568273474823271552534066877326005776170913892097980344949350461930991226400763110996940568016431404869062280821105230887713921476840664890142767459646825802534072828715111848518660335137271485924097614897905361379214277415776222549491868944530959290096060098504770398312182178894899105877162560741510405556782520067034420383360672449845755753442945240732068536820397947655991897628360200889698728701112301663438875590596484126464095259526015836493616443250786031307126692549331786140629771966058388813926783172721464675855753649771304444965683;
R[66]<=2560'd86772439875643829910398925496118397644980468243653935060421426429664515755318921277076319127852733209416501908299711696988293155254046791612362417364905859213671160076037874792454705424030141217605867752265571596673279091388578242339904622948807226508094172374206979659828816627040065658386017964171778203595418699048120666526273722179861250085521321631827114139636645351247058508734844328660483161103400939613095104316402725829987722071490565232703220131471519471833742619738063736289713065860285790535071803837714794729670655540030570216515072212301518457315840292160111705453505079395323573524695057602471633360235863757830713292934803046751506336292998519798034545184646627532574055541187515475645427487733407338401255389523827162851798144718621981054449981156700979;
R[67]<=2560'd86660042054985458087035474402317333893402413326148309711117877882198346765958918604498883896507696349201493982411126336264983311120353329780628280970259522076585839190161340196052780052272702927357595588144135085971782012684663860040659695373083628936331308657386616372736207541477925778905961528594554356131418295754555260146073787186587749870047183836210510475546928155366597090915605920686847072020595420598586263036594295558097469765185278054424251982078462968110031641042136147707119349572170574474479463774153810344382224282566105999663074957271343742155430541308348270187540261280617727712473453207825173904415429569151288666051404525816947021551567824014165303694515042605634583345133962460045887232992844557403372643903270488555993541902552633377734498691789619;
R[68]<=2560'd115433884244441914755544033004845702060129319655254954636544497884684051583106755871158390810372215853380970608756650521416183995433525440994104438595399282130233703793830956420353798466302025463956049202229838454074693887659010366504078669613136436235580922066392902297560067525071717831955055077265766172131253511771424446119109971706160633869443482446653535600584880591978119114706555859493649384918317176053472624900862214219787646542041300985919338378828160265584788822067836393431602800347415109408073047927101757206828229614490020541130336169572949714558359200679620043118713202427579325246095819772539303511437382544593094250094260060501326831077326944427596161439949265494841922048010288207792184670630323691940858218424388644097573714993642159546973423173579571;
R[69]<=2560'd115539670428615600854643003180107845207537251807109916959732824582815566427271395598547917968864052544793495271479965553688657493680707915504256453562814814528764779213603146567188314902671688873704715581623206600089056958493805583199900777686826911379607969289809338350955768423324414095483759172663231294763466140149232149521791089033449641457999281042250281842277970596425390052440037577276963361436278081065153963360882902132244271911295828693377491363199281809848481364146097597738230057190829187580323238688326697363967124141235999340550032970368346837349714949532798935931468183337206968590851195012267052177956373537295113380167334668689875254952154508246410313055168774522490398770138110060514982450428959371808573796503773431888037003914383980739999172400460595;
R[70]<=2560'd88465018822450516566516897040131128408816384258197055583990176216686477470385370003621016644500249789371797109528084905006900751745624425949615908663946453703242100018982957413131577802895784847597087230268427118699766740439322277514110383844563647734773164824272915508756613062195675622890233367432279283083085419530208290818062108440640030640428759748922028594632356258200438266006749952874221193225130195536651237454981467612240613469685944781973896220742725287949990298840742252805568207174638651062710709059300610408109035384781074283799409500984450740885940460685907050138570707760196335510137696179632695217423968404565979044420463618092642358165838716817111870430613006512822765288749008145716514000045614592383629683616788115758990863978296358059321242357543731;
R[71]<=2560'd86772853103345916837346171046543093612277487282210449760258829378529702122627592600945798700767238234642510743069547913744827939432382791101947639379330579493455350259506643304783041685422067580176592658078529580032018458678904275980890868995643142066568373746826726119462364420381808853944874233467748169486267065731712377268598841991687238001512177199057803860643671163718955167490691469905673838665826197518929478764577362031340784773721992129964060395053934854466994102806527767249491025855903969578238283646303594712524274158477855760484397457622333609950670220171989684426139581368104585328069295151173431262105032957322796638986095926593965863552997601419274785774594943717503942632020494499642253310261930603069458225876940701839313309784900960154413890334372659;
R[72]<=2560'd88458847961286593167586226609893460958720097506648808405713204722629120778463442721518952812420090890841436943606901374959230399889008643794754441389226150310001042724382020728970456775761892270368502888426454685644638801973023570803934373397208636922408726576874726566937248758211374880677894757815368992894624330278529725462820831765634588183852126291221659255478065216234023077356417880213390529624413724351110640890119861223924788930276561942604988408308097775218561932252421346349514346903456813526499292278184437378221751362955756047027611972226306643760907229735414419198057581988809996000078088642149349059935853989695728427486294428278509551647620883268842474432046037065570917242873907852383847893016385740220518285339694132229022691702557433345525409731785523;
R[73]<=2560'd88458434626813845760385081100673656115354865026685256443379080191129654180354548134697886455307814339074762265986201557313193278218803681810795960809643589764979270411579528337144758374546580327395197240779562147395696332979946926514586812151806826595674169909467070013556457990123073721590723461810810556114495399775155241687686308197047117485552765944453710482975869719850518563021500195142752937966046517676976068176842234621519392573682186856185494619306685369618213145239320360397891284647266821866438343616703927611165614151772573755600399513650227868915560045888478287178976106837505837079812932979785064707687100102581692874605726911060332628134814480451521446600574048825448803418858975577637392074241755828835027989774450130973888309188175418921914057916363571;
R[74]<=2560'd115546307791337021810780710264363309586168621823507030534041888172833681207658152146166617857106097449903827982813714985901657893079269582988416713806073451484736686320212060248346391874255004003930999462437265457869584657266525687728344287593003326928159168579087645391908330198872592019616990057629039958439426446964578408561275762289250530717223718744823844775385604513924304526691008009485981638067985493527095413455493497821837007212068540488733082189801394910079994557208587339651915639641167655114128598657904071892110564564885259153206337917204218575636306632015687598601973939710220487803863248214178673164918084337336493658013995404596291125132701857954961043920002214057023974882173345751937889938689624805328144370959448542637918490664078508519772922559279923;
R[75]<=2560'd115546281964213288949324523725287038195812116436194190817975462262962644549633684176970772107285521921853065353401622324031650787026003469644394778121857159031569774892538120014661163723246837362208398052341150453546324960877193483280761124841687127378656528034096471565569174493655754187766946457586601008543110879275314694001147669314969676594712033102445336328052568794062091665789606618307509933059211516862228307088751444735584836066907845955699585503725335007111528534040691636316732917269007703572467720294644127583628097987883082356590946032776496273502373153133487064665797871116195662423460097268323936011287266556336251668015610467698033781458144388223088809393039768083475483537709257636565865898777422770538083273404865063148989794961586560187796737659974451;
R[76]<=2560'd115546695191496654577102573731276422593524994144741432958744638491782414474052740259893258282697512219741469268071001186629828487915473188561862396669655586644328922486121088919745184815226049629075064442977145140428397715499793282412145348221189325762355799621136702917927498877264818473900579177218367891041531346334006821636453025939521075987392287214770828027633543137147285822931547851468594658722011516174150089642091204563832960417873122410822211227604952912257390750204118638552246599322293501471574140859851010051459605426027009701203345490370181512266884265417980904864769129107467950891210615951861097221442703293319741740303486449079755244239345786998859315548587104382585857547479040827050629888791316924405404447321727653849374790617947307277971290640823091;
R[77]<=2560'd115440909108233069408532241032113690959029811735111577758859172800590682417351064641362718309402891722622434518926197892364270270351109678228120185681647338195171722347122818263978535131475036768299642782889482803709288365985545758514160173055456087517526748410919018361618552801494117802495118967413886682183090921937540812239499074019358920293060296805446624445396935781041559095324948441997386208570491463599045154986825113085645144717970545231351949789382564148863773845118920936562958808926925133392017094164704147007098170147580093353125805351623606281527705619942455700457079108439395871575030598096583958864254931006904656227193129151814939674435906390078867767231564172552243389848372749252810709366572539478083578200125297312527847478840487284135115113196892979;
R[78]<=2560'd115546722739561759969462250653374030936717674404759527230838407338386477947148468341457112550273291040780727707754204862061197411877253444857409417997011239732541484812239329959179914077275805698136295956140834589329686685719319716644522387865054752713945459234437308020983374994711175578297037005386304405000992209190982766831093824469451740223445438738636299829112645913130121151622852260971418523529298082725498604763769974599882516526441889201355081847951150286244329594275447823440524057183614383429963948914108492600426719860863600664922414781143981222059815408681271154605470586668979399266590901347670015466733512744392957287687852145415490168768627294616011053298330830524785981363038884641561803956973219404373223499811821368282624503114299528529967501108523827;
R[79]<=2560'd115546722739955838201736017003508257434755359998303641069551094497676565616142015403273461271889747252964039748628340121821880065251981710572826427443031949752678347249141731180748785257762203343334725748464712928306844004919169512435644332311121632789433343832090879639707579241217630013152629015581005944983620500135741693953834502714004888934545310889017470340225562701129951469677676606324902878992653177207066746190943034230152855037836533111637183381049977195623297187597202496613717709615106482101053132796062948744970311938163700178155937763044354733757122309895303843729627463977421679299464042595742117312110743043371591936732248115285708226068981438552579697030843162071766053976267316108554717087290930992345882950436909717750485501463653624447803889628164915;
R[80]<=2560'd115546722639094907626661245737804909532591966489781953084988522520572222864845856601620043491769758046278638297795353737255794604240466418343264751725281306521479364581765221306299608273170082722876331525555328207626501762453420469461543977334640100656643504890236585964141730521417102813553644177418191268038085420616886341725459427834928812510531129022674912771599794289563273028549085194336603310660025998747138877660475630809890762328290397353389498319669392973592640919974637355747712030718785870909130775201301094332338858540254644848166304599309797193301197132738002109096458674974852587276715224521188178491869206966392523707450311227607053647274219020873779213780553359525944119269601041375508583437066346292772058810941534049920698781146177247548220920000885555;
R[81]<=2560'd86772880651411118042356841401889421067330502551073696255335045086054605835356755382423693666379619922014936694799007400969445752373298193184674309332317308841794651098074706250031436859901107108473771182763113383727106460607201688663867874338586330943876970152824672763815484928233464655414222127645441452300120575414264003196335530427134053517372567682451079334348756323890519344323877843221300835198017266043354492921016106168743948808404961163608727732044030608428793478581220306846575626053874787450662937429900890155094163853787986100302283579730910700146259228824742549713000833937261179966475673914433062565669463281375616531378313949841745352354885005188756673977057621280339987227834508003209422679253782388712785861428676063871268925711104540347082415644291891;
R[82]<=2560'd115546722739980474480329526131692994171050579650247833373191615019254092427119445517310176276560891546743632092093093285297460471957598038380505136090695016110329231196681510319730670248312049778508711846805380962608222186120750590090759019560260036747727992059516667020894636350785014329245056643182486752505467281333498880213206581423687913280416709984382189596263465577943307389727131207841117367794028895674942581888499221272597476951112171070666938704147273405896324892528741294379418578395477719707866965282037934307401729339777463824313985428628216415009830348111539661592359085508868347034694030245697405022808567680052191597023986699605860803454159727551415786112431110464776622394206673275619777240706882131723136359522760392695723210934243806690037728191656755;
R[83]<=2560'd115546722632789559698307003600344956711552730380179684853867416640160677182585550402986558765102798430348498655302975974935889900171084812923433740653861655268576435497148481088905145795576118889098774356629885266987004743029065098611226164816719865701576199261614524345651292095177683408748358318177142988163880406505090030134346665875841569263558049920592589856309966928592991706651740118132603422198258207371392174339764892969209110016976108402852050416322714961852885822972098922305644467452266190343496856744582152305123538631248766425828071743637187810570657567134675984338450310528971503699837649795379077154365649158415770594409409405494930755291645012006958079302371752498118743236523765970167093120708980446106324188562886137861622536529566493538597792484897587;
R[84]<=2560'd115546722739980474480329526132034807767160513150230760675695873007655051263892547225604825473704876993313810209424888846869891899021097237122688469462902129448370901689052524657127397382164174266815572343777905027632394631168336019187767226608785058710162320946983857242986550854507095624842170426887561307795368280266674681447719904573561057305481797246622313270138006655522757633455941218644254198720074123103889468779781616381602035368768444375688870611228938057639185293321615650308473594546678547903954356191763530937084412744963914688013710399778657937251902022891184223941217750479217410692210184618722441273893761452411438952505388950513773571945520046608677100728612946543287190247161715159086299084557321793893938960584780368038407686634759553025936214008738611;
R[85]<=2560'd115546722739980474480329526132034807767160513150230760675695873007655051003325618910933535755320573574808379199379205032476999760926628059568277259571367927111757030014547292597294403259844586270847469326425300201400705052749329389101448446685853052612289783682089883639085086693813359716856365435355865648476312220880385844814775316821921128361409133133715126993320295642174301284851899695322679369632878291308452973354735448889115613884686904486279076429002027047458404692923316591844756621262174199540105500490264214513197336055614267812850171478743918822353537744577935447445833964110674590255751396197682986065236183756911453331615499336143181385332893707120153338387201667854469442813254529648540896785191266641125265208224278123980690035854537379058964365155971891;
R[86]<=2560'd115546722739980474480329526132034807767160513149935515132330253078634144980767869227522358556578761931483629438364557992920428504703971514878329640098936662197950288386386274955592069048049273126550595002912966996357685427544594431174848824049307127812078132197943135190335117955744973445939684014325680224682524603729763910472553639593359721390992480090438591615525260137754746361222007753170442248828528809133153621330024590212658336673249600541434531915655226077732205105635104810127927062329504875269617024218897683507474309997132380708231484771652947598801436392065017148481810600789017495980082699719177607018524744618867903517693653347731895594945438330271014861119800475692111153341096066910381113246604797197599456370251588522279984810689491348072000807496790835;
R[87]<=2560'd115546722733675126551975260100779040857778286802925929017572693996570925743012100892605849023547579316137181328429805206196121622105114828930292245291825525670842756428588895395621555674998289243305562824111801723012267170638613101915242428081528206282033422420116238960957830084757744880409654481563112318619068813498732108528237176182309669204476995215562436824158086875403236793702077412113898445326663268714764978794696499354390151965993264959044113791114988843575537440168675724220135520895298534872190657503493263850015581789518028448565856653437338274967229617683120556477007123071938432830126786583600363458832859516139960925008461372050122324342741232868878571329770958917450504036039734074910551667663301252548211013993067755865164721540222615944310897452987188;
R[88]<=2560'd115440936454945755581025183767796949002830262420274793728727853277328389909550471150102206324641010733420777309765417460757409479490560898787542382425964333052708911020347818354476630821911748612858782900190431809197250968683684198116805232445815776550931959671876209574141889775058271223768189111415335031434192706587925744932080121165943329462272860789889248806925685151270379665007037411490885357710013918497730733558513737938189517808493233160637800178501561366023193245251635478447923306159205930143444216653823834592702118151355256294979996613169756356266868069439177793016034046551588984137978271858425653070603823584214887931476828501204001630077753279468061098549998587914649162436681830052816964340606788438078739867700879988858607149844747169232748154285404979;
R[89]<=2560'd115546722739980474480329526132034807767160513149935519657299989321451544994279597442268315107011040432114759163771117794431124489707665092447732062328527125201011613521112007826368151318497042586954290815243422170630238120627428772259813048106444047674346164856050517890202126637330912956113488879538877091017933686156295651532484127143001348190715859477562748929220789193597015718357345931450694025060028758026248525313056602947289929125368950221277294938334392667680172923651481464810399917905648143484709011272122177543216050729053394850400421722709254071207849786473148263989228641620332467989080141636229125671316526669268709938463888083262083875246546216602367880580705678386058854493582993059614876328250196566473086790400857591860232652428419031183881145983120179;
R[90]<=2560'd115546722739980474480329526132034807767160514440199223063284829015232741743109381207115084245551490284461812829567083701948735255751623475903397324184796480187870748060309191323041765990221273236431646333906331843522337427904502597932970465014777386190628997154568610625978044862922875810648331172252588098602743510958379540967382055852629352487853166734967639121151870379775444749392554580833697697506431710091087310977158295527540397035920016417094506118747683535694565229978270594275734915551244526933373322157708231022087620721092635107506564907267135248059128926736562869983304583177732092985661834871736314911944896200516204080771410422063063137473788703492508252649637997851900095020450949796744322793793002089024244429433860699958526611220971260250011675264234291;
R[91]<=2560'd115546722739980474480329526132034807767160514445239315654714457295286574527582045795892392864981951282730967140309813909046289827255895982900747809421731016027386149839509354720351918455185670917861421388132121888838549041608085821626902064957801802130823403945266942305912448000954522956883824750345368646967129000436782207312187438805818010834205939174981362961792608852384700921999034232487571366721617168349525152081356015409887359477377939817917387960309664599037141410649456145894489271809351338085735281284087755118964563712082851089244117621916399570329598527010900415254902503255359441222908482064770352695031610908675284676177607171939597701901737449814023232751491446537614092973807625971623137078729037798357658680706082266804704297327367814270136684189528883;
R[92]<=2560'd115546722739980474480329526132034807767245073167305730277168628939812777834341317908057330522244299882100426894246954842433841755145637102101493941265907443765132621802504921296933804411247709529457209601730452476685002518090004936694693392228961031985759940704310865126460089856228762423727657649161077444908032672705242830059754554745052622732164453746947866126676387889710881459320066063183880108907494494407207492607453574835819701515546910908150877504360297428389496226887656980216571623806365976897361291705762681463384272658246682093601393113018552300155626127969731917461040913614770763784732859735409766636446068997260511728150610741895539411280825610460290257701122721879625485980542354453594276408595071930693178549484807520278809188281621207486165844633006900;
R[93]<=2560'd115546722739980474480329526132034807767165488482988723828040602644177878707693484547905581960321561829035076913330861309311369049240888737382203644851613525439239719332939034491975061053919746871998295306058132029258734070987497583836898914790808036360260254111312783358359373543886992682387782884339631473703748711559190143966510822175591603046301187003820293148580378532717725240728014649023098404103212417626119061263240633334079252660040393904666417774639424084006231748526588776381448808785402580764457212886754740208638419487403411683451392915081222972124535175246424520087309352933710456627001401756078853216665610684094629546253086997226834708827820820574253142978491185080697459488419982355199182112185578408550263801897359485604392797732564146987060861421695796;
R[94]<=2560'd115546722739980474480329526132034807767165818714598930853925161917235940977577173828490825478336596308664980578025390538837458796619209210749880825397011756114698910025979427872652791322008026506615675365875474273838763268146487472399171437927733859127588540496177539696923013354481748669126550641792411157459982730050865922983419896009498736568391909092659888102359226242469240298150433500616505606381146782673138844409449812204636357870083131673312597010216485956848779597624066257864452545883515685718674634315020874746311357270343408333396281253013563399579407550158755442832820629996771208156625769524367552254885729865788742513186962617938692839068234493483415785404393633101509922207175378876172709207017045204065674036423764283687746289842678320871176243346879284;
R[95]<=2560'd117239301686366907235464229640909611626777714585478885543984861841796100246526608587217789612380334697553239369725203069856406381647719925662112771961636012172549148947159257664692164890253599176622894888860767555413302883560725032384361458778814404321837428349247357439202141795166457138770999223154625405421310383462381198336146095537633024805827776284995976400334526400327715021987520154734151282401399434336579970620485543147316382260886186593181759072585709669146078737491143661985022991755785885661185717026485694108320571112540780853484065956280036896914936215457846779717050873561307849301547042833770897345287095967257815599727763994344555939640984154177929210186235897196418539620561430376407911060752580008087025436561583876161629545643492758281012542609503028;
R[96]<=2560'd115546722847145219605422843945967965334700497923310313381834172213292348366676753675077193410919697237697319405030479499143190657336878576568652339479800263231699733112198588583222529886736190744365176005975037684549316444622228801826092979977822912375269938720602573337913796858325867771309552249622639694765823940175219233013237181051884935358447198210422939012560603952953494476597964654955720118971760591409547486226653769984377492762268803146564411445125814724377676296314291546299106910381324310383918070920645222730221670011407957932069615652811861464825685287546657088741630515058470863213178448670858286752050736644514237640620688557905106936205195628555881942404319727479611446704126293660330515986210133454246611367396246825760991639581246160808901309230236467;
R[97]<=2560'd115546722739980474480329526132034807767160514364597834191840421667136677749563116878101643028990179226678281562086452586772609081356127322283193205296512809460151686158533332603986639936933669864568694234736822102810734228436226497852019349863049119496698375962585757869847199960558736117659995416338875230404764004978622417673350567124568454539381217555313745488912293411967216318156341592445044453886154851888323052826223293116233024446347115952578619638938037837349231077276349520101614219967145967763383576537263327517094592325833108380556140613414292326744953125237997065288066329577628846451349415060365495025251695542006532805235132063810564981033948755792658518295286713354695263672724008171034954924544338248354935106994437035024784058619668936215922855721059396;
R[98]<=2560'd115546722739980474480329526132034808093144645759505492607490535018219430356551449109780508415740113423485433368994495714470197997021355231629738858816017695786336462462627049574252664440500090710228158620003843579000229285046831243712902588615073162973938683745291183014504810548079294215481006072450211740804414130088095265028151995627082496574646383688364914842742363509446309576024534363452211057678368024614025840874779373644362177358745808580846995838706545344762272274427536056426598045914262327489291464807577700603159277487805894756600923041374805814656587748281666372701486596679234360878235491590403257036592144389447667103960042458807053978490220748488967895908924465209292127754029123186180229495206894092371003145050567647000008431127093061537577429997139012;
R[99]<=2560'd115546722739980474480329526132034808113597908414647371037991602900170213060117717930659335852179630532720298908904228234955007769298288550225240062224798463240731230418350483721950572565486904127748026986411020204376389154691030269433630448361038050655795032326293762812075205963493256871380311975130971851264663330368667658108395379179067652770846373717560015444393871664494400692991768656796525503500372063298405627611194144461344839830094035983680431523848583091744118077121234585008527396758799329498473226646030928353015018022739884875034557149622863754798637053068215262729017541344315586281559865891951052951654636243824460347309433736831948216112501261426700496736055972156617044292321891612896660660472300093713216310082471545232304728681992743650553511159219268;
R[100]<=2560'd115546722739980474480329526132034808113518323735055451393328835276927933484029269430565592786566020881936931725556268515992638496069618319878554690150868293213505296050671526628971800473999297645304959455240914839592511726069422654622378836566116880838666667410744014125324752769609852132552173999766124254911468560320609955001918632099749589279719642391572155903057397418487943241348763166633223533847423113283411335994489873745701388734477003793057788873532626183270312409129395686187435933096315933092265147549392157072460038588659165643430752376195686068450659237792126653983989227141147082207200402783530527842675998328880379117726270642863342482886555323311254447851360477930688389470153658693014840967581318647020287279951226493406555299090648606392622340200744003;
R[101]<=2560'd115546722739980474480329526132034807767165798075123292914807376962944107273801102489161780434352513432695057102991757746280351936769700359561645778029460679146830904741630354040346739904212986319031305680079464176356604911885059613132774733708741981582782925306875367589030823541539685215919123567355378859047481337767801842903040059913533013424987728803712275460328574768439713712722212014626056000338978015444712983691675004456323737275800069165043188957724305077421690313079465441564143643952067740588580376257925222523446184426213861414156317352787277966740136040210135632130854523430636413038275132777642057389641433495930585786287270112445624696064193458025287356080351268479041888471264945309550283954653082034176194215303877969458895249669500111601537050837533747;
R[102]<=2560'd115553334376489796483187516179077580145977358918222934262383407884859609485225263792852240876112240920704280388042523197174281245397166680213252864758774101980053138314881243186871233999346968714510291013416445057975436946686220642867762329159483979478719352815894660506630894530251618572733278343479246746842391291602989608996940577633905578311554873278753380416590414500914368205270062015239714363685819025340442688879785541438098203329878896705418411800777791341626840990597898642910170249919710493781656181324515484033395186375292740088986879627875333699151463459442550282910794854482315746135381585254661797587448837467696291665371677703923152999694673238023197933194145970508504677370772956977900976269400137861327149816565748488230161323197215149194472760526783556;
R[103]<=2560'd142627985882163398186656758819230554505193553130597976292014405741628603189146361726649053336938818653889077460289028236613734069736128282393932313794882913581432694977713523266023117019903757414210492099311678389766379381878741578394747346720723489450393191728056943847287773047377225170807890165207654139316413149015096673876767457504367785126338247716011669929186848894692322839718716775207457746566433104086281646623787906607298396355116719185961432801377588532878423018004790381315134701419109963269610829174930873573477807821309659287937631602701624546120063292549708302073423548912729250181164747637776067540542500899585310571544742576316064722280638708128427871537366137995915159025584694855760738618433370344658537422145018461869863640289196525023115449708332100;
R[104]<=2560'd115546722739980474480329526137868337807856828698470564803914481822959209989099126455590824417461061084271124328819486685696289722649030605633838544944257380633693445765830322164648973159608113501774725188012904249471331866779907772889292009828916059602161886248683782806488690256209589825693346063756855405763294498121717244776347993838976497502896306535540734515980339413384049839674571430454790444831967013022244292985688970213149647194759012103758583892484217204814147034367507273506017774131880767840533402610219908601710751622750204740873558047512531770835298117793014253174812883319349262197704340280627345223047375492350231195221258120382727416391101634070435612951734265140104488586162426890281796150145452654874449402140451547497452414971360175967520410468365107;
R[105]<=2560'd115546722739980474480329526132034813330532845668383172466323087411333054036379020434573307127829556973479434202240916469833906844901959562319486953251423896520576263968828042304015631493693401299381282475468950855878081535503036601357435736529858837930243690116739608096653876161577494833276739809490658611452180281130119400951198522562897853147313263993759619191201307736053102234834586214190395254674696499432576675320914972108809311057074906951835242558436393958819018874827323281416705783727679305580769958771820196592972251354533377274573256857619271176370846271863092359277838957270711452894271603895564137597863778388269593262852046046597257330416079299716120365991497694509469295375569521407423621287491156874358199014899211307018296788996458104594521370925478707;
R[106]<=2560'd115546722740006740349232757680016847769738627611122503933025322306276372413742789929425240083119925240553915601508495477545885420455802972341514810398782503823827536010459404797888559189534530206377469165730855268229950762476514875401729115137043964870486418710940137457963932947039069598427325489494762861737243507239496063841261882085202244116786779090189659880480455025832687869727138084670907765283559793893241499791255699765186123488122744890251264933060167171973873051631242953802979115223106512162596923364324311838717958687845114524513100661961612130046757923143774987084783516159898827840025844033223147441116775311278362977876070681130470582305283125207645788183974033234103172033139298887708540458424238760129960776337524369260246110674553608377959362898117699;
R[107]<=2560'd115546722739980474503818801404957826031202979563998549025184451467707579560696365782925605850506030826066347251824046713250646357839070017150623149715639699314939074456869761125855121191054444771694311591878632090626694802949809147994985635141119154405262911328541875641340039415870146127724086439733761741344344015921609600740568495541137693803706732498063013630977145794333008921925347538563316172855030931363927883901939628677179318893381386711952993298832735140868771363119170363270149310238422614856903511107918362245720667826977581105941691673165592964031367032216859726345736000776911965556422417583085113025606231572980491718901753654788340617200152691896887839690203327922188082107684978312358973519472358093591878602576829080464703869587331916554854339609576515;
R[108]<=2560'd115546722739980474503818777690934605362589700973338545925379247235396649416366876356707467572339371732264572444695429562748785855677053249377146927192772339727168669802815210531545318800654814227760345531220570931810054320498795622182941091176130214633816061005461155340389813793640139447350849543917079482330023808536807892915169788554718133646413600597972297272111791295420708355216570301469083634551048772170230671462254120104346079806021806805540497377170434382333818919542303067165101998476448337012803129136064583855904057582141605185287283943885695823177353904740579630507414355862212773044663408839997191041831707980923141865203743472670844627670996453859801916814269108438244806743752301762140766189821569956422307014050641856126680042747274057182417718713992259;
R[109]<=2560'd115546722739980474481797604354146930079881579160674152826335009961085825269435585371156013299819629550745441151111574592091367994879127497841689070576949143756427359865234249833291129279608277791772353833120322632455784246290983012926954122645945255851106875749883759631918177433369920841621925330688306304293718512187904397017113812880899461725921945379309080807721650405876131038761087893466261886371367480752667322655116042459103438596336928989776097960167162235616172749553058629291759007892705073927958315108772007705076529323513437964301072740584567235404038616637354539190664028931850152902085187229870273576877935141227617346140433605003787369140901232709603272770137674894275207554304595062577097663509449826235263751221462695565175044776615756337018956059722820;
R[110]<=2560'd142627985882165039805023042501880860498663422396791064203303160961961237334925993027784854852020654107635563599517490556537056245470469757695565892295171032528694219830518449703495305710995488047001231376780997525423666159134093932205262270536278019186910200201358296347279876039725731597052355172993434579670316161804333367368469945293128478609437339333566535106330833382189772332767084808178836576813246767250462087791508274707165072267043589991155740002917993666401976712670686975174677454921526802259888555418580784714662560996295888008312831068116843028216121647545468099637297097171459678959142105781396915803084956695645087383555644083304748953246158890474247721477910203264519129798819325898242037314827616752924085939911817125383059953413246664785712980701758532;
R[111]<=2560'd144426351019398421528450960115815473095211824883102038721252844377195040244912767434228808197389984824031856138632205351113601123726760202701809861994276133256926904490761163258235699001389548692706181722390945932993872766122921975633259555243425378820369820214427999317710142284037256501816504090232305156513408599961799718064968211539632834813638332281385554203676732829354061889875513179749519202298207023755019014537032779310663335631412943598024626683663507336631269907825331457405847535943826282072425730245254741772505836147613111483629037516189168960729932866689035976507664709202372928995602616260439744104791883325020203775647284595765132412622291239067606979641425750950542799364664151396830203415187297946204652270745349305792423568390745562662108671460525124;
R[112]<=2560'd115547163408162660961671202962855970685888308194562997654957562857589580848392093389316305235179687079134673333747495553632852951316531057826236725804773602375925958783905513945318245528559119067492323822857844185866119024965962256464156417280436733792474111343116316737697874178979206636567186092896259810998801030123362420465008308925498808831375119471974487797564465471091159783184344197315922595619117775345546311889505842110799274828848056540388393731242110245117751459003089903722354427496090918691645042324997254816661359786750448876346657926017636621284299350399817318837281083001236228266962463684475101661868904650870372512457605802802039258646273654964555574270521511065638111186727718706935512493575353971317030138812885064787436724199763725368913163916166195;
R[113]<=2560'd142627985882583754715213709887980850299487595130662115957630676454773297757872314649669352784309323842652991594838770209083652497251975745928287637886041014388125902339444242980023905800902594914309610952257087252465941041549288325585936804562459051572697467787539569471807292375271805769406398010118437620608961792509179170691828974690080577295085183793539218423087282079112203690106160122067814448460404662986932460295260102220549400221137393882062972213558599205254724575740043381025487542094077699426935799128778994932667967994831213229028568488275056623372339754149682203699646877313487242257870026604068053795452412788352641411433497599526655176318090257409878258591395729579029078176647154132829240508708678432110407424439314792948895195655142335166549113648202803;
R[114]<=2560'd115547163515327508312084770870077767016175722486494715799242805608997934874789241906798501978873595107764903875265879627774712914498118907954710239141742967195759431951433380057746832065597150058606032328167372435065845040905335516669342309267561862875626480528553161986798411524571676152838753920077830561956986810718429409311359276142883394140796454915859846046835073004337923464653858911666914803783495653759882917018731598429852552360543978040164125120563768577057009644655197348323425617349193740415307615856402164309469677176148505504638459045305571809142733493910424537468690521951081184302543778386954006512117590910025467391551030392565464991892716235158543330114712816649616823923907275565920757197677178400039115587735522372991380363426960499581545556608304195;
R[115]<=2560'd115553773437202448079301937109562422021819285224365559214495344754319147242996323967421518810375279384165408128453566129576583905947756148553911122547101545215247032955942976435823211250122552878229604866677636430629226751948282505270209588933112066683776718055439663884621807033409027064434783381094675930863828260914502952030788694331386711229020506039684609437577669222791728183123791776696166477144741060044546078700516088291560344848145603952421018728609615818269354093592305934570917674338622023537163402101473787135291529619670087683375417818332853162904482016468184576731042268069501199500220996781394214607918316373744672741102686907515628305479239862108788470182022218256890700373995790030854074464460033490642635289067182162432067682522597011411046927939421252;
R[116]<=2560'd144432962655934009423799258761913481817087189460724551378169454916430329537415369938127330238956957535350054307954980192057309892802731161955170556762950303702440532470395414545385425733340262308740911675156593772867188976114154799963050812401190843870983142402082506241235852259016627164486972770654369739574108960403215433402435546002207107680901664853480623888706199059773928451645671087857344532323815002005823024782270280262196728459027264314687290174999563258525269289819841557251949922141122025738919376762719433338006853006143854949530934096147259229133317768274103024610381091337490790876309292025904848206599960123847263332398992919826654558155436054372349557922982936118716555467191398902204488077551725795884305706872709317740960438116743624724114758183433028;
R[117]<=2560'd144320566550330171887573788464096764348446084982487975461142231043860008477668209640517901033783224896215823175735024825203746309506762992910959329783208661193628377684840512884834775869080416918001116301121929384235931063936934436709109991102355578204520519196079080944397638275360905565677218296086907733781904676493588815118124105254853979971309494881867286266921872417836019010880714299772647792901488222411242065798534031071188430043624831012435504428583460357469582880594068734362727126981765127564645203358986194189254435475305062857808651865854108132181457726094482149588471224432519747036729983006196227357509404296338235408752058442867331627000001741275959243672448967988776841706953578721080274077837766314879020699339704946165363758759868289827265897694511940;
R[118]<=2560'd115546750389351496842343024257687691038032807933014068924189325874721798118881536711082970256269851292054875374669135099546986132371005441041000846997623547888109046908988222569563185506400188399603945182812414258254050502302435657186962139433121135871317363318433504224395459460138724983879529055825491729686481134347915229964338182940514199403858089786277894105447256104524931565521374229666759489243792659707265031379398973904395011493294980318086117417716762571241574924283416408797787305964737019003876335460725575477206419874172918235277462993890783542840687650374104803224981527001067838173447578058333787357190235821492635148903923204358741060630657520570610259596955244078830016252189938603012728200566973957809277840540065716911372852214436886438656675368158276;
R[119]<=2560'd117352112741032918342650650545995890768122785768016538242282075172831471825469853540029827770640749868314166860716503918947175950551356297247218947690401441502860704171911465527624569589756278717513067807909833894782660849819437527880657349663197549727269335450697026596243233909429977792769896683511201110456885594594651878870253735081794871362729885929251421578120725499623244118291627543686927010041671467628096821195013081485484070946518245905349362749931797975737488226366286932697601513528547527281668719834214845027348705061368502038691188327184886045889946881477567304339625179655753329390984483730447785886277550428422353580269877218526170555340290003297536354081615294124130693873992327260957840850254296699080185451817326186441051504284349069927980166823560259;
R[120]<=2560'd144433403424975593100411907670875793206613286745847207965469888486340017206903177304158802770180597777086439110617160652345325937397807810600879104217621834972237478022690170630635019403501214652729094039533148478815802634131054761653198088880579233998826893722955771921520194097917714942703994155631218714391245493714426849352770897039413246579610823114356742703706851683651345874657585013467569159355055198278645371982859379683738810496742715524507667109200697066232592311672727966113136400641458338646995567474109860019141688418391869535550107733811148204635208560085986903976810969487815518482807044334629641984606211999857372869231576375997067640261694667434119862902914116922016905635991335615980200108612851326100087541224588241608659364331777250261604075600888900;
R[121]<=2560'd144432990298579327328901539793029225692417966800785526481295308750655903962650331855163168258449713116461076791358351573270824964479733829227653119996296989328107861458660424004503723513990404812871768661106928966802404444599628871604619381382509873359245133774336744165712573952013719280852164902150863731761419446575471760007837303221115587484693452386542253974457619661472943937576264501683408107703472185756004188233935858487172822102457831663436200779651847599810285783319932965286706434506931449440372293982484900273150658708170117933580055858516697459558393789822434722865031925625801877430841810549815732245664705565515577142810039951240978311475088412381035390571749719050660601724725106181030691585837308138360659883421914140971627735933598885808966410025845828;
R[122]<=2560'd144432964370988645936159619356819974937219550194858673509712004001447739665203201877991273019824126940310230754353483621907419182223891344657938782537711202570200420316445911806614605580803747208860591330144182729190186020039962032080327277695370134459453769295530637709772144518801768694064712137380895443482830746544043596047122956348329347267582821397297526173727893720468636601392465831889774797653892016332963067508102969162336499771175765834549720860244637878571584106726475116381473564018069376685322941250083180976435776120454677715493699042008138291927223667018011647265236318596259444678487001335949481055620114493845847747826015825333960190412646240780594661114323577597905621850031196078755508638019005786677661848785201448043276155609969186379542469655413828;
R[123]<=2560'd117352140282792669394085057289883430192559164799873108059697277707069248098626386198284940603799589147717747969332831042952857154440066642877873883900315968046193892227581435133936926462506736509442608424109085231690743010902568470275505793689203601051869087983161871525897077118232609952894485696969761777683520957575375091782587748663258673500605409588538888369112965339624506767919382280703594437032759171265083893484803153601768335997354164589545662045147454650799029547216323920290096670210656605924274127722154722685837459125411202856194212097300459059122282568842609683427297102701524830465705319713687608988393188251750390025555920076559699469729464973031243953857514210989057405789280314581229011533344894787564054232628591340167733845041182401631226425652823108;
R[124]<=2560'd144440015162370482357821379137659872103308310178443096184179827050930344109832846411377644850715563513736104363725432091571951481950528198149488562188233061471448518455722062153002724607077362072787374113916186730098438077450534505717875721905391983547903021256267116078812620554305958636410759339919709644178803655979833802873649147083783957542954645907724956647686892486052862104673970734598718710247834679439977544689316803021936317312778977961071582979722979172007698034357510915167111685788643365119840550092616558684601035866667210205084030210545605554682157319442452667578142202907876683221654065268573227692454432947856347704583295083037765651303241070245493369238226247729218823471253615861648636862995583568439563522812864793366628176745780649278434846643077956;
R[125]<=2560'd144433403525861166368205648961246794457169662129145636369355824071333312582072962332293219772761129412143383689544274757387352224000743030621791042762745210895570289547837329567835683965561243584486081727476828853738725423645963983392400008133878148935898197745328262891844338820265100010770853653507733656384413382605820219823537063832066572370246512697848640758769240626068230281527506830678739804518389698403192495717276290596554133211746166268950377909780439216927860236456111447308993778251286019079637830443200029750987780031991697056352182115130310087988469602540712608788000686057322588188062590155625701170307600808864501397007634900273407936685531745764868315393620642027373046362454263933069140051456024015158562532649342401860757740498719385992063710207951940;
R[126]<=2560'd171514666567158619432746897090015394949033252295904903369592862264929260578404221342165231271002741113197575773992929122405448041799060480443137379486015580276953419137778670956043851483129279366830972253431327859961544091838239532708096912420501403382071316625578281436446861468378686312964587458776097283424091712271333171732253831674357724150696835683424225251781106331076078637958398263985161317536590283814344947074736234100231005365304279761630697164013636173664611295339205163285640309183707715558815600119439687315539899273779059337807719516016610367302125518085506057582294886001694819611036765515212506825857762827472073297561008393364731624902676948050279074646940141106919165120926790214605318337967034947853147505235357614336572577027640986191506231320134724;
R[127]<=2560'd144433844099857314380267517075455944653953086777659327679519731529536515784270592549678741747183104720193382297907466899756203714947211108239033326360635634495234154401730217190115620161571912814543191873795532007726360658018887288726832445405555043354865285401603772093272390416080908892087650137102845312146628817657117528112737210544717667455895191450712707647290987756824948298983819221880076014723478587734936660930493872199997139870583157302516290715831512634374313612938899705431127525343091242047332620281284109072673629775238678438522868100682380785854588244369792078076911169072722916026233690542446010537886104224512986510146400399903346121484478923166813745221049545923277679493064352979912223071434797579870382283349917519521298660957991987657309300893959235;
R[128]<=2560'd173313059245760836192514000568621645237377902137489959777603858787953704555580786030255366373236039873552761904031949847124769680795920703237986340241073742596729746878036093207182763619102270655723582540412514370273363633263696003504330198101374882428403801824058938661386545038530800437143177746478239372739508541936152139116602575751371305174383780998475008875325956370843619917713878940172073680824107864733436704001840406076216956596704768241160537422728676880055628772921841564866571182062750947781714100712681784254053444020627513561654949078662062705611028029280826553718668743342875543100345615113999784513108774328964750780155038763227961112112994897355022280393104670994794283933634828105970760295132671261931049941156630909633219222015062062546160588842878020;
R[129]<=2560'd144440455736366636383125507215130285375329975355420905829923206290564959666151378932832396690383499103533859367318477180987375981939103059629437424527305090509231126009181687396351619413105865339407716711999208515820234284539032049617283930648887764873666158021143491173465488386602541108026077674878162624699951634482706335069665904874113907017777148579278102556764967457430548960245948364681649444386447884315542710850477870404188751321036642417525673584755441683472825252976508637238546801502683879856804537909196093243159941064788551124105925555237213105707665778836152105801223589313473430569487220872621423255591521307990987000163272532837588196957725055257653182212934900046882061940195681328026715230795050714651172984190752103689731098289455094770171387199112260;
R[130]<=2560'd173320084109970711720396799628981192934865035181757460987426158999377762725415753269057733753966743606982627063860151752543688009952234547648777942188891156743126990810830316002267676063423292384712090282897995031066728954361463065552404717944690456596853868817529051030173227063852942143099614979886345431520937095536143418920228015925095033769731697677465208663844534782685360763564445136844096822719838966541596116662653377340455138813434278154261582260216094655941595504543640187124930797253718979458550671256830021177176509802509011351023177524555883206660336244627418072161504159720467985600158251555826617913820247836023145321206018690454158809913312783667540743679892487841037728770816157924443627068001616690746235404905010577659248356329260879617983396079486020;
R[131]<=2560'd173320084109970711720494289198074994008153202260196325996383984686929621552508441955920515081812264465494085139967473131977906674132816907423851132346526042865427651591517571432043495695444506344847031033755116208399056781092165396374938082521403502995187687195133901463739816894763325125742643387672956901595406958128283997107512325861457903652394499508431896518238418955842407154572797271302946896547458732931479479562188180640440446027137870021558681091459482310034634408694221805935564877918049787856275742559932373576251611665215065085653664621840114149169937800508438942046689339846760119558564524087656180854584845157398318539131272601717151505126779670370880693440419259191401365367582491856828186135737510802453917393676623775059822652813515368057138072384717892;
R[132]<=2560'd173320084210856278574162545698167181107678864578412910053064726122052634834212296742538362384380440399396159168830900225613286200587859364199966888635088474614252110075556414558500770178398844870624250758796976288384657953765912664137383997137627837944325177812225368645524902528535042942123499953330226027316998622455400716097202403762934353187614945121580316592466746113863345511547025847140033402135466963589653298159988293448786206897583282229588008421238334004890352867775972994515826364595698567410668505184935165932489420554080779223890001889860704659207601923093209339354539349319568968884849619678957545196899663428423175576954679737558681095697227988064407765544498443166283386570248063179624115557611164707972701130695242552991770013871236874949290991190033476;
R[133]<=2560'd175125060984600617528270236199030682600872391078375281485491272839826093838626379473351642696343189420832235796534899981755137158486092679855825505578155810093650166547750066102932448756027423602461812577312684687368799896699903243788676204725283770990190747619868586359166060970595018726652020313582330664791067097820281015094526227867214906555704421664521494817613495847883232542220460445393373924668879194709910755652522819462991981790643895470010359668245640205177777322280183131521867790481363609055442579970237144934465434726026877785564621957671955771620171622764286402692422239356725453528513130353005986065193822503302822080137713789851496363509135946893235708040400333452493029307329110493185456678849769595614950853216985557430125174587976323360481983326340164;
R[134]<=2560'd175125501646475916688205496515813718363103045239186188284837111473773051751615462976974803588759400839522845650604313900865608879355796223582157169363901651953382004474023928015726943208358027840905489906008551728723731010675430563277281936749081635993046535564230472453460877997089489946730777737463013379306013288558647580550396410521764855094826930426560667327931327371678116626567286435772350827244903664510215482723590880850408655229812547546765897074251079501816747583762251443554572113422950333376104435275156377432084207430196949631055160793631677548576892427012380988675140327903129604476121001519301097893427755493402713713798619158523832328191551081083928269961388082332313772595009199524831089025672362818769518594605093290551435569919464503277175909831164996;
R[135]<=2560'd200401348967628628467732716463362203381269480250126773304218003278717400219152949260187768950452622300445165653164173028297777373925584879619204263558944835818646274112751909109620128551783507304069118965804451261723037152233890514538051263442539357575560954997308615248170028991677038830240842461451892753047477766794914789859206178913459160772098794995396658037673203446165641839039647136820794043935318773149969182735448203332442951484278424232704130951716250838162400195151202915400797304851176681083576030853622945326432741384464387128321913121623003198809266496346033726448936672079654461471136036669232242746201876922547758024740258815937898371334835750466689496128203733899606602499934148841965821174528620575268244736264085284612634868178886078135031777647150148;
R[136]<=2560'd200401374800218740820735295750230321733491766827305383932756715930686879948739587004942294816933040229547478833862965257738274929750864440853402684339600441588726133607357560241755629613854758249087267624673065566208840920161771278668707372845699733001720265203127709547612724205147924632306633545192187731451020084330882042284944239494732766606567521779115208533903743662466449079683575062025173707605741115817163741524922716626114019950295959858765557000376683727062452029860847830138472086892068419389233522856680259373065815451972386418592703715571203603701769623970677480664157060928420142333173497652070367919646408310570339961049128637593694896166725811210241531071571535568992899309263337417418751097000325188424944826687203306420093346972224164792954970309936196;
R[137]<=2560'd200514185747693830755262938299350315023706051820550619960365347801903497843993803698964817235690506007116942222623321767775921016185372206256860630520789958912912819920678746408511472084632206274997623235933265084223302447227695472801506286437949930676653810863869030773151756177736468907007244291784598999421005766832597191732827728852277739632209590180774085820214985038048095383576906927034244649516769715693465401331489453503417143263177518831799124766176219845471181145734518638339507595159215754859120874701701025557785037691825609325264907169257207898599835950088082469223912603806244650083244683742724824770648029448605638123699514775534833943364764202334314805454433114256073729419527325900247070914428758983138037504500424471077926321871539509703941229390349380;
R[138]<=2560'd173327136421361755003213623428672576960316163580955603374763197805823053999638242235390528160185084092225507335742207804626926390378668556127359110297022796064359361656617703737138794868679893620086666147172847816712873919479002267768025771599623492832730318995938505331567223022438608933889927319257200283878852279668863272021234349015093871502087508632178445908795565552747224399261272204465971430131443060561277895799565252879796905480551794997922574485589786284426195319193445766446298654640405714742653971137516971480635355265883474554411680173566464445567737896996730230474953328492106162380964180287147586775287585277632003675720670800702075972455902403851139010075628684041130184839996216842977918436844866884647973616124436588218572319993822484750400147589186628;
R[139]<=2560'd200408399664430245586692629395904247967357521980014679215149076614360461753894817144574797788884818028862250024356695769153854422924963947358490739454760106863659586451196687767684693926217939310557361093320806412369541241898765510962074404004868498171406673753005077617310014125162485019839733053363881225165041352751363848836286444428757772206867496901710312689619222393111961197500927113505764017540448714227360033343320197976225691978727232415613027206095545770868485896879902858895440479342215779833600773789789830711983553318170252745687627163528271383844440842820399057410332134951994178096320366167635044348858526437164247809254197277816539453188472547779879957561263867855237646804044953043639586700208467959247642808962322205805563734297833310887123504028992580;
R[140]<=2560'd200407986437148412938024753557508022563329563090833857872293383066573107631720508534235589789434306514966549530130698090826208561959107561339924996903009172048663654082928908866522060951637251101399620597593176112602590199413662126636870887071309514180443291489529562568362723171639625334320244786052769384801578545273241542500847905801213521227376230828117955421615782613083977516530485885019163603861669098168420993369682174309895600480178932106744150786777019123604316614396013122331958060569741314834215381913923835996919381023038288625291848780684310817897543185915057440392243299871844969118461489891443383063638680577366596214618223360825488708930418610006517269991553564840728063953134814627731202357685467724102437137043976145719393458515124187873199617409827908;
R[141]<=2560'd200513772621297564985220673926882606130787714869097518489467990658559594524837042090883479272265846730969959293501114540906331786891367699745359180632746959834660504628099401171465047824038548313480497676526883266487024749508467769130725219292537673731759171171656844109811559929285690808083590844775480558333096203541602481737542620016695625378065140037965524413815532256575886297119918462320384308185798797687508472806178511344338618972080050565585175746522509518882404007712507379657858759827126588636786492700344465863705270788644252802187532713001217631263662200479826846603597055105466070510757824178601813394837819402336749419585810316462801755155466842893825174376476774902972047806573864328459516950746688683796498076318413045716933019611960464893093653969650756;
R[142]<=2560'd200513772614992217056866787319656556323108012397043977953644306317053524025283297912686666436075599250092585863580898595495340477595291267238617733271829939717252738811143937759949743653490183179399444153770788013571744262365499867190568185164352251322932177174997609909990088300750223745902239736121393158580728583062824549373113098288886198742209880143782156788754505220123882923940753925149326791435420178619803288680548499793202899250315677803586178242640582169398398469779500797590454540216001959416844569864815972040876473105263396875853599284484879542583678270123869070479809627100486783527691077173002819343449950926087400254527552384967354861951475798867383656658498657551363379574082621134528105786280087378130618568813670051391926121086716832019485074127078468;
R[143]<=2560'd200401348866742965777924976805630368212816704232532351581111940308100324443607345958213553709102361684172662023645703709531840440380783677550653289315108938864317550773436509514990433933070339882679101426571834910774718973606755705206251785900899705337068732209340673399955265723348322729224035411525843407202048195448154929240869224925213783098151879576936623397760431355417735973655547348421941958926898955701229283169889160009403073871409561980526396499356934363707377680110881888152971215910363403693298484754581525942030684667659981823458424021956560125892477325211714697654780560377262355481095179320691140593188408309640720105179327780294208048788519436185240997552730581681236914743745962582609460083492982444945478593913887821143426516255289902308607868491023428;
R[144]<=2560'd173320084210856381176778921363167702529155344943423763233718197188477904055661905342755545173968698556972540426378951911753253628117869030485938066424601732026816016809050692583113069767688989031506274378937889352913504877010316999588693447751075461550887023284695568445828305665696770246672277150982774430080013564511271723932568931743910093053239393583328470427737702487220991903947274497870504685202227827321988917371627812999226041288539609584902409631172203107405228898935335387770179286074941380580446182880798388430891999826008710239438156340879176592696405802027378463739383777812645216950030659495475745375361706782074706676587861461017237615499377117527512728731650880069215014874144568286642553645319297053606045018889941814852521036527932224723655264414483780;
R[145]<=2560'd173320084109970814346599893922435566018663704719245323402356641894366784551260783104026938733051462171952834227672510434147700452164322940883621700716720271933754137301588502233228893314279912574025947509791369695019825607904712167958147539038573028393723111455281475378552404000928774393953102417151493164337021933672837208145110587118009734258135824643295412363909512561203720164417019431080043954452998894547837911526029068588012740497650913540188836988895686065064844060744821867811710621116686704878082092735470112783170976108992524092166109250250694566149014290246760710570768230252268572746516219302582521501380827295480193054742568940924532634478335280752800008334832050524321857538066742164474922893189509753910762716731779204788960069981672628597346700481545284;
R[146]<=2560'd173320084109970718134625531075792733298815691460631983178726589883017839195417704471215361514408003163031713673989893860950654050558787187183932813080739985397622153175372512693265554405312223991233485752060794713537384851621658286083642461888397925135754578107751476591633022589096212746859477605388788587976885735327151271619197373163304795517745797047382971550059727788504768337325204314569785859630230229961302993771557315749643435218294094381649990566300347362645114545971768545985449969434600018495251504272592753531725568432711204942570912448376407664583280784876410472184215418464201770327835081570053836780249102568838664942590019022590282533296349496167889463546841129255547207985687491885672143203956877243108060789100481382398044702204908294990991552059556932;
R[147]<=2560'd173214296311652490041129546007544938388449306845407150614215942535672371340160117128629715526315991726191476550100993344951558696135326629301181651448180620358020427138703390599775593814766070353975095507963043156998866737630118756881538912309696379314780227781530911939470934537001469984748943778876028832801824046074483651517105514097463270116988536455226513114028282303170394773385518065207654691282210020028168272647581411159950066601401604234774354132361107975537893115807872147585606282769174384306143142955314676154835106725371140791023966927487121843534624554212886983411256896957812175155718648380360042945634121588575802068415847512151334333907026284009336740123847098519247527333297899195608384116607627090268966403290681117097714554489094886130933354319856708;
R[148]<=2560'd173320084109970711722059880878247195429792390127949869287941238382666468414911119108615778059965539475184691547192761922490948515283210802569882700655128218655121432102787055499288065747074105866428903185923952399449619442041345462436761721090373821256015624433175101777080240318403865992325352138917674131507904968298817814668130718142972512301945920318941497052162865673936672011277503693195856239879732439805474069416689571379908132964670411962267010280113167082919602414337149430306901452086737605023350197715813730802823598392120473335168383982939942251539228415547225081973971275422335568579015954174213358510899680287007406237951418021727664693940100373010838385542913949017338263364307059641827668732262167231233399740649333027042451304130160902267050657158808644;
R[149]<=2560'd173320084109970813945808806104553961558041396985446303460286969156580404314533844458724650083954648390112433588120102726603268507039989017357139355735062443893343531625272278834520596440070118851959136391105181100541826556377098031022871060339774393203035815364295571269763851113300529208340154330544976422096475765221949467683204076994093989116949433203358536623735278984703004879833248500907497388558298605708785617497302137125411354737315076722809497175459303143950680821329837075124748468940726597710368961753945705893131959502785486953216209473728803431146240474374299069254400314864909678345184219237480071293968905806743333252454133996639158751339345686121930217570613603913559263106387425397466018387929731768574043146113291197008251110521534402519337704438907972;
R[150]<=2560'd173214270478642027548652531381583748392246053720238493498107370779531661049130598855672651135166585561294342651991855695674277913736894564336145047125214949449108934150023282637709923900490966041139893872965750386032392780297188436965206652149893055757687311599141620845560042392057487317381317143247283044082160311161979541697958883215073898799930061772051248228247204600357500740471722432107015890734688024962913646740658857109041940990610952748735295566031512775181280609754770685641749583047203647564774024963226946810573766908905054037215460083770113298009176609254054703642975786694265376611843593152637337428631642683389157484740764475833749549103450340591785470042372162772033938359539498591030056878774244941114210509030216016280500257069004907621304421794989124;
R[151]<=2560'd173213857251360188910225171821718191344796229765948923970508061133728845494493839774548343672079179986079993762654632804679473166337291453242751109618529718074219608551104973613763961839238913264654163618458162395190604945028680461484561150667077805973965308134854012289021501142331992559494016828087921591872606199497180745229884910696767826933565426500789247274897623791548781079377741414606927028170669467295163969409441941921306610777925589939366221998510955268362306005996367081499658752698290421260105400620078382246553718747762971110869110434835098103322705432234110456249840113152946253724658296518769539285800593722920687114700096513766604897542213119526360257999646824968637150129129867653971444689534594340783430928341937259166034194861227721232612948923663428;
R[152]<=2560'd173207247234906569607712495879843005206999977939594094751079159209325232996594703205596029005727169424953987745136601848311858713915234396677065739781817524673717571743324633948796059131315757360945894201791903144767807344725511558621784029050803965251450793098644348230940253834287504022383903830644736480215559263163552369104617449674875059430301281421851787221547438016804679014384841207425525887461824298273361208247409360614673769195958632073508362953607027769507974747490458171027339440829730458064660763883233055411140907068612214545636613519829142589619511681536797026991788179926503537760923207939712026238591992117667470858576111663691631451393235099007138495202307539481830223830336282338399185658391978657623183408796487937330106819998791542573048313566025028;
R[153]<=2560'd144433403431282577033207474102567045892699993648612780452111854615336952267106437801156732353709236607809358865141213817041379864531916934168891178896256159898208052939991267810752008986857885642063646778434900735633663314103517329428342808920972537560733769776532407790834196280060102573342699078369273566870383114233574452373432498000963737897413762452658687147272320712569482815710693667956816916921946892210164734892198165261940869459755359275673458756613806457660984877767075960724697974613225709201061332714387914470345841551050036862630112135866228757520170512340477209487692900781566017613498350813684262382525068787157810917529663047527462991531871154231050908864821879526223324936158849407394544289137365346332854258888316416860059963252140085226721346575488324;
R[154]<=2560'd144539189615456359342812370397341046218377527512121058613238904464320235322375943098637151481551602761338416560373245420339279184988381820797126528207983596754059569983102094660976868149540598287537085551768786902458032636907828938457600143056783901112180753250884822155050561821425191433897058218971443225072409768275791760548052731689722771343218808821881113133805482520399096134429783722238839481110202797201554889353975275379752217271858643563305417313116198686801495783102773170180482292219452279188693462397661012689210647109324898278205095420711532293990050358209839468441002893787995591603774529207082247370662775164480813982840905515503117217818532732166514562078931623405696663101052645857478673767145911615600994936104588222027788533087995823937242584340321621;
R[155]<=2560'd173313031698114361899135546682356408942311283906184218031978682263461418226310674853195281509253019889519534262096297795775228922681207924010369674700256053996558270413021029930535535577429640566479248414067786104990290294733752478855104389691658521179557364624363996953068648085954800518877377982036383789652189055792980804738046646898396229761941637858803394122809058346115581593631860581289585492621115211767063055576621497325950401598181448368808033063646044494057444113263771682241518545483718895529900102295043046050778730255817569477954761864323568637594661787986076281179414977738349720920386390770625474732150525502425828343349811873206952148341326943035349926572690286113722887600539342561576686890206880640236231166661271471078990328009681529431375209766933845;
R[156]<=2560'd173313033412773374774481449580121819229847374525074461276299045989538362139983133790238018926641115399312774960502459638902286673442662385703304281657952764929385492887203976548060644856089196050831258243451520585649946629942689756190957160661564022007875826471328350901456373395171966539476760364235465889845086992491599699743995524560051236460129878126858068020124407886866952964171291894317163775519438197569084597277713612910270380028992381181198225754565095010388743273422627820619291769725715638143023928795223017380336876291220802509558959632669899304232085238549460517949819100079329821624637184218312115409497512439325986318147110015111015997562777003645374296985037842829890808475516339946885134429622270893208760705828518025582481400835015775388617096243270997;
R[157]<=2560'd173313031697718731851017401598123323291987635240277169199855318346921654680171906267928562333667009149531924536700047755639106435216707043518132990770038319023609042475948952783986409390042758965044075156421233196539572516935646328443051025767993121698398631160818985094826275891084764427797328305106369634375993481551774918437776701409277168967890884673830514717492218297431896158707436123132933790137440872249100250150242426394382310266786863188407238987990326530498504373720259582921688411433667826759641255508275768561732060225915562180443945372163517228127567679901324713892071860664781733595595937886018400549446209020089566906720214317915355370462069175008672938798082665477020576951286202991235473872118479534704002086925299893795303054434380723490654768208368981;
R[158]<=2560'd144433403424975593100411907758039595422653194045011173311101083279919586568225187345136628646023252880863018426035411477691901501098598018069529481014820095735845612135527626248487460854535517217721039747945159246734908255049688382434319420476232852215546048995237740038899230324790781926864424811330006581072744172247429159429841437296925101608418878503488831945774959506596975783591763503019391409176139593557321454024020384072676648049551424212204157861302310623591960893920028539329179111187765523056089796227908349797967092305891915187218796255602148342377310216857979549998037188049128674502235996270368806443783338873811216883000994972706976479557555541504042757270610700608790692126644196659549012940020280244109150124591824814659603678976834783569896195795277141;
R[159]<=2560'd146125982370968044211074895202125743789474515880658610747565074959448935246242687794428600344488073909594642976063119646787933464495565945542002880974922190499465496340087389983318109857682075358259766840099701579637736419970986936066932488171465182193045986180789541500918595081910868869619124354688359035634542822742148918290241672884028333141990868620959894501810338283972883167687030018197142960826650721374505816962848632322709712422266383246127059903723315424767370811024221435458463836071569537471121913364510831043809005761131510899528630581333489760731011444741629050536487099974430897093185932190271968947084400907246865861549765419608157830979655753033026029617509952250047616476556361567654464264458153806992232543066792333460235336356557875831709686639711573;
R[160]<=2560'd173313031798579674850352455345015744002956392879401516759976890537605717820828697766572873424031227252724647526428765112065974818952915310937856017576767796039904582768369642129290118944835001334109112848688727856912320424535386746982192040446453308315540449673028147740108335994030766555341397582553659158147868997026926159623044105600043248868913853904783990081782548188049026837925420236128403326342361473459094522705493712744099952552702349368557069838437760606588875800595050940431968350649966284014448200466889175887875478240574568033102119781651484462760044079107709700506652314570406097047518636616666051055962604246727081455687035918560453193660976838116873142279245595080621927287682558241467958564450998691160633821578893311882811327200899680351179985363752277;
R[161]<=2560'd144546214472915906188216184447917083267697661374914236183806726765012903282706018956612086518966995107303719134065482828282725031352832013298405029756096106349485411232482599908596175618948964444752960326754658288097625936937715653490339693540524228678689558462070802763896790267995523945895340254850406958727910171837706633489454569955303434176397635234992528193960621379848900149440994961188318692318639934318797740209291987550226936397143813078432447810126667174882968672311017424707956492843578775411013528250259407150478744946022344874953822773699751200193921129674081333558236568295261400967509107834554252537698043135513370112051480377877458672904805123516779540718862270575862101205188873912140096676270128997073297149048441947926368577986478938816138341290169685;
R[162]<=2560'd144546214472915906188210449767406108712749415733807029176397498404465893902998279016454565788261122733269004106549394015469230269095197366971443567668501108595903952197662463938391751089441751733156170555749192084733231415116655948829101409494605503709983684189196662364583783636878618359421026894598322513809078505413493515761657061336601809476885471097236706410774928555179726417396792774063123980196393975455443659175426970896141925423108070099172779697944165780620789608322413879039275724577260995736469561543074916633238916647457631279837156838936718932390426446639203443039914407342606550580387009150619984087117844102590958568914739590746075248296794852674982928764831868478841212316778593724887475098932924874991263666782802360345767772194651540448710299009504597;
R[163]<=2560'd144433403425369677347402127601611979397705948792962051861017397849111114359466429641032757431107781046039574320161191557143067248607113169376988305386093989693202814488613243633248476872597978315209679885413676895558820851068004805940651286231397674509681589155188261541145663887477694211455326604031939493135485311334748805986554906424720212900482186635118395493023704359541703848240825016760456781884112654110109778767510312750612643687450527047203246995057622388133973435738779764369829049211565800258187614993048154856774349375926540861460929541205531771807785095480594288181004872215251988184184191555602780890030714630913679868755805011956396829285356438507525860846539493882324703763049415422673367179575108584526147727426709401312521655131196087764084567980725589;
R[164]<=2560'd171514666668464337562858743284225453170555658849799169398219949079883032495388804372092277886627564607958240351674115780730741725531988169153489695176591599802402478901635164087182020495216025592693801029525380817488162877438648659098922864539933351840285113560582187798839460263149891346972398383977406466344237346110397430311777943006282166811215862371112392707469783357164916479329204138732860125680021348519757459216595094109766358096847548980743093646638471227489874943917822476388655722681628235623275528208884800813208142205931978535703825688060924757062700640981716619865484923209572908666849117704071771236109585254094022346778405287626541821250831387636630986432005277846343396856625194584858489893982818815030156379143733650150333778394591909996058694311564629;
R[165]<=2560'd144433816652283697983570140008654153158987182761268512460212590145417612017325149494626871985292369731427016730550613411572617942221599084677548029020710547686349258719957385648518397636579459121727261725088042239587415159226911135944398191702095789838901185137871265435684324565789199738087464612620097947995891763401457293415090057411702772778427237011605341763485897527129790215173698469971973176222342364204809480459635274251562812911860170812164685480005463838801475995220260235232427971442419081650671460268361846501678592247101290402538009761650776902402028438754118073870496564674536480398973016480646708158165738183551593776146782622098312004796986270680427013675347919894898228243421864553973426816411168529657435912506211898285589793066222242981842188114416981;
R[166]<=2560'd144440428288766753741702632134906372114042709993845511007040384941832224154562950338833782783663071687159285604339854903227108300139027985994681930652072149493552890701269694410557360517822047461362693314749294563713513524576113690805468479318090681968809625713111939055128750239557637958879784048472349246840725438916407449885331287413994503893821890776975620299349391184396095695469836833140248766600974789470001406126787889121709365488395852118556715208095338174402793750453038111415747612369272613793148779509571973590182106104015981661802433601030982001650990256337083551398296968598562067523039423808163053734709801769462665912244287508660510683696321392813643429743863466035925065208129536452733683417625296744198724341445755102919529472691286106250112892449150293;
R[167]<=2560'd171515079794440349431917764818048133813697858416410792227615998636538846533899964659388560943859315356599964642081383188820108219977907345645881670169119903725773426490642976874107609155687036583462177356584767979502772363779388887524088024134226473187406691021516564582959565586608071715672519142733374433187843661727362072354985717765338162632654929693145389785649389425828590021202775831615131521062537323647897051869748174320984872823885731292685434345262384967375671025649726688152322670777454088331340690455479461883441034157325267659657931422513427456636068376339619879164821122216498849294790301106731181316272758777193938589183026099021073885959111337122158809908517821218068035146733463883171545810229673265502745757805506582637743734166662192126006303550428501;
R[168]<=2560'd146125982472247592685725616208086933110427240655618720147005366433949296225878942786743362448820075159665004009042066722909108591202641530017955391604595554629199691787929450743240415895265260234194793678104904484695959213416971936597950650683198629966879929250644499485404630565550869198906720330441288938331450002680116184478107779023840707473436530259825951493487050617842978070181313993770054807568521005992795763988077958218824653860051790870433647961030406939224701148198159711235860530316286276757563556623608257172035631846738088812890990763479299492439793882515566621183565370367788502567422259815216046005748103890565351673532837410369711981859243820712175810407196423895920198795149235161356024328711617713641413902420040021088490787896581190522365732088796484;
R[169]<=2560'd146232207609498125042037488862240454357760646990620652309270047383938709815642496771909542570575061543384691497706809424012309320223521682936240719828602433042205123965554570866202874051887106061184992032625229928245030403551235159576267554440120463230479300201231434971175643928415053949771110506136777199867315267623523608744815377699974098763560872201282752044169904354044987566043951448822963656568942840950978787841087967438976435558693957855509550706650711199914381761036410850304499816360039455930347477820190450692600299079598733257433784102497786823943549927395377847479957232792726359727926908506462968721336143970318375063293695472020637226168182924256213396879608592788321271520933698983027270507980017713070387645434576368678076264115415056088013359946224981;
R[170]<=2560'd144440428288766747728448522090027874021298136381128323939839399165382982315156219310310248927835195444329085511914178382806721415902712330469609974777285359147594895410320192342279918048345772311554721404942581009403974369809778152906826618565567067363740582580151048332433415162527232370421148975680408834897067318077633818379865650324577623375529444349927736140354061159001131266874159059413965223830873261961321677504970369217083510378053380643602912938837844165009501349161814445221395954533331125195363108626896603122384626942231682280083241324522231598390170785638040157104242105487004573770731002187236911052733547032248990440533976544812358610124495324928519009656751670962152183983460705121965492095466879154089553051848627559200193267586868476726706888064193877;
R[171]<=2560'd171515079800771867017201235478850071306248088221851286530788370807348448931987451848768641625154246661138144240485220747069912367324358912980900039243862276776784251278180189311889717778352614866199212647682143815134964017217583846502572737799176746152845122917827693948554393365218164844217150033801872478674669931397596449307386828212993498522279408714422341426170833465899900184703979414099684927446183359057494767469031015060695908752993158015267079871563347261681259960748162417429723987195687449386295399959519949414553514443561092808370972867316081391601725123284453562074408243752753805066312382561725727125930537315501251492622312733185381749794275941062564155558204838967924951770017397569941791338900943527250581932180759594239517358107876851903410989266457941;
R[172]<=2560'd171408880490226449199963026848659629679832341481993226099798801334938391680489620867737639959337982464787988686013060157841066211740882905428752205716912568589145210722299429621319635994128749111132152352670984469451829878623469037181543526705162374081193655093108650472308921599622612160959618428891049614634568343465734197098447751461590565290875795958463251272715115401783615158968521639732689895093715048297377788542071502078144786925750387952911972202641464670528084914584493974573975204638918115218055737964714624339226647491869779252308113313974094997222375731766155584548763712696904674622331297494966722764763676786541459990815561454161525314216775645051177480854948000783390048438799377894507417256385531374052922081367185149273700760232754431459731002239571268;
R[173]<=2560'd144433842579848107118332476368203441277481655266914415011360878649905144345951942799600684414707031128162322050403171081732655950882199741220656813095316865485763614510098700707564465880866341444552943999663290615004875136818362156025091805424774187782043208371474283382772809565100846852147114363124356572827822953647066834196247161635677536312332769978156576284484760551485931086120560484758402089411960346781671278039322012112417993395907910907678936785073414963096662031653243520261064676107129751545517361092699067858059457467614950270990005384965217534239611137973583916663773381053100155984310635707420678764410643341902727973397694801524216004650021000341648386183150049723704348808033372919786123900296356313543233005861076566691500450565461458189747337911686485;
R[174]<=2560'd146126421425348973372137693965814976745246505703256733426587419629217607338838258094809677575320983737987443286785934439581132037885518644815349674861906300129067236930302570410978307041665429312087438092482891515111543036624151870286070969862084676597561321644380336503350946524862174844359435231006645173492428084568513182391767617267636750824426140375899795824364331827251943990534642317093105222940004829027058888551495938399515170395628737698587113562283419586323088509363365982881664303204766991485176968612510620424951543629620194801417483098682639355117675685683498726619921480602879302663524469804584791258912018333479403847922738472298760593012100132485552296037071551788128940437619653636459412732889618336593081914157343945036634682748584740436913977583555925;
R[175]<=2560'd146231768561816532195215865223917002871826787930079209976062517995603291734377909320259610942822183987080034852429714141147170380383733267624660306228590314077297775413103962554315785198504177021309085508932003642948928344741417789981082126272264819270864050984872639494174826795226745392627045034950846260895307899815557049670368584140874069803722428943838700152528108971626310385988908839686803772295861541630297155411349640150122909501694558471266305543443960939787930128620509920345973287921329809604874505026643789906341213293914220375901968964941389864438945270108183234425637149221147606670377551033473223933275444100745300911651977908027082199483662518593631256157966481425123609494957094561047955958945243727058058340262662308781610570662813636215767698259662165;
R[176]<=2560'd144433405045450016700707033793565872396068793531616241346843684971733325307708074528770536662152971022363911794890850501935839505317449392751151118911742032698709272615679664317811985666573114681442189202633958913011886481575410824877920644998949103594767930217896226110928552268222415263273985819659948251070969065203134684918446926654972535081311578990807429617830622354036078106690923539550663098149484249429575588556256079960341870984515029864043271157516563772284994417646743790939665262153349309415654036281449398281949159923672552822040204135776997500691068133452879661166879345284680721295126303141358958068123369110620266135957277159757641937983373654560269682881017231863919917613181457169556438536518477590764964858639878377251897838103587955589121950608610373;
R[177]<=2560'd146125982377667380149488024564184584819922123072713163388101920628479957696382566711525467954726784393573788662415433291349903421840170395775338294053007692840677682654161315706713232112712834867424365669459094419580828482364025398422015978590144832658472774316492604929439075881354911716756201902911573409619692276710565009459738724236944210155214909089897232504503822526761499325209852483023935688509632625887984742842529858108933284631698249451747499653515265306873953178741386862728451150218739719192286523208818559790274811664040352085009248185029237154605910598033590622555051036335009758292425993070214882720821990216397235852121933636410221447714974912677157287950412197308562335526734392482734361760349819074948206743917943234862893085597397724097719194491376981;
R[178]<=2560'd173207245519850303880864343222191164668249746769240691338609948596228974501723249485853012113766969841076170270918061912041119914971084650978473700639037840358621053408372986434431368515506546303464482617031174262651603905806464341361611889981998716550199798254292015909271615384500866190862854800219477044914735912151614123021686769363944313151548096162647925538531812891307946593222017580536435332604742966579717814963288400357606614657229207490208206203701548988659092695439380442665273505907409852299413121198412964887410905172344632906999096644152156924942521699562303742023639629142932425893669599438209564515860028412126229900753836084679701421419093047426841636371097972859488848641668470249350504384730178797847216134295008992697200053880362745091094559518446933;
R[179]<=2560'd146126009913542133412048335301570305688323283698599916723338460615483885970148754233787057868486525380776504791298705723401218589902616103423086408394712218580686265279167462523777585370059276153178779874804988648652004739308051672917291590493347007461973511504731482903283454690872188101268177015501003603766135664302441105303106990224978165614782253300628155032045367168209338891982278160673374044344649596359674222677123646487928606546843977407284254345424657157326673146326718237860136133194630700879738026811565622861753228428203116996847576968247487946771000742018523439320420637781163739305545095586702672945636407063292361590278120236787871084331605708745202239687478257651025445703936329136626823164714400949238279592069769937349596362599568487292982848415679828;
R[180]<=2560'd144539630277701118497641091889174195954556622639243223635203991644831604716889961411955356687799885090883177863153357273632907967369113925470161494559630772216734204280645124692443513076553587830740752463667703841735998865832360962843038307468009860682888354393071971921467227717792020156001000735627411400085275514676478551020946735082488277416811363713845163716045549547988620582493751038697433915256914137633219367951982765703489320867765698117296807451088618744597999525355604638888545433390635489591109531047551684392371761468107697048438813334468397981631772641783459333217690325444884439304242466267334949000159663901163155998407479590305558791034520550936044634455302047239377537884218132348019481886609622809251793030549296453469586971332381274818365983053661525;
R[181]<=2560'd146238819246427803573446314478527505815181386211839304478886387738239865294643415080430412823799068335750800090102798109370240980523878111841365726357830095827953811541836261025638862155729072455648257425227278466305721369790477121015435820757173255155664375799521032125958926181479226927906041994397319282214822913253725569102024318163218768052247856476776403589657252077292288158087139626117269688440899959340043066897615301134400126875706216617667076947617767878056709510718894527003133714434001173462676906561445234188455928429135714031893740295656258199884520106791049640303207095446783120642052189035616037629465814471869638124261576616500671051189823162021505695965558604882093242950864939967908341773901133056338011131004082561638112128327625349708051270121903445;
R[182]<=2560'd144539217056724633800816733542831520082140599106411597678389114764591980554187172877656579903042914204319140747224267794776391478056229363822411357234659409290617814749727141968410905873696069216439042268793706164385562645819856308229577422946267721962942541008112238202303665381856824675217238241244809239316102681778017099801170702236119891366514899293347965144348922866106285298537276693534839853845155737528973406468371675766804325632056162698394636594432249289210742191641601413798230519176755738906195692503924931725126416724925284837563848489344362848028763590093794582498567726964441466772948137812282868843443134969045759740375756495734627029066586435898866881050971351622906826644677745311497095594307447287168809547168779624563042929108738068211786824887391300;
R[183]<=2560'd144433430973434782739853940050741776409004291208131793685619248817035350682958668546378141739796133524704857530909216945534931302659980697579837368463027634094528753101376496498421547472985909711380232049343171090267349789626883038902175637961709430198123327955358686170817403171709172435073530166377771033941267288876546126533473678494450256410441728513230244489253720364054884272766726463609060356742761290801925808561300063691626233660128467012160949559086943486543733302519803145570263779863063082453642338539168450554581105716570374035263773198194266902886346617091355286034193710460589760258597702129303100264310383100660015287859330735007847283801648527583165551887636558300090838753733436763820300490063263868290925934881439808282619294049328282023534014311519573;
R[184]<=2560'd144440428396378019015538744223857988127819829238411557027050780662998798293129690354306592017353065045010263282782594907718657232227350162187249611477650112598507211358538212226910289832111840997970680647318844563459805279963726271953142678257993950956786026659147098608667626947926220505063255017980250534259188002217760734948171226771933829917231784051566523048496247758313237561111532228872491010198328020954868552155496879713276508649673431918623956695574555476676968870625589004233906183663657078702233117858056123525963829263289122727834935189259323673861636674755572244392403236080417600542861616454884308364751381540996090443404779015937141201991740969195433954769584601037633828416975066256932829436235256242560115683504116145286825783886599938472137152206820693;
R[185]<=2560'd173320084109970711720494289198052122658515372603599642397637122773103141315620273432717243000144364019416400419618651223682556650883976464891746915247814524438646406020850361443954626222233086648376274847634417262639087498702508604992251451692423207296086971297530777340933661917043296398402193589008793277524752280407942280544505974194472900260482465284865781834148929429524479092932303019003349127568467838036174719864961552569899367787301514832176302681621471476224513842407376491767288926705437480951875645162043103187381255611132678083738221722595507353091668762524172757118170445140843436621049142186970520043597320708326400934755688614275525796524381863259888599088074161878165643403258887873967717484625999905631672795018023778223771763466692385812246474748417365;
R[186]<=2560'd173320084210856278574162545698144476659215983222750045244517858658223608634412594065705119391095953715537752061982471990827293916943276766978303014578323032402756400960304131087651002602389190991327330748116561746771216470609092070859598756482544691607908449131350366642487949933413723462722713683586222255412219265655139923659577952058013626889368779755695217789116677540282423011282354881423332016228329416039091412366129281564257185989699741590248281695287288679794114053233741849413210914829483972670494950023417461707323799876570602477616630963253068325498278851385874095414203030873771267485769660044011022565111107455262647891106725778629145772270239067656854349653739275607888543216773918390107935168164666300866638036725315233643958833720848059354537726630516053;
R[187]<=2560'd173320084210856278574162545697802668603473104194141576818797060828323519467341683979446571103357221299366829679977120362883560459545678717228310529993296221384673508952908330315156407903759902125721189245556657714128723227964884673571674262067918844123926925384359559945960405580730493848602143366806161494449517721841442061571521876416892410320255256237268784923178866937687736687752134768223964963133566072620045038194001722682403059766559476570050336582612745657756401969624981093716194144982595813598585756604917549161844851130171224245646700886372933020204698142375886945859060582395147098466974573839166908482217172641535910311827238994763037282231109480309163341100405999483297353629143116726772078306406658484303616752332256947305023065505062496647396800857462101;
R[188]<=2560'd173320084109970711720494289198052211650740769724901421685276251209038702342021925711395615016367082689950447673075385167280463643363111337012144158677146554699106612921750959259439230256088782095332729157391196905391257217807526622010709004588437296856857648171036523929692625785163057793868924578968517754970497990476174901885537259659305997942301617817261360358765232153192088594144676486067665103959594007136819177069430365352150310168168468980087149816202636372026358739343620276161744017679756946429957860959601136856386622415623877370564394624441436167429441908355887630288329980292013874866954832151580154352005146893799436485722771287281206755968278119688447847057046646316869382945713836211426791826419583361569888888478384059673754568418575752256987875457193301;
R[189]<=2560'd173320084109970711720494289198052211650740769724901421685276251209038702342021925711395615229026274340695297616382874058181544847273141146399452999920904365780999589056834644103884031514913375675976706381858999415059431906745875352628055033550305827676820688765416448889182272756215651910047251384328858633700394298108604739527752080484084903738718767205240592657930631886447366157580453594021415459423561755979176092936397289115177880305290217896150743027233839486954487452535275610813724464893988372012585461094969532723707144795896980108515074669060630998820688330346216532642367416247530739224916775078018446774072065359347197848635287677059025061776952193594718917707543593842310675676890661062696025874476837946843623476893090034698425021991874989787244364387669333;
R[190]<=2560'd173320524778126728543438681601089974555781345407454668744764204579998851484515655427933211469975501703259390263991567365084185945194273589957944376105138953954551706345634624431754152784111813277340589292299649453857766944042503157274718316710324260434430362043507849944081164519005822278207191498360466725905655046863301400032114721075223049271862843332205175147706575000050576009800942779249080761999769980234956278853676302417019911746878234538225439741807450577418820198454316325909089583523331857850845742994032266835743824061462698548003596649104347428373994576698285196699850981885054948254212874249651542871309367807695134907783578205538402210323895472216511092437716515747090189355249532164742813403138574958977332290672578216709084192881274747708850540280894805;
R[191]<=2560'd202199712281803653351994636397410003041686187264606973412797670864415967354259390041722998015697982118751680571256872140523573580233809908554606201832801812493427306734977520211844769251312482141824428936150955057582714009618253585845399365946914557888927495747554547383167260987337145497835628320604111358809564463310197983184007717048375808706364382837965324140197430778247059429205960078424985612688933514346092789324295067990434964590709515862589995736793641333943542423631813185606770512745874227200961785221438197333458925185456704081236118199300446816908465736871054448134519390769089172002390723974123641763541390022396432659881100599580330636686763542831935164713138270633561157065534239525371747198943599389472769182766156119548938845972725878575049383859279189;
R[192]<=2560'd202206324019198548596129204947117961654958725193827525886045919089470149186524003168970028367220667099761071851373270516466266998956841590430636641394501706626054533720889232109143420218102369197417127383681806267688013994437535042070019005420515400021271325759078024146934300336588350980096011699210098908546120105363063493513970137430226901524907090179815472561060744184988920112613053072268299288068650629552176901520292222827764687317838202266908329126341433628443510774328919524129704117989498933610281746417148332705477550035183556838037670266402233785830938014202416810016184540859815516683117332135065179128684931041532133352853564232110759737819892849465043888548293480010066172346880664776616749053767567464530168594609413949682501458921481235554086656390026309;
R[193]<=2560'd202206324019618898712022633942683804659179326937720548802019962733131372335114447527774197702305198972056617537734045765523109575841488552945818949289213609446124777930120612707055094950998667173052421757786641353691045857945519094280876190467846812939292185814190901967668846474487474554061468544926431625474758792426114943575903224133042110812648209114272722827189180381491509198930004363679706959928838683521719734767695221682154275432827054089902752270713737805800399220887294100799716066667721939803148757637298825109656813561273050614140592782881377711566912051278275579596140633548055085158867542229969159223436980375301169275227452885853838495608625889328791722163773592112277808047634880990721604720176679347459808717962935244198072008488739326430831658520630341;
R[194]<=2560'd200513746687007355205154146199977222683523948934375648381457558878148929343579751310998162874256400066981800789206283716580870357292668888944215526438733580333877794767937065270858123916367561480823192923616103924803084695113826985815295200982524755944500242342859314474986208551110625258060656808234688149963171246656068870513994376781182227755926486437070903915188789379148406268581210647808044299234564705130117110552140702014692278175921090391098624766402067063180813207233042996122544886414162934896273884282193815897015625022246040690653123650051408359624376663841683870255801082914901491743209425412958612469766675810605518934658776645913468293129923255042833709152723042398706685496523544039515477477943291183360153931760887188861384084853172008096442283506095173;
R[195]<=2560'd200513745072836740141635330736485021009477044527586253481070727969096995972172747917705737497162173397451845931195766532943262759903850999958790286134310497162347444905803915130664297535805000009189559578997346235336949374689955325885158969269135059040115226757255538726970099565512459937041381077403805950996991284209767608819880807939932557041452482819098687133863075226197786710240716960145919552705816761494318101628754110070449743642711684107592258844388661126820948275428006778200642957312215038212860557976296554441397798412579253788953014667181159029029345297960579844120715959031739805754900673636049471265403601721406982330047765674080896643930220613991195673132278701206180900066356628894424922552637461612920592543781162858952419062100174190933586217618723909;
R[196]<=2560'd200507133443028491929460579737938379130514333516995792728971986586778193367437087988753531183332204614620189336186891257068376760836661672048606335885043402119263768624071456723396663003738875128911587157180049530804294185765036571082835445831561558518732238709828089620565737801842280171586116684696325380991114860147609468212312007231522803218258880547875830643039888809484276333338115470788815062453026696328890622586352443988347634535279738224145821827958136730820627120126501449929886103128457382236267134670224994868852730594472224510921708585577608343773439571986677093345456360180459018669245306439747150132812563689943836082512710224807164148250586691155630161671799625686015962097790784724620376011379190604549599845802788866173458454353667163917984181182092357;
R[197]<=2560'd200513746693682253325665539934772887470333125319503828706026769696382692038672876101620391017743783129820488560079412378865822332748877874572229318936554713917303834792353583673395569895757050331577291412415098445688695635199238399270297959146713270132791186416790015873981021086851942377941874651547867380374807032011954840658943710630705013441427280809157227133951932158120089672412072398436227900894023097810195947839986265107613257751048608104823176089319843640552180854906938902900371432292895413723777780592863839557878822858778920163915568749669685106829150634482042812430799546075855902514725422824751625112654253321631288295831679656790066377006500823636238088528593801501427727610761611276809451709343189449479729696025317477222825899631728321170630875383419973;
R[198]<=2560'd202206351567289913469973394295239698174002001025897663857751342825274035278939060692284661951104096048452780342696197352183273173279059299321200793684146494077650555204786277394096374475722991394418361174377492468876893311768430134269860932290644063263864538054720449199433315316954698697801448908749723300550482101198748459291560492250755430873833671533130914100873554170121635399564530642335407045380302291689244203636368936927769558351041385930088098153667043956654295357360175408410721813167300664783761323121378726536799939080749488485426776958227818795261421830909553729927569317378149326876081750696702460173378469966277604929620138047974120266666148677974061894357028784251559144006750201536170061249900087711454312911823242203983534961020505174625111918813467972;
R[199]<=2560'd202206766409134900024323593984155077787398956223044937586523579378548076017441057629198146392722328158775493619911786936521159324583830722292327237275100344354223541764202920333753417506084737203281401276749054048523756556643558788467992369214308581875467289311046381292573273709699892791959884971796387183630485126306725216677596166910600082398218215511403385329529752221988453447773743567470043419435708147802698127474451003937501471347915229794940199396925064580300334550317178248085805518461171732248751336255941981666899753090639436006414953853972615135816369996450741256200706516592848274120456366753026104983838088060233126941805036825752209318888008700320803478373772866025606256503384043269068409112466703116574527757460929553242033856992523093237005936875623748;
R[200]<=2560'd202206766516719899451185915369384928085192955236374426104461190825603111457906252481680962573043139834343031118754856348171904419877820835648530357755086411815401668734489373727667452234845133751127224093092302721356876861959981820557955379217468977707632178017249952316442859261780119307019513008949217634579085638354834018495491523709880093786726374431184923621843173417799507965359491983242022866959720379067633723840511697778564399279967367972260643434048643269694473320333318763378191885096167185908487012751359654940102425132104633828634294883160853667396670775321080443136510022676857377326385856286495307117998030954291099004112181031380401398838037236870926168749897895616409578850169677017742426714152154667540691136314072655880513540220141538525340479371171156;
R[201]<=2560'd202206792343451285848921912356234226584986966910278940954443196802088781347327527615445456809617784341029367759907246260198780251338552441241176432092996549575688574191462916800594922833645224158012657657228166657033456667972596520800544603864405739405659892904940910375633832095227325177837797091457382260320765194621607778787155866745947322248552914486496674302521451257890840006273718078164207664217172300961731091496194250893501865037281545234084095635055634121326924230613288759233746516529385026630451395687605127768628064853555489081718646322801523880538526401298520347002170010961533471741273508561158089938497795161136924579850675050230995280530688547658961852101038642059751887499633207021666078651408800400055931488136461273700987001238385841366774381351880021;
R[202]<=2560'd202319603391417858767423717034479807361179269733937683751095823233507567241319699192973619204283765188629988545831419555714381916427970465888412316477806599720530974058890065756378230697864441002803797107833692735088999507986511888257119461575192074452377630818342520357239802474285801601259663001982112038484876577162664436110990413865847674812726490952056721384461846709570570973696175385652540105783425517812248313005350017315197694773329220280734410499818756711992976721073299809342478680744662156295093090526802684899658258484707408014899254652793100620784210054690102128327872123053872877690694905983168283497718472941308160231611533436756984572441244586581374932297677562055337561719535968622271652574962300459581074600341690305677877567326869724177499741694018645;
R[203]<=2560'd231093445480381203263993623621058979413425993388921870127831551738451259445594999804530123829691738687236964154332414322542438004518761865947288654448907492078731933079052217202600406810549136494010882833635165703182048063470919635556418051891640694508187581747609018891859027582276383783738673322596256567538222407346924391714254175467072885734684171652300133080376821977238409876387643708926138917717129106867726510173506423030546003049340138253598227964427809493508058750167264725910379139257173497821751058016573198903775370290278738933829428249295812098986013990371771151064406251452772440251562346952541398948572958551647788538919144499308139447429189188163507132770530041000857395545912271697025102085104456723202476464063118552606503809854347313588732233728218452;
R[204]<=2560'd231093445486685017814012193975899437600000830032229463762776901697425085144510391107474997392217010810952093779618601723346231566603429843521174326371251919858544664978056800025877897426363253023935338608417593916342371875392167481931458394638463340622099143904166485738268004605917568662911020393596008003864510608757743540691095056040917675312240118432768729643274119001309871741043753689148304907973502032597048660560339482853840478179459261473460382401185134131015725791139420401340895592666190387173415937317974761043610223319274359249413433807966339583014523137687953984269846426119473589582353066596072826443763220978780457677794168948292469553354987362522739218506320232115482040118630199374092764421233509127939594122337739604851365081569519811912247343693780309;
R[205]<=2560'd231093445486686653417570269276571480757192408376715153781166454000783438632986432318031193862789542269290164811071951724778772391116826738657837387514077695714632844604711265552829541280694487177255886690626805379867614605835239219709001952703459024749909854228017107275495272716917869674283367063362178420722511758771290676803661339474230997432431595367389372552710198778940755085322109960472216073611891434176580889783174226436781658230810465305826812939533838371281786240331452714842387127479358038352830698891189065059234486644346816720359055142059479198927676235214235428917464716993440962193970171861615298434639480817608034916975242261848481305749817808760695095407382190936573182478206769796843422869840177639726062653626961011912617140747355888349750994308257109;
R[206]<=2560'd231093447201741290305758653320445569939656741782839921620271365218409893227912346060334196738116389164500411640439184091006487581803059789740089478161466591771276377178028820096541302973204098599178786906364556018330502949117375831623232096836930486258714428826363030747477419229703497941929068776376473745423488848685402208628608679330065460543666470230733383045662225194102504775446922370130437783750994395821871902210690604887239493551875327790840221674252590751205271168621837697181172271539910883690380465393624016549075893154464490845375521812903667031693664596465063672883100916944772931439878975950751433056799378514244495751825597601568649618446930793157980150285226949612167578353051246038477485173904216632835184931154652196315339381503271111906479905151731029;
R[207]<=2560'd232898863022773144275199554247230590730503418352840988261825908378662432628237852946159413953120733378576291860877665010101019140907646676481296205818963101098204715019308656124003663530934036914220499007131459611276712815560359714756901375466787312680644452152961474367486455027516652241348898137180121691647089936199509817461023501703827351942386468494280752308269136041681849393167827107057979293795650313242562105099958238072537556392827008928510405349063038302264953678276693605162197754852740697338676320625422432191746868152981617236818123142363262204512216584549055089935768958565715365500448779477566220962435767654578787217378246375948736687809122602538157736712993470619378299307899490497689076575260285368581405276132362441223645228039933168292046092602004821;
R[208]<=2560'd259980126164956073971285910745319102858448164638239103743228011280356530852328700893664526856863315756677312570636786532780712504789148259307691276202814873997333701713021422996342863272162984962097988644846685646627386082152453067441837808121547378996757579450088973799508339849299395277783259359770085661775185482669715390140207869620458025933396162855251302485956184227096494423030048724803437079866673731696476751601023756261352962745897179676285919460904512766126755799591906059280906124677760924203195938031818685992334137958224787942821068409691266533831098516458308517809758598195523985310351483815250699421208243588009556736750601130013194214610104894557291850836297297435883065512767653592184699318616455255929909859612555612244254710443524302214843054381421909;
R[209]<=2560'd259980126164956067580741433797442918623563490787608399311008499870524785041137364878357473688936247053395408151968988989517889745979888136221371125897005172966288515940071934459576879097124891645019876079988264983043510889390860650400819752361127686704285741158478292292649631889271471830286492701581612548522021618813810198281404777991927921700870766615009660350577410642606773877943158360222236312300558586431287535512949920180635187953157388194793746508040883548979021618479719854089235606767522363545950312448978388081658255434267969760592473756949727157941480457372549613824745292473538259711781080341257599260862354344527277206753514005218887769018020833023467924016938339939791884711957230761278064959771271682435817851277695277014266470346939673688932556905731413;
R[210]<=2560'd259980126164956067580741814709045406016154843366523150713370052786860623909174897876281192176313342822908885306682336734262150941605961375304936591048108136019085937124686083266542687299888476663669102049843250843947859513112142477894246181428053715008771808408518660788716632386971292345877923701816958985534204105201327456881369827352236887587702283346530449915959022075378331699333739754752689643696322914610694812414649833004169803315832539072405024279792458033590157084621488770698211489335083875865318039608154839726104211285186726552490485484547179311114762524595851495816198690086323424476619878060038531339428547094123010909789010913204704035779520512435491945290367073355024561931740551903767450733613255529705103285668370232615590584928565239994350115216512341;
R[211]<=2560'd259980126164956067580741816103644878145956876960715041826243503432032175870694615538801825896705655102456217522980311475153206117430809467571139495401913890471530914339005246294744509261031856581234189950326926538420834287762515289177263221319435931676775473323566053232852396521714625967660819608160612913735463507838926117380871032453369500669876340907962139902881632259753224188532333516578875592367805830098716179537320236457535521273031070055406851128479968413919654831822767430196825227320688367707614726155014382032846596192194323695413437726605094931751206134019442326002705344835875497211348259219840031946263576925886244282893180541865978031376118466398936168455464115153461364255166751697806180492207024980730069098472492474752404299188817102754770769247819093;
R[212]<=2560'd259980126164956067604231067569569953397814060995491342011491160634224165084929923498678617974315052803978389820088964391307393229647295583424863463458128403079774820468606354392805178952717087165612371147980023979041654350425057971320900800170443122096743796054104685896900707677580122292812034742355159409018474488080698551284382148974547451621703249846252559565582427126049238954361364315133095291253209471704620522903174895605520141518491457649070957524611830929566321648844180093400564919201548258331786103758960976239701270116196216859330629293223621372359523405627929336227509012196261175316693690762665602984694098299389263377207261716232404183240473717726911161137283229917150231505866523200334021531967582676230495452386863913711162661813160991737179426852787541;
R[213]<=2560'd259980126164956067605698764973030098907314819011931001549072235361553803553833933244320640053151070090153917049522186591279188389892456615155667819092764207159179744594504622801667963870049709125620765362610568978993641531300440060704326800132014460277008487239217524217817530807289362338731506121791499567133109213941016870893951966573056931182211592628043930272789617581156654979336345551885524528155854268017401427077601392808589986486758914832918029567414589145557980297477918219731824310731845551870087654894428331307584519357957686420231465349331912864484512067027746885002691658054975327988877442351735317224866154641157443174672527642791841955654144248883138457668505789595594595460362217648870899691491922976666194656911639066685405801272096214870393190468707669;
R[214]<=2560'd259980126164955971368767429461309409077509466238789482946040296617717096008836424607579646979845865145343637015420384701174124411348331318392602433930369979188830895705590897952576676152618403197516775531492168954563134517997505052260401833965780820552543108573334715101117797263124078288976341920343584130065882167604024575492086822520602804518918920687299000338672227580839513280485597959157715565884644256348457679581545161886069590850155593926211905817679596048547387569862722875067950275731001479136140084752764058202181208243097313781252029249987951978229030425462557779545921706280265459126987768195146426111482729732772125276080288538531534727851178679819836367518121936495982422411791579615035292881030894610423144702940320690760196248251615293756171836430116454;
R[215]<=2560'd259980126164955971368773522559376525753434106105885465491424310522576070777690773967130273182672031049193662828488745265391280577870004555602801259157582532141237543895082964368889354747939188902604378733531212621005851105622573311843126047835285050852804799293794673499962118546509112488085046215535631435338166329544611576293130700419843642610408438307368294255337171958524341466619955412547292537821246300062995810607707463592280769161044200979707631132286102658085044350523082893343758170665183631687864252350753708476376391232171454029444250650125988427516869261987549443109505152575448300625448351588488960513463887096302213538539530472076150732248949127857864025969836344108298108246680310306215318209380377661891179595750374568317563452281317621793920137298339430;
R[216]<=2560'd259980126064070500327756284688296770443344765322255129896105215054077674446191986686434620803479214174811695819629113735079331175021438294768789313385701105536876021923954775322013385553980190261968164190404239662375285635644576319937761133196517968019542501089995257578629120044345991500159027012530884518413742622508561372889151046005753997120171787601750000244393008027912371380910086159498078655428649074517441309299493225778630478125031858736420924257948199345424458845169004557873501158334410821025076187573954077477867267992990691630265108878292109658436970079249345295973004198651573345138407083034431304908368441974036128119082983543936302495849130387653823953835891020161349590502388277929290281005382316147680026745829153158805648638790107452314373059693078118;
R[217]<=2560'd259980126164954431977183359996010877629421192244503329367372769764495806793162874606640499665065540474996085301961269426528065807620462978259196017914633807608546851118066112326600664798051300528833466263834599887572518117837387420032705600748461883822599604576809824218862243654548410942892422094778120903438423830532968157530915332819088622281438456538703956559416342855390223114036361349783879830938707681018474347897672177957002770347238935022813616681375245233934111447551911444225015545434770565002861921191401124335009039003211657414083312506049953527276084856173942318336397347374187848753932626387616462209596910532090375160615601772751053880195719654605526124743103640148595053006436104893004830394437953816911938830714430946905241054502586442810571469145527910;
R[218]<=2560'd260092964653770558452277774085750361431981691712236324700303810517494254196782366071859605259460739428365630057657772353657958753781511040553434627983647360372117274085621673367568406425030194296329018820293586616800862201872144488643497396808743121105066501508195995843937950353107280038550025895234030487994558241957856111462235429444636232612295508047469120145117678392949692441262487086142872092217142152345137589394585207782008201841564913529068767162797745945154761219130440230210673726564257171991092572468079465474728624920041361685054475656214045571581984256473784736134636615254211194551087460673284777978576549075856055205056878815477232828937639571916301355688370795983560341038702279275522618271314047342959678826556815352798235939753697446964928773005596246;
R[219]<=2560'd260092964760961473234392051505637168737056096965666500508934836268148935080672109974453136808369539213208988856366750408840732455753149342860490459305603026366604092153781270547308642109485615587577546609936689641036530673890881012999059129048210467216658085650006450843004825776578823948601779877651627722800265382622666507625438365234695449986127311254800262965192365087703829488807455922784721113190033479444116387824568838759818283352514158816570475595350042169372815745562999732822296550944878778013161759066440117049038690788902977922877979359150352323794924066431151490810034970738182971861739417576862513895777062884371037817268003808167807615585290028076069354857065420155885937073152403798318526194090131982356306865572381211137549728111270261572938922652489318;
R[220]<=2560'd288866806849951179811747416691804456111910891650210135222093941230013275430551075512040015027203316166889263745587429425862643610805056537274627360868283353248653102949154551608227993555987617114776977991638448842998626293354707238653871503284226902478435243539672903819457541539478522636882263761267500857251570457113190539796905848515743401515786301586907818752044785806040087061463504454170373849304659467424768102578455015596077864905977811548657173768743939869773435709445382621092004834399046484794780696043898099513186818689361893899067531520939793833965531355680582736989639441626291211950162361876241658181062395997719324473418862178152773849306226305178328095704794603507098002783788458893065006309086523733120721146402277639153556166873226234190000537247110502;
R[221]<=2560'd288866806849951186601609168560771520060194280524098096799299245751029776485362657104980773109842804323327502384825478792929119565744880778380060413023758057255008226607358271468892211564652477917475595758117213884792267785211847039885542496991055010042742697895121699254910786296136188213015963176130302883200761228612117900066221948855110602282623001514085454669436750361889071702860645658032129283923311477213703553783348371486082642509608564352192357962477008479705174344331553747132366603065339710935884131110819999245635683738556101819391720568918520249847899679683764285909107532757406208771794359359965897335263778701343113974219546499379001467809781342523037181201518069994676500701077510411884869634585822398701367361582935379375047756538356224584948918406042726;
R[222]<=2560'd288866806850345276860477198834781031691906707329246309259926668851178926335078966978000488631266765346253362653625733012222317850303541257672467204809011647705244129897571899624639556183562614815883219734292093863115539867913358174084152186545592821825084168019701430271118071600524624883189868989676058708644693076305308967644497145406595353646473119622025056367558246984614765409875188986721544606741333561916300130619345980596194861844856390357717452096022738340268333443560769552990713089617779270396245065971148580162783076290148831893330647441003172111863662817013543078100081903364068172332110657384654678914769442955275540066596947149744817170713506206296233977220085277077964266977318337262356323534064279197914864131796159226999013070327950479510488116624778326;
R[223]<=2560'd288866806850371548742629165476820992702587250880306442388068874052765453673619125515665958028427245181610143568505238536686391302359750906056337479631264508178347526656193499009964868239709803861560440693954919367017069056259283468087830608376349490592351372069567455305668290820402452945530084981774944308344367006208000208169906533576280779750662421708957320261611105305502480032366795544453203398776201610377403618830277132832605318375695221846973374193707769563624573567283977124102165533549379400699511707748970729353421997035594331581253824609453008219485765281006813790585589982498958481091982421764251406715879288215268417832382744361544560368680440116270474279985633017263167275466035505871890025094576281225985015374992654904566805038514067593738856525708227654;
R[224]<=2560'd288972593034520694775108629645955495889552051402080402061686394862356776562470063143253449167647901699458387384739900315611858247558314868538078722657212732160062564345104717418468474622266228593624662814947625209103336475338416909821021290985720562655380353081006436987198478173394231321178226176725773453519171359070107494122763113608763356595007230840293116522952390418317799955881158715364208730554696515336084934460332352249446343512468242758522915364939850190286561945958138676024275149064067760807829100637608147507050297838059103401744763432078485243216320767397242279612974044886479646249520267866740162944313270329049878351699338930764644896411836846234418456246680504856232224717354459522467015938071025364575678101980342569109809138558440903916168944928777511;
R[225]<=2560'd288866808571731527170095775243697348347479237754081687937993293280355524437938833138344238181879482641664365100050855828402115787135161435137230177253404716688368595367804727904898945838050769406667359075854528654198418697894123393291213699916853854958577453025160335544098116814604121485875657590333539150101447973399023975031603448630813498593399265221824055567007243490986722118436310074489657233368949880853022875344970212543455829736855269594307596007912999099903319646218498692609582641575029328791511227133572034819067444270004328802398805842808597377012503889949998906943822507026391782424099368002673701299981057168600783664367216967561651660572202122579593196689237179293157520376171385863303399868920668700777778294215877440109348064301087619247556768552015158;
R[226]<=2560'd317753461708241190682715757857929077792345210412485280142085232511938858113995079814748700851396477184445065885646317285275665206236621139928606289603745014436265581735255689383707325019340021025288083384129161239968896232728235119992076014633698922053399515294515993609515865915747875983005198472846596181811953529169001368198574672847671142827941537139296490832700353921402223713079352174335991623578988369074673285233738205628383525865588593982226805833746052957688234736197190187800229468400085971887179732821622648784962920942095904714513462212025573864267502345225874769307636705756996018869022888243685673479585943873791752841324188522739456689445926301933674128368923004565752814146588145019546101759182462033012437628218819748517606317006083878601434190535021876;
R[227]<=2560'd317753460094073762640830104428110437918814671191536033763068920764073510811271834649190867405410742973198387209777476264817598161610480729341899937345401536993621605276006289492648309794453613997106353699045008402342909593407683583067425754999321787414198242363244344541923241602058660585653467169272569003812685531098193644875076590433243872607455100958186040625538491868252174403629552556298911580098932232068356514545874128538981518521129373411407703083334821348706761816693942508027313344500505572761035544557045372175323312246814407841777081055767049952742469748764764761333484890008254086300365048412561488244625737091565951770236561406512275152953717732843591702841856053049588561517281949537343671303511072846233671602750956487833249323191057907152926467271644211;
R[228]<=2560'd317753485920803507445248902303416291608277572438086903782679358997949219473597823054048260535017432959417566769871018129864825108146614402582845626766841424045038507293247499070365118040169997139020850926327939299100022805044504062251485014452540618167778501428229925769623309842993915880125780696442787039102097163270416756034335620498399107196972351671628532770700856221300498860970239785690038002761339180361854541756842752828840339556063837440499229058191249423732880415873108112600173497444335715598448924767199102411600288337723334963005212827152800200791432317499130513672727295744688822014451183255065134428475226710031010508785759591943248035280054587645089523241361195098197032179479175636090000310887995620357858263366816336804785755250244550367538553640408116;
R[229]<=2560'd317760512398763731731977620729875566385882813267827127800869075824629602041568097705392795870452587379712346385105496464807320475974054211770590832137918922101662009914601694522276524368004702350004591898508001115290547974075574841709931007178000110806724869618867704651663951859549046996277294566269232037898888921946152228200507734520372687419590849791872076734552369478385796921260922435317503731889817044456382969642150774420859684379559689906760071324095369114024811058242379487874749273540946369725456409872307560000312927827107456159767959438863373275480394332242852008234512239098152505641041143277290222158563143905910500938020310749329901992593884593117788212266147891552088935566959778749138506065517071355227841016269597409512378421674818139507454278852105013;
R[230]<=2560'd317866326023787067975471229507657514056754706338078265587332643916376162997662236499336137929133595803314363541186493976207549592176863977963190959197098235580381014477577621617176920476074723797191919221359681094801250503164529476746583780416812838733533037436672603782897915864846470136974527444117725938706827521882514194464684027888752888464540300491764728898716691553481228445241123979947217841138590836424592817160452466721181577217685584255169755381789712632829698992349147758693304239404547204848899729855904484360613987352875142953442411362520275620964913696605042167345034710169252930068821680841337069133840212129350878470423186445721464645482808861199325827000453650622438409660557716300726942693738570767292910376994111822459751339072315514947366616955245620;
R[231]<=2560'd346640168219941423440988578401573441185677891353718414498080865611905406380636536481637617189009231841741977411133015367221425895156304635619182023321294562637043669680759209978464337098926956626999795712215428828167338954315955933909437895204994081424234401887111997329238149758784285770926145409544037258562911679829804700638097611862095441099458119993524589534487360636226130679761660743754292538190740136552503557342071617190795019456197270238568378928328444883980957107480173963775500325158058196391917365201321355157511711947574161390990643213096903331079263555572399016988920377305348012874374459881454112282369984072928654279369330723949769785189579952893478468163265083436150696125816475493747902248432633702998751314456638574392707447839374631787194658233607475;
R[232]<=2560'd346640168213636075512634312370317673931216494215503767680437561378859213983180955464045677203510228796939888441075445805794911053064076979210403796873104767911403411369908830534641595512731596310010120123547061817592294097220652806238556786640931325440663481316171181998336115682528183749304564848789650887727461541454542893336417596848332604350826870745034692644164974433911901949258172322500674218476564081791009525458905488759924918918593015245547287733786260348937605526963443656030489274128412299145770012158718909619696018581614500749253645764666215600872261340387642609188907804755912458421588889168146233994155178238974164532666234922148485349645904400791606821268435638703516751134355996932431257082506883222572889382513828137704710305405549002889646237305766691;
R[233]<=2560'd346640168219941423440988578401937953016199007389836268946267811580470554049938471859124309452907060889721301550656373323235022696392883544152659542516462690006060005898914736444592788379881482729021028080701829148763430476405175151246493154817150119769762244752301771563471069756380790362340784553214971661897130268165881832482283932933252527079830435507599887003008173366149049360540615918875990379376122564782206735259189951988025706090003957689611518263879983910870228369057168741531602085422613663192057101967977748588791076492177664709492002872213879564694436071521484720492164057532912601207819569571278959526566523415747112740764961831915368647286271163882498844679575486455191494404058127344396709801211770261524779020300738445898254624590980364228738262664255011;
R[234]<=2560'd346640168219941423440988578396127121882330137895166597395202979872110245050396659630518815617755026457006939835584069480493345207298704569277835815499910533442415138333137449552089878307507384189931987473347250509694640040991757603803327723395309019745177302692205150249949720473347859772471440644417535705400739136220121272286404767258130380439972887398174305225975068564247247892446886672447728886891104446624514890572173647426611827798894856493450530194701029170482292193850274110516675863864081445969648512322309910852178451082854122974644393908532691968190346229980513353679099842568500261592697464172501883267217568136738365906524584364074209471177360982317273000632388880214196513265138061598778379634284891526636433677131661697201452793269248920546999639523612979;
R[235]<=2560'd375414010308510779878961263126249810023043473222563632376277465812406393227934640416558362353085354780297539891240582719099080239180227344758327575341581286457632923469561611471706263574232923937689621864429163056814215836856630090076462973561840865153389880550660679530192550722235788911904888277988152190478699078040925751167259022279407749544042229153969327483280711197881875166195359647782900075379744978319863384897549887871351893826402277947884003358122305797535430976144643478325547820149572933309998172706206185174499928028294881707734854668347297209794270999506043136331059548776306649482026146714777751755916328722454283041344480254025094417336971702495407328652120630895088139081661434822165743675736505893926937574106501613767779403789763204065706497767905138;
R[236]<=2560'd346752979267881730114753033573771727013600836142968452719872259537860866669920231268764186648718907173091916032667176997217903813809589531799853860593145785372152384965171769829448106801681667896762274578730264012702940992372507925827314503207811043106155882763186411270683263636868931148644894929061118563710158335297111007162414828915403710328319006593151136968938907958072871020551033215438963826771476117755376706166864044408987540529975733183368968977642006401688214754619278239325135573631597126480090996016761913904208871498217208096943361230282395113210187619207790703132530572071500078284181077494739484797108510277717612484684130687393525175300590184361007752808147546805251707364723492535512445323620658142740234949077141100848129390747434655747885881414202243;
R[237]<=2560'd346752979267881736128001408850955581531484518720145318135658992372941514221398280997532052675476112220368474164723028240279658363697508544289384397690010260456353557771093499217486923814886482899099706000262718478882735792474759699681864840570292662855108920068952026950612790409731817636116274507548751322570993348837747157335266640676284072354053503501595039714557012239253269068051826152037210748222387720251174752947427642546441254246256464774740705153012565000210630309635234192935563377668192256266156401811410151964279870086118405173042826525039443187617790854534167037733914974019827908995465138211020852983859040257985324039402165376652594424871289308934182067462464167603020609511670824740602745120158149141587662838940054977729235000695685506749097438946350165;
R[238]<=2560'd346752979267881832339975413279699128866447205061029218773492225417117279689890679187763740326349500839323429788781214499368524300878386789659059002703924859691903322371999282129924105288102156819670871733326782952021120646337030686399130881816255110127220118072727759624565405948040214968520133488003868240302858425703558411612459027995512958505041467778494296056826116784682993099681081715981833231742947816957594618230154843727265593518838509545863227480037201434183443466203423058350356370880583124139251873186321192289724643024485656679988340749139195105582291084025559221969203144403388202371498823215305155700887836452093698785317292421373399005031010896810171455066390437394477070231994659969161428867415189767175497314924472125815496772430475080608497350951073333;
R[239]<=2560'd375526847183156297303773386756646517462077648882823798936402796929333504685096086611402442103545740025517529657294045910742877449674815286225510067995295685365271526936685739240918788500735468673703217310404066979512545494532240897920761917688920730212310835344370728052140902955851624680845659231844007848567702783109448519369181201082596149217669981121941422754927725289011694406196036420685385534048552319291590040055155592559565096177323095709747330027486440226326604628052163188706916573863079330057181757327594674053043160601916974022250024128758158359597088370829754079494944514210162407437985194245746702912283384434842260252608887877425635912592595352495036208206308580583109761459320757350618731805445042359952497987089606873966699837373049746309539590441248067;
R[240]<=2560'd375414012023591682260224832774341432186093865197398010940320241942362720154153961071935164833015641799541224985852731732429230911508687423077578251346881531034246359682208834407349408037865208405918173452377876448770064821394244962280501396365815375635687343343623737480358904048614727626737197096760116982439180324745796194409678730479313828286351880557855928476782161305357850972092347397041322595176417451452513901498929410614115783261055507607300786167271855648315358942085611510019656252972054019314920785928182806596973937684895917996797343109545177790245310315631945686183866341392599730455047000569002688667888469464748521148626439641488100220909542356887677661478832580647360044240181662088774571371473106406511172515988965889393897680821032911031325335647123301;
R[241]<=2560'd346640168327552592125462447271820826084773664378969846900844018080690669578394092945230041385578174169046201159586290676886551662658405419876056804979329405702440277444505891753482453000858821703842749495293245223080057521517685740424040761660015529428806807302058742924890391888359409814973059775733221887552150534045109221942978367736661677105225692966893696889986826782954381519261578132044158281893198059487283816001353585112469349349538776330570811233190633354334483718851052468962565563785511483866557108485320845254106388959447744467907521510622982111916904412978056648126796570529194373372978644249526835046044236947848761957594681743522729955925130844661481869568310852657933299078955993005997116812385578842241376526266395979015602226781898833569397353203718740;
R[242]<=2560'd346640168219941423440988578396104423301481540664168691521215530596532020320214926219256465504328123603277944993230241713827878014945816548538784772281203823008043340230355727922373748805171240271668878609145185129932532395609721553022300238814971960564679953466726135250832556613410515306744993891261978506951962239067605697661912867556342953553374938130734993786189468702873871815878768843425409621277733886857993397145328975810679952671763320195035950846007788349589188768982706267383307287990957130747610789382527601964618726349283264040762558814541005213849532079065579997703016303104140540545969322772083357833123020630902854911843843005892534375101167554306414507831103130093736370523788867819523405170131135796598508433482935271221936059406069539252101235402426710;
R[243]<=2560'd346640168219941423440988578396104423301481540740066556427449932931459321772011086682641403584071797330892669641883462085971192065260581406729869610551400716000463374945030304202391679881295816859551836664587354645135917971169901786736359708515092725250546028190817885553122566332115079741038386556453605262680486692097171004212428169589184212085038596758648222098033725196683094219079912971534376210725440168407031023881892996420870962409422906782467271186876768602622762785098344341085800664489040468491009442933372509279966240123066358087266500973374437426349942578362485871119206254324548050979953724019315947390538667360619566311426843819516911800739326334171382749577363823605403028088678740143054305192539950494576324350595462905114472873649337094989193213265655940;
R[244]<=2560'd346640168219941423440988578396104423301481539450099329056255358987018578857490501569753145881389538556823091392520756378598703362771203259048271938728907303361736039775599115424191606342345606260906801800653495800398467544714822363626343292677333271592288281379394204244566673821124270096571295241872063346207429129335743477395227629981672921642507750889869214776791718136942452759132200126416995955874565094280815503506425391712014604621508923732379226675227330252539409315248948537554222990771843939905259662920082863421083273609940366241217617522488887887540377908680591338215015498275953272610769438116140529853923686687763134059212023134448121571767176764172817728936993018346506910513062265406745632107803915252614103040533318796115206776420884010821662780923651430;
R[245]<=2560'd346640168219941423440988578396104423301481539450099329056255358991134014596825157887729950814840567191644553315481216764193635297293123177008761788330874507837511867348893734752859508526272974934544324407182116288839244844953223952011112299904206950660720857721317647779210306172770061492989086710527630760115125256852305868088599229289115457181608958853803330039208357475753149266487835078467746245912710533971629260823491208862367924706229349191061936369138921882032365175712960991305005753517205245632537499419072440980545818829063865337129752380977332620389037137282977330369901397677883197680031399236759846604571347609788851471174504648422530598435444038818380311980845182126984110037504056955840752868030989953771315012583662916625443710949360334223696976035726484;
R[246]<=2560'd346640168219941423440988578396104423301481539449802853021465380857286487650759585381960538616461536993778354108326053582830020695411279391354892743376928182121733169304164684145811969930785707329934532596925435500717735756284989395227554901626687571347057018973536335274985975446451186579738960490139171962817033845062096971095884402770898534598920577790373796751311797024990604716119118703339738899935516738149696791771844233130632750977144234982972164743579651776919616375432483589425957172719238219371063911418094967442000008583984846000687926549481953100871827430958612355598810956423000359937864370815240723219905685712957799968877711263951862807281429772588896707666512681014705196678032001409862197114292493943059719577725081893271450636608141294311714510731707271;
R[247]<=2560'd346640168219941423442548411501263510328487993179637824042434717669281223299693561269272373840162765092198665858539017124411282378308309600923934403297949077132998236916744908790519520833649470798322793075128151205710986185645114388608153922905874804250656040509929111008138475615707326093160542805901839428870177988140413475216918656803489845739762408829594818447614899794659847968450307411584169815163997569175980954774996827749297616708726694002762463221116263765987974104467495217794488998133054367462590381614488621082393260561784988648377487165971372020197099314097551516790761707893761025978909926536126733991690938029676739228681994540245964458906580566553245599827000284310722205169134384897348673383730893435952141280540128241241227521334430921393644306859140695;
R[248]<=2560'd346640168219941423816914449837511424493740794250367041995311433540574669379976050846637124737482801859805459060756792853555551204919278376715844022157024355508600600035415670149795419435383541576324152690860612624505255494501714010713915272221421576224024253511881988662597281592854658177985043837346852097249582380628548491155087884404580307479730233065584105050210448318382574061137596894221733378704446684616859433066916828255584369609623611355957869591579358597193580284436978358739601996487106669149345015433981014240457586451761892494960274560540061385566208385804499257942397557620703479004442260687929765254158229813213737834330793688590755198812500408834123034523488887140719236273395906551155552975298050356053971047395680551017725949718664474089842967433463384;
R[249]<=2560'd346640168219941423440988578396104423301481540744810172984089583077666636050469505723613701656642900787330967995585649928751640191056635342423168778031306540625089472260971810688563478533969047228680125817763231132322263518207713822077805562587441663777915422731486852853146967264561757173931595859084692202643957112894176464108834436900730473837761983499128684647481617107423073353886022286795168782318514851009682140238318103071834782163223288618785375759651513511786818627038045536930631371271256726007266249295869546858820753716842403375531783941599462872490319046333280892271952640276798872931671644970598473780663221849966141392541338759920838490692409370040646329331375528568438770005097148814539215395580426439717046226593354414466921835281566700958089593205974372;
R[250]<=2560'd317866326131372067003015893665959036601651860453773820427181990580597103168479708809591252460959792899450647022352480106934496344586445573979910728184975708004766906887654418499385757449478570231847337172390413813660959312875614541313811671587009149686819045210006618574526166517375515000114994153659888260795659117783855648883744355925594129739580635784245275891923675381903747265734203373228574132081370798749133138721175544910240311079122646402235943763350028607787175481551887923163558424374274786135100425529708114724117792472704553778950265515096769161298503243984277989551355792328565167091713011294640923562987012115357672427906755868329885690001519594716809072602770663560426390230403527671888696489041894887957320849177634735460230101816662409929488268714792324;
R[251]<=2560'd317753928310713592954430062866231906184860623517346588897287348537535536440914349190523847233279096277183259356242109249073790272779382659694526592491131195400723399521442498702458067228278218056755434271344232027773931501690098403664978130903152780840288242113186711826334962581860110272769137601590013791285605419486612824766678038963608902264228710861671961787491859432886624016917716029402988548026296637624289836821431004839499962327952895858049804058742722706031170188976284062120680806952701227331040442224439255292494962846309984295219320625661959483257283935041454195465232522549626210018962537424045065260507924418754852730294865858117494170506177828506246883176417141944848091532377715884618146108668121088720536892074693637637108916085750244692378261035103017;
R[252]<=2560'd317753928310713592954430062866231906184855649398974233554798150025926295222090958630954009424383911618501074202085463163259531510988125115545518276667966119024895609992638763689429635520988842017079502891361843179649883972404175177170418527358936384252446907254807746436633785953051836137622748526967826502922116800690290301404245081872838309149457517728091045972394892505217442809659997103345038647902031068102533274760353727975321318238265381744714134656521880564651408327733629107280122309477987618293906019011852302822380642919018697275260617645810520542787516375795756003457551223231327033315846061186113381469886758744836280957151564950240719974524942452725814233994672059938047126225359009056498753298318481606484561052732803001536071760848522957877495719411290933;
R[253]<=2560'd346640168219941423440988578396446236897591804476423072381459814943617731880785219567729902852851297666906412983414223674875956366531466564388402286067323730830457101613036638499421089399912468449519092639417597816451786750947870374558491033789687847456652031368860595090151799924516586387643164752653043483700253098216852089083734787440222260990608482582544859366084956160361017877615661476428671907292693528339371065065350714343987916879070921901970187195960366076691867597457396953589014281939255673533418726046211800829126164065329284284080934498773581119846982400717484136198913921411639027848222668052554535796108187029276766033407910425042215575341268691324886299179383230679663325222625255260720205213646496989383849053405821942040783735807293069263054871790327587;
R[254]<=2560'd346640168219941423440988578396104423301481539450099406263555797928604699085286685704155700183589463125443053799153322378797192554154423873363176294533308924109919565820666660490291489171502366077644978386332783662099048354769975383360286771000443511880431429263450511703027601284176831867197189718594785064788462608899094862091020870085353803578190242402317493420585889826532770931210368655729148934818785398875580520007253529838437975729197750443660618919150691282768572632580417586426151510071930683066943810540202700410416169372516173880450967306976329100083089241141453493760306847801637629920295757698111835369892334423794192937941231440095280891161529444733586500421709157199167834701740786364920259922358152881309899717669437768255557809525865663297408472270911572;
R[255]<=2560'd346640168119055856587320321896012152751365916607385772363691906503165932558255657593098072827561894805854769877973028264784505679840867025868497603920948253313631554116307334556192029329430152167700189592589369377879519736764341896177265585603977793525686678197913440086458778297084729974950749548471404303581467517097981555051722461303484242565959677118189631088800880084473024526957006213855488505570988943760135033845316549712060945863306523053489820372954468645052967497794337048001334423649132706798558945259949182444188690219834913464074151612519621857188954137698952500833308194398357458013167805090190645959561545590964839819194223831840061426939657600183981473776837300398542700302124625728390689115097789085227954247104919214113977686066687078928206229177570613;
R[256]<=2560'd319558905077758499734661345708908765231053294180287005130336638806846699821861687082859233781557305103315102975390802456067302611928537268778892050096585108684502255712305283503701507980342454362877601604714406773583421284263420220462824668067888499182649998612598625682620354414650651335605978913832224805451392992444103161974203141044778677661304552031020259452925633370411533367356450071726530979896246040513538997046847907632282846758900214733233590390275226706092534419896112191745167385978891157149596111723565045324479752893113525508108161851891558005125724480518023438851272445240747721048274435489173308654842500573460781770160476055677211361784863474418254246910781400444767596623524015050681301510998344064973574498504213411635863290582468226544466098569626195;
R[257]<=2560'd344834752398909569496505007151866130152092952942419983009574410394754862076591650713762946498655616471001756310864625577437103596013672230327700391901177496148444344947452554669933720019807752394050897296164834535832778862324892580784089488709053160083832129597516194538820318694146979807756042390097057464237415914211164420053444710946408438406467834762406734353008168971566729655404247621958646395694857970934217021971324626633101966331713039429818845950476959378852538032796377206787999845208001402972193835440673360699112590834974781513747550162783183657014164431312312691041397653584781341925959714413044460785113828817542467128736368608647556091590625836213651133461822326553156770539692958805900445656793676466283441778829740750093027744267999904398261273620787605;
R[258]<=2560'd346527331345296002627467734115542137695067288429925384942415688143313311164988261005874703863726665507281898541677338931008558265212530831439626710991673494520544808182507976493038577835743885483559650818140715973933873087538471276117260024327304569658693151953971029258882512786664211782439828201323532582214689552954392001164939315775254585790758464868554262623449817064234518404678373700674118095987095677130544565054642094631687310914694599259296033777477338381854642028942308206027515561828572154776715130875616169554079066038677482022095521444667022462790004872352799905555560203853245140207005123906407746780615940647694454392150275065056714359167158857636805701791896667648015813904375457874072037630405075672300131361284046861419372129039999341347959456631444259;
R[259]<=2560'd346639754992659590815809954018164250374242902493492066808991471967671609634816252704171384903121282769294268400385981088695138508622740234549717508487202569712794995349737797216897115252946002587178663525085458495919055931779792887320350706960886472469357557054457250565324128636786865263217091181637074704363883585131124816580814444580758470493247852625595835464420331470199360098882625163380040813066669102060279791831707795644997951422429637655327754857453576497276014680884560643819534394404664575657326793729288425330552329164237972909596712769459656129441610069562015072577160725859841802266529558095412767013551575771843575355161481752301009903646220811707132153856050489627274026527313326121780548181194669343935469268051147041051990212946303169908667685750202931;
R[260]<=2560'd346640168219941423440988578396468935456713452570953954374605331905678270040827841887686882805640261629055024316367123695012413901429867103507181483117186262712989058236037905425742481426553020372911639356188938600226845142865566690050800967240112514660669470918729945410790499817413537623241274882923091640535132957305379994359501949865607202979700119007270157474511503196088712725526686140353522445207348818950457825865195399282231283864545248607720830516300174179545859206332098937522350237382556380337594974905708352006894488267862905497326318467838482320233713991822305542846665582451298495648592716482748515382511758455349803731611200485416922599522224921564506091903163452662894187862827051234319560844155892431273562463216690964200356244300403455112227661369582354;
R[261]<=2560'd346640168219941525666210958102395002469637075059692229665610677603992878884479689264433871317288100800609409227400098169915240241945251583963998287606754324699441618742948380799998992012687556718825811032408979869046038569316185988505552094686904897759399519762211594454374614547470583573622629091719667421162933867801016384918921896027648937044694018037088809545483639020155070557745629568430462702052639150743654244648115517090239142289539574567767507809580978820941332938310875041362257210095942737780517022813762098951747949443200482374719693828854361416774630656632751375418631436616515861219180119859265493483339297626678785477921353796867014076815494936207211141190090927446792953295577855618991221594272840490037146439802521001445543909926906619651799674547381300;
R[262]<=2560'd346640168219941526042038981556833117873379239206184651105860292714730485270951161360754554777264516196773895614426308072460336810988995026797778461211508975947765576279917422673893601814298396719001333370438442490281568767448974825856902070072421065750172397640296778423154945519056963198360492191277470061054486174002430694906308252023247828674323333948617075311885472368171293441204265708184639369035607602933136883034497898792385735245339171146735671622779658462289783294811402032988408499437241139227717680949553225639549352540676380264880915740508076205472417250845440447078295878782936824075475263664786341386860612964210023633853197402004598676921158610310328298503414431542508035482457531514997563273990464401274871091607591915483689735632773632370582487013120838;
R[263]<=2560'd375519796492659931924689103878956955612449801074922459583807820680529429944065937547164371518790184775380914054370421262248059151490795606485150968366594585975344916122759695389410013611633961543057518962209404908495740981385895881159423471859940915249027175420390450896173020443414919670363849215956925161504530104308738987789450974885736189641960691372357128918100966606742236840033063543254521834593349313210996471279771882357356932463262451030768909193551902355126717097710251936931546740734173903045255950555498315492453560918869391968167425501614667741250151353100671465368273109194187499229206188585097096246287367021174413814027918726328662339483966471721925237504823274250207314710270442632675076217385310898904464441729325894306676842715495752866697181994256453;
R[264]<=2560'd346640168219941423440988578396469024470665468516135067705844012299696505762024921820213269354270056462395364231976543028095455260452211640910563704682439370937070337990551218780008943061288792276132708653222795563859161402852199316986751573259768854171922382688571835718750073249094294234115956944947837451695952537130786342492888952835910763455987228063862062113397145988846739697943215300976697228934044319652006765663066070493113828956296910529646867339775856097260739890108289860138494924311189876143123667370671243376914154555318810868925225101081367919123548228457656894576833380518366768516316835127034588763760690821379869659759462542579874911220789863567532414012921581170540546628279938886159758203244822796354602053938608139467286591613826570265123009207040359;
R[265]<=2560'd346640168219941423441086067965541467409853352444396337399752057404929482015340881470650229423754210114080212966469346530464279422347782588341819614535274894403426242816735944380758864370089342081589791651581018026874132367380616466111821286159425939109964753503871816416316501015097523718650393258997404784014210727659506103293249540170587020377278976579251379294510655969807018227797312043562388873280978675412106453095254665599354709825445710035080870844996289021128183134570740481837138177944152753536987636497677627610857389519708612697014993564196880717614687076435403989791780812961435093261964071194242499209651278837162448106766952396608169325360714874380117115708039447101981714268120956177265505340843094466518359298231916982777067718725853933787996220241237354;
R[266]<=2560'd346640168226640855616430936152042013991380831774920154475346350080875365168619692892029723151421497078485303936227836728583275720325975516689755591942993410380756555900912210105982597721594211298341622931841671621447561003202012662744375410682781715640834923492402341385225409524010824677242745485434968366410665445588436727953110007650508149017080357087270509969114599829527198608125416075042688289370756323284629654176805889016906370153688182317997161619702431685070343724967198003579887491563744402884223895344143490196411178962832329974496683939028132637227038548603539070385981833938440231869708540912726426077854139074815614662520927787846215053205525940759153314505223025505442510731292921859025604849561782081396257472423479074852861015146758034855277262719972453;
R[267]<=2560'd346640168219967695724023387837901322330270632059918143010196337897304302099973974769569402716286239118281391959513111909867811035177906249876146656078119099001605133430363849160849321463586576732881461655392928802294311250227921516246221927513037400522764080473502807225316407945945709504433244729046824027690698173574309481630184908664307375395762866103159632965803036373898066952691724832257901718753735581386439625025066406045929989813706305400739396120948199229243746073917322105775197437187316803003078186568772368334008877714378258640786813809147051242230003159166846032787113185601994659966501439638076133556315814831641026738014354505095846152901118229160205757509778099920413106894036888730690742032660380748623383679731791915025401320096265468966739965625668199;
R[268]<=2560'd317866326131373709020705569256071342791035737463972512754120581260180953104973912248487090412693658973698119485052389126730321915408114693447517541964137001876916986879100316895249544718831125774667537838928659843114593275346046541561270443015770559574229430607567049055285205816552018972058978197392324045676314710223938027720523508000218412316355348425626915866702767496997090061798412156111966829163820511080308321493531552024146807450640850014418133023102607900484661131489312684008119505572341377652342245424184847264851559240847911740976410349715125628764223047437730776400845520510432123185912253026011841024644493183169272346032391026262052074836214833024480616490929136234084130648508070001742036221215121456761954087348903343666655066123188099622204488056071480;
R[269]<=2560'd317866326131372169629121498390341055738567626568848569981339298389951892046496115004356882737688589055998903270657606190163513676637972636207188417938703645682483444834394364722585965776988060468320743899369830133506987074219835578249421631182462614616708266436014230465984609829624717937885000167921955336587567376628451032227460720024559105771843780165248685847936334463326157791382625726603931309946166145166227693627379257772410171912449268351556723628695626249120869493328870661625671963827984107433425468703993520529852233472311282272693679506875421850789874492649568568730883503527699593995230376446578526787404700523391134977636291082700123132904570453742502693992010677247706845959746446911210506224372810650782885709686574592630142142818430070621860730657215542;
R[270]<=2560'd346640168219941526067094183120486442460044670011671209123748445162772901709143233992884231559792232401213712773681156733321058968668291373374826935322591310617546755759528449269275972079191769536278729910773580764818623220764100492753879688106217933475392077176163908940988671669068407950577317279698458944214578591188069279120783225293551455851372445754976797059000878335845979464958373628854440447687068270106556536094455097962092496310592783076031534755830048116666211961069780850045061854595218190496903626135270896241214988790191835052127516458972768672940807975921207619765195300652816575837717068807309412178176700573345221184221703017274369348364618613008729308178904727731185604394090156527032181436101913417257810207853131220492415345638324305529405505688692850;
R[271]<=2560'd346640168219941423440994695388673674970861538480437742572954911755834640999677859370017120364862099573734273079309830555978080254361301302454799858915400500694080217996506126974020534749002830786850960670707935346038938648816460456413020659276252177828726305657014326792903421202708944826372484104943692036883251152148729822891576343403009659668970132738173260611618405632461647333494866086665805238532288292699559622362976660645775315482603585811694882271581824381451802812016984373543546228767749001330322636902684761846793767298328987523054000664236572890784735906930263137645038140819568494002797483743850899522558251917286438263146109494783738933432826148928853160993305338607921588837727226466871223965708273646183298552369817602657386150157954289541985826494564419;
R[272]<=2560'd346640168219941429855120178691379718157478282116332341518685644960692343958946307958976030395751752760495613564162285873061569569864894338252876610634171077147950755385256405782169690187035031274651970417045622035183479509786633092115102003934211530264154399232103328132909786176793211571149636416595498816974219857648635898233769469642928300995276876790785987778456452209328162864986406740948000055823008515738518620623291939154700078407654049433747566056058311476615557313004241819883869049117899086193747697224933478238583880860203342608423678508761344830739397860081520845201672410087536219956293736512943361873463539741364629472265484127319188050357392002362120167561706655043686391771932815450985636084725779456222010653679717726416352204390138700923321673549042994;
R[273]<=2560'd346640168219941423841871803414559040563734786353701479427516430380958370776710023909231036352708118859362960048527409719703492167418760845613875918122509418934288851741603489584840401440520424916489088288072869414779826743530768901587257603101409340147502736592775863431637164237763319710321739434795691793823246584612777465541296265255946276384602297945714315693165187692982342161714417127330247528815026537206841553640521410999960818004983191595435716918992182096806394203707800429132394287144058471525502799536282859712274430817238598618201313505877768945803556386301909397947230222273678186808064902795038024780627908445918727534414871952820279933778330636078893025994271535991106758235390847493389595861974191244621786422618612360190490810120226235092965701779773525;
R[274]<=2560'd346640168219941423442554528493832761650162216195837371228787610107897164055741749848768909835793370228351917014102222296401549235537070608137678544614061035056009340656920640978058369793007942125711041897883746106220231316947130568703838504893789354381152385493340961641265413288694435005024734153353116041279606019028173383921056465827028635277937911816473240024690260864377474331848239091738319284594308708731671779827227271696613535806662780481490245167827303744980855383615117131871108870877539979919245437055418308241569862042481277287327033840139704678965974316737148658231003848654813416995863359367142805220413227613662054800311663854885887941202298855349536454189413114628699363937400936683384517485459160749488047581556952408513270721165539747881510901419523540;
R[275]<=2560'd346640168219941423466043779959757836880372367462252932057512650323098710441307137612860939439260998008591484665461952330007766523381650147078312537097996550591354997599460635126256504254276236320567261547677870619668708558184419885022471639782072894073626547637716027768214289712155694880066482827359198051396560678078223169015923276125939992180440938064306292323824919536594448145089016880329461320345487146599584317409678387389784708677081443541111396054744808007387106204112522919907870646930052205111952110785113153282302659447571427117067454084762494379003776300913489825073316698693972878988612815288903496121269180834761046211201583575328316391395491207055773408083566388162078226852189150719726642203947818450156705974204319592174761743095659530682010332164610212;
R[276]<=2560'd346646779856450751857978168738421071874992090557683622324565210425275210824902107483084426232168323000418237538673577926862829091447305975004234738975272672962007157307755805216826902103928037330185670953137955312625427386399346680032636279188940785223628658084687297921614266310723560844979225032463221870856430857689235671777869826206202762767745968297663056418962385407954731809166460001515514576017149999024529491556362555326544465242723323054840639047706462391104360163183058179681623901523631594516968194026194396507001563477898573244789836890746870540370901034135044480078587511872331260520277891031721827833121457155482962548304171923978492749828773758205202379331033063279226959217487262845878333640602127226175877665589749248593555506393448423453685353828149077;
R[277]<=2560'd346753005101312549110737914697399139191476068817335459430674301700374147417746109200476848300060997907357385864042801900679764472376356220869380239787398120109603967606963192266681130674934249280927336694072416654930238810052509985065311740851759647901859185116247204536499264916341219726560297961751718618645262461846986089766860208692431850682575168378563573389593463147989485637597799076553766115362133086260226984758209663620743637861192329662790925256979937900191107798877281357396690140405254271563662852718467632246016212293903260805564389601588329439105189420643872291666410873369347553251668584594532127269364084083170923120928890516875753134928693648067075650120933917031595245641451134639573461585248047343832342830340246705301223176125174891534938743140693909;
R[278]<=2560'd375526848904936542061070959929113125243271667737286424408178202803930490995287844971989714220149860767566764421489704351953446053639879187790372014223643969715948981547164145044843857816035041842480247108442207248299442280315410681276497170162894489448953343009515494897462500667772871280565618207090033629991508283636772876879884438132367938088160594969179820330049294641820226604151101614504897671076869059531353715558123214624572055853501411550720390292325759990059026058840115196175379185150351571696399540075118847860959896885529761906655570018114836832509907012531845653993422297274358545431632051578409511528860607101053806734476550002791250115147145313254626939959595440106570453269535609168472278351082246586744317867697853513768900679579740803581754791698038602;
R[279]<=2560'd375526848904936542061070959929113125243356558062184471727556469815282639862125110714749944170053562055519536578148746815954351172453836391371805600201614639656413806221015631703404389589966066499783793091037316234243978585762600812450467054081537582666506969361034581233065856581076184976639205191211771179141350362215794119324234944626159935943372824555028088486825481234783283387075694420092562555425979101182545093399766744762687790236148667594564401481933433012127005436232854943235343831589943567212530606839972928961232075585952349651811972251301620612259312459575200117860814727495801586456759261726362072270237063985931431684423693354626862531961591163706666570047725022036941474113539195629417550911038911364822201303578043022216002186650253407083595221718969156;
R[280]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494853594973324418037622686313693593358238051170012062464041867230118212483527281286864788416228772874639601852980248998821199082686379191084733823742999823656052126846488622488741790480602482460006261545693042112718059375236352043337112670844691002800515041085323731352984359013246360278557436737379394237687519771289690459630515509745233421572971695529101187214911111841472825924538593736903265524184422899911093116161256489101373512313358725988873129685561943375946678911072101634962642841521818381033463991759447827022348103285408113136603412568772523979541130837124024;
R[281]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494855063361131593037895801483267854389997255003041355006999126353976370218728310620279818993590975721927371185047246354939847082523495707082547002584755880644674922467693176241950503125752531872141825561385964302519795291444193158007629478790612182980570581024220511078495508214967756376470973080474830453173243363727256261740842703831907329384490362157787250249012900539230486787103887151972606759287571168994147128439276273391586815657945377932731353745965955578239523714695665480030991725041096918461508253874229067344378700784221508071199078332483573573113480745674351;
R[282]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494877175553992581272394017848683528875632357189770533725794980943322421076844486279058209504834063973999053813282321525127532605613062140456722339123253829199702771355682227955809910237209825411559259303336472022448147416922761002429507537024922826379787517886068849446060909047039765420767421319700906159391410103493572730010552816855815295539070104458412992571153909747604925780042204381948401650639319522959325497489532385042146349269567847687988228631949569074680560154813355331920319795927511663128775987844321223226763957890026771118316853488811944545377060095969335;
R[283]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494877175553992581272394017848683528875632357189770533725794980943322421076857001336697503031653038868716243434050234203525358684628095887447890049855679068587827060340518995435530845556785934640923981192220717886397523854155240364046246960885172841661185834369497533908589683788491700555041500200469799356172223100232742861828169960256775918733459861669754927482479591731195437587015241057983962472110925595411507102218322991528819467677184882413330145175115580959336527665133649259570925767148112441031080054342233862335869217504690995054596056326689228916579854515215010;
R[284]<=2560'd375526848904936638274513042574841585385939390720155658278129085107062466460973405550289061933033461629854640298297634990751872741010575431502700583342397701138265397156626527586783838459992523631222579702706463348540403118359670849941038229269338287636559792358013101001514962560101023381525290339120222757799010146001475316762347664082567115526842535024904775625857086810839616856214176069178972814887625036175281887941316563485488924599294999855526243361610523152242576701370517185613227985363356266553645845212682348147101344382460447759609608182784378487848496863842309184338579166849177072127720536522904776871412693935903890858813951771340582320337582173247940678295374674226140455826931501575994438224997635101970788891130484307906553103497467597984044905727035706;
R[285]<=2560'd375526848904936644287853172740199614144856102681427696213128261632665700484189713031357621256769955389002239107995907746991765745071346083533367056390654680314511931023935078965120736956280927588092261406964856636747290708534894661258092120183593800494161464679249624444017470690907951630181418347394686711796292517121015156438989369162518590241598547615056056392628121169123314926355737141835083358565723079887737236454323284970885854774148873428864839809947895686897307647063740284422723094381147263814585899869567732793203251145445230303917618378716497522255806002186604945321590720988247827257924476608712912361194022415293971172672526994295600462900263577420523375285833110604810238983822570348281163345421266642133434065409074530824607700886407595725747878318489394;
R[286]<=2560'd375526848911662246517982153134617052975304416381590896504923851151332796304781635856389027283550332793966679240266554429603083007597096659450916058003011348561872845159795094992562156833156793872937272872301359058512886443561627221479831225149912647365361302336533837716967547142678569852959332098967882693479709145762774094466429997123318803274272410096659593903171572409974652135466483983750632287283187925949530151983012882033301375766536535641232878354308158945295794185660977257087236882632494274159454151658712937593602219041110994940542372236952199859992588977185824163478011033538955858558549739284102028501016049533844846347531638563237820743755797611744334201056690747920570013932101402894492425104098979764557730484378272591698995743323063675389911946208177286;
R[287]<=2560'd404406917953422338678295327520918644765738169333448693901246192958099761268385534562352411921086031334826724184544445157628807384759159267423089530407927320391442142725679662140427581561749684960693807719528874284810270623158308247948934629463036651489843851814143475510170700392618020734429135306178452932773324723480878957476221233954478965472168072254980925851572435637617322648423178888072247338887011719777440854345857986430647686244632920796854622436879686220912320364767151529215896313615876748466984432316175992525821023686569894942464055092259455111535404889841644334794284823618324530274775855406100732914016245091150903166936494249944929442676210137180584586619866231882112019515461909341298583647950156793273249228079725574836883395698097604821267972366440551;
R[288]<=2560'd404413529589931660681153339969057251803798294552882071480317662181396680631593414512921025891802237229921890829520912143143387438132091166917410186123206365618983733026977927446897035443097079799331147974738889346152543296373643308062912169691142721569695538994623060524531230847093599000205146838986055434479816355706378535943935117401811853623858475654717968951389078516570809849254673241613551774405823528382888084410886775976567595696995071589211699164450181334069603966757953211184340697574865791002576247347208514413290913641232809548945503087350498351613490302432450956671197569473613802907147993888217705555080633731168314728409518137731291110802092177364189240660673719034388780967093339207847786681769709336116665307868756181407456649977518465275700279391467671;
R[289]<=2560'd404413529589931660681153339968715438207688671930850276148719930130964996761180373215478956642378300763593738147011417367598189972055709499568907053452740900893048967382217141932486495272696734262801068803910781558819925499954481574867164776370593874483303062618752119385049767915322959482324192601067304652085081435561852229586872244882545535930579209298304954394129081421400756758874575884476976607692363963428402784776185242683018632584868627875166860896160407242500170798797879343454717859425718251482352798237041084811452126964118395702430866258525033814463615471730422846614352540319111451645646523209549835983345762881790419055108276608730618968130457334899592726422189869199123171773139236377435543824431924269692732665243848841591501848427138712595949752926381974;
R[290]<=2560'd404413529589931660681153341462121827184982211345178075547046525660889453344265628440907000880542374244759382731728703961258427277122136380751400891741209860574247691838276737552313492740479798213366684542976499548679383671903866549740177015631899596955149482697733717303652067881210853607779269548930283865728105598045612017444344079128790154766612888744906274003005022219232220398282974919405365541198896209064383904190641581182195561577526556834478569806260991319809583113001872630858597779015181333837461920418339622318965486937997636860504591205032914603565875002590659253550809338374523998895462825553177761925770536854742206013667369524415743177262013714217582986982562597358488998129678933277748039372657201744909472254953817493332324041797580987939467521100872295;
R[291]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161632797304173338505320360264687648792156264386749475057482385742176279422131287517768371354204537469586621447702483005860541522903143097493829280059111038401930075963492848979250059492526998407693639130213459368257481439999469944450927663258385724614225000101666458721295390321395116722785825634165992356694083697437296228089626714022808571889460093281516487842991837958042466605864670641134853478640159108262083624156593887025680011282893368620576538741271222416735161634439360933634529764924346172150418711096566024701490607207823264589050862751628250571617184000450575724453;
R[292]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161632706732631379897511860480348034033710810823793173432692340833814553048585908025066517617754971832937943883007598349334823992839664322615512264293028367242808123676638357649479909180341909490090328835571006317978425332954918686811463900739822437072601074878560220462356132725811000458850644128372768568739385669387531225796056256381514513982994977253909854247356884683186563232523161081071310399955543150575610156681558175646035157482786663716294103326535245276798005692530654105447317256744918871339630037141154454285420711957592097414272582845067560004784570731198322356114;
R[293]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844676142733623174940827834796563416718013547270614521238759817916105108331283439886616553558245742860461898180278185985465142785224388588716628434724255262019740193667104000193024377774961497329224485621471220682326505291180046918897359852794380948366306345280520167420503641409945266640313228756897370876384303855036024369114239965388963490460238977604448809671178230844407620804690632092610986863113583368508804442343816595200311903772140995375140705612176050217293330779210475253642881166681136915087561905755358628676289744768980096933487485918956873881756878499;
R[294]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844653736913811544692612081942423866028625065493264659036889871519715438371601485240993626306941381436679663271277777485736367596314558173820325567892604219160749256865726952466264160709125536926886936575971917995679237469213420309335162174530313899817110737947230037191794200605581120715679079182413414314975448749131520388966955185416991219994806043812127674681138240798391783686864739504238546215658569680400485547358388880751006896322416388823125330623052442086298591610554300011778947324319130851030758648329772449936806356543306337760376015633336958614426514903;
R[295]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246072931639215390443848271533286048834924596025928654661783643280296215054381330893291603834399348136915163182286185759461235032146674305013893090033664028443071675825710842293151280235025867366856139856005672335579022400805886215667403854500264178505191106733682106482612632688337485785140013975890405545244281190809606978035883853798216891837892603529666910396820514811438333137492392068906956670670154112913797422316986089801411687345746609574264012683292582380322783314236626150809727514343016544167582017600491487222851065024617417635661678692309225368551849195947110;
R[296]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246426640349237838960509550446830345975096606929751977480177359356807724041339168177124908860167697287170178778982387692075336690182594321175979117171653857191168333357378346917526828941184638801538925922326899800810784054115907517498103975445475760335368140951674352552864728184579919532538239630534247404131197087148663516348606585023260962098586928743765170855990330363482903134206244768574089370720101608846867668523874076682853969251551209316354369042672782999950648470207233866140792826686164472233142526528019326394708274321469717493405359801580429766756753234975059;
R[297]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448838917852190430297572083107538019587064486503949825140062310809595008755341407523250826429426491735622845468864822380140679601098802283362650580983060204029021490553945256118245488681051596068002975106981513048427293811887830174721385931332253857531363996959751079882980199187785035333358415295048666220592175000598059815572658397745234700449115923626238814766517131784244210230475593092993947998788878581835396027901457227734960998591877988481907966512658270388611285543139947224815968950936719889088398949182509394729585307514976922430579248362122533950491407740724;
R[298]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844316336775632503259831559940060471529686397760996388758986123723960539895947616719664172904749838482759663600543969309502601039572168779708238688985330340554455575577205547516230874362877110943701699304768958093763791228025320195062958053733413185657354192572148800684885280399326397066358230292564180597431077892713156012155074289150236342508573776445522460934827473506206260508101036068841100135815888625837984504135623511492624216850718482219884081354793607876137723051290963180571289698774535415119558016304478565194052326189390230524514339607314160597773278612;
R[299]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844674829892618587231283605607383497904680299009768927568811248048903997053833185832604125789713988795172249935638794286551859051928974624350949694873637555454977353646964454129466334746320573493385922572249893927569605311366339451140063271112796979829846335666379983470351014844671932590818978424320050513793320605267599149265745189732100905838274925569399963343115827200167422152865702361681716298393696339490448596499015564591251495399931194950407318063245989670045066083790190961829692016884752710697747248808273415318970305610928661319757696753427085360148026982;
R[300]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535541563654133905800754206988663969067049801960913146019697728449270502074954609083448231962077513974345785184468028484289379250268367429475595505293878581160075811266576630711683684781921785098796244870244225628583825261750181999253968155271096271460772895972753755295761793806273807279571574173842552598508530817312029542283414791206787015916304316716760914933574152861304574526432528183985353591187742106873536171944595916593427511348441189116797927941777803190742776981946900590269990945014936980366832002032492179577767255364757035265949655876982099774098556889659171052191790897781;
R[301]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535541952655944566313077403875600004954645149336364241453498937755187716667208456536884651027007902291689519079404789068466565998593154692378926880264162728223744986394398752962113521719869885249051322363515342208021626983843012073333218370413186730763026791250575931239347412779968060258539737308075348116425753427607020616586340992432151058776294367380150743163907205556764369915338169117339504056060586646429755014655373166214539121432131776506937088459389847201664339566253310517478705603538449520341379972076208391065245867481445098585280144369473802786691889188296032177547243320883;
R[302]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535541952655944566313077403875600004954645149336364241453498937755187716667208456536884651027007902291689519079449819817789316740407910720423258757347631126605825200585407029541898255443844294811222040611150727664616701891938805736741273562927055820348013134799549628915464347276415986052048088863332730650600603805666045050863275322472868215442530973765524297454878968804166625452077077155193978544452696167620954666989720043868545223045946560376915297582976312465802062537773272989354887750076743894104684632080145926526993994408327371593237189888439482413568077424952443838917198376882;
R[303]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535442368192415475158339021907805228676352188988276005872525238499602416995884217956468028100870434580676080525013723908444438088927202157052721183284266781942399023806495100232112856950176746455734626668115375671735225134862133450728265228556486241580075413057631594554915586915951959483231511073902325612688312768983658526538923319382770444743159734128301207212125225360993263307102420253161764574683985175286934483670602429568709626885128287827893626280844729843119869206164497911755209380730952764976736895240998711785252615520826932643787683594531266015623842138068934709523057729433;
R[304]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884786918772746607248630063638125591701522177586947813585754063763754119526803657654198388038233665292022769214421311743688426508558495535451173978779975903949971957786458063996055333194229874637484765107585092761714103963865951395485150889251432732140175175859506490182444871042385319656985626487240037775155384034456472467210791457117291804199833082825577587295172264959555652468120986492478922377776573629201414219642458551223195494021704488755664777542795474146682811672253774138269371973114711125909138662209312108017744008234265230824199820566030134738185355146330487799426904934787643751;
R[305]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675970526915284467228490168625416888505441888996699767798197702261641219170657290040032549711697761062563939503018383178442739468219722906316537220457078280513378718184247729520441668702741192181174309718808179863229875514513615139849634486853993223703082858185040903056651581375775934442247606531352321116180198555384837762945870798913482241542708356182119994038885497856500627660252751848190410852340435378235915724111359650951665662219753201861111542572063044720179514719793476025648750940747870043830567790327562662519171081836105584836992003789689061656157472726739872046686530224952567;
R[306]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675562628952669309858681756085329484869553923410930354858529430110763831716913208814646062206238745260680521256028418760838880638831308062801231851089586049189443561434854342949528286366516080085752767401756087043957649476334537181793978744266246397429071335757943377170860127453678585926200908943424929143604529809489095642369962512811771198504290340357855872889900933688202518531669736943557659463852381278293804927004084354305832616264357369015793586582456788822319769382271730064119461525050633526223236366845818290847049824525417451021957841162924737501115310027500470098840917456055238;
R[307]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755167965559517919196475625281290551872680513179379522030123885103672500482379145671718424229056075155498202413012573323302031836317168123352698286565592609570543656776157225222983689259941952151287059970039694941414779038414590882965184955264434105330885337288534540578996387938028590730333441960204576323107197754350364948204260047779421750526492422489894097631570377003406638009891237305352973564661956860761999725075895176398380366877275306642231385177220918616463867572167202764447156865863003994010847802920469060543092400737812016396473214839426107974666888693022508868808617;
R[308]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812139508572253375677003716853745000899127754906748380433443460511189065738091329848456795018665833920600786440269700206694275226284331302380107852731359265431820903647818783597571951136860503942982543211022443623062605309041959371621396320950430829374619269505677603554630189083588661647807036947321086722380781837777035217152538715462488553605089233959226550469198509035197323046384257489364191830134214167270826092636528921197630969917025546996370314445777129028334820644793872536684086971224207113948031625439012192774077231295043450107731515891772024841476003106313158829085760625390204440450580560363;
R[309]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812139508572255150848937018018618407110502215287371764859672728996302502058491948238655489260158715914224540885598980540752505679797955387736641219187677682346200013104571035609211456457491277970825962791458203330556481177602775599305416065985448719225145333244759887192089163217983936515132713837309498412937050448310623989133632675915873779188269701242610398402537875057088611847456436007857594336550773620951325665347424328750263687455799690781352815782679291787177974497140336948697187052373617179350164184586129974440961334236409433854148492973691172910361767176876073949755602189314994960418901169515;
R[310]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616781760445790646618040839865459165372038106739100361418941450962204717301885497760834754816512346519394863179203521381114723037035913801363634817494907872434297995279201274298996159444093766275729196060338852896862374770582400413243630151920722123612327368949584681219983710922798531328996284609923855314978922612065551930961798510450986946949382887384955037431016490627578746346622486951467998372090395389751873898398749291169747465077592831582547575358148934597579751785521970781364073527007553315486516097533455910640517262951824102085786791135196053940806695101814009162912655019394237301511975888823623643891970907514240040334943;
R[311]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616781760445790646618040839865459165372147601014696432140017732814663290498104341781313774052165590006900585471873725661042276522177816352662397657932962621343939996721145478263058040764099214063599051126673645006989337860732446277439783636088613217638013153425357216929690004644335100804335469183304271673727769662034715356700764623240752357140142767637814632733730832382553406435502824472505506326977363687196559395420213840121245048265260847974711885292013428095519315024871179355608485995703307003024342698236567750050015845196658268095715874214029928103385896792262367569543291548229883499054788685003458076556137886616402883663144;
R[312]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599302624438591986909246128863467631482100141953692261112452278383727508082112759455340313904636544104148941974123101011438710890249284387064694837438888345228445060892796927760058461083599318802527780713105705423019782426119238169411820451565317016103469735053499552426109768074296257964114346522453177306389675039277500542925866826848443877266806531417001610064095443968836669023508344287560849699483247924532267792703320606525527255702352123871401837176625419157093858891128072629753970584765300449922276457317628444955816050502130247608975360090221179912201691260532443277467106491185842927077646583700735073516446248844916185947461279791042794959080811059;
R[313]<=2560'd404413529589931660681061586573583057359943787621700564892669300699875961960097390194786178283224806505599264804503280588086674922657743325713196909931691566316229483773462487293911375321863444426322534560611297044187445398426888869199527686209227041187697819197545697373933634981122225389284758903164504233284399218757951127125295704850142717125550802069696633508274554777737870032817120502840331569999358733716408135757266075777176319033112444318006908757956383516661132797053426987096340984911795823943672452816783070548019350060933253294656358833249543264191059651590178981132132783905393510599979629627425739840098223582345637903165393777142977340146131796712761887229214853113245234103881093450211446604003114462996504706308202251482638507166133903735901815550225860;
R[314]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891333810565158570704129969518314848697015724982659879427559746158009388013601955764841113616541325795220701273398285045762641026734870647355774403996779829187578179413675872955426357807525529716092268747229050198475310135132741863480836042958211061239005971773611120887802878937606145157391085658988934394112569198360798466675926547108767063069102947289009410275711110880598481869944744252569411832250103536446211883100976687584660394386078852370044331663572593532672070029623769290963017469501148977488560804313771305309390590912716141021513932224152490978148100733027218185942583159357889539857457674159913416760885256260563514521090694199818594922229;
R[315]<=2560'd431494792732114584387480574149317485255490041294284684974500337501065006291637059915277668864186200872780094386098273983693941536094621403663692779131675953962003668961977645849894000378519049692837155687305256672635560103681728419973096542336738908224044584211322424620156784375760909532583189762209575244450287752245065469035097413306400416931705946637759308027901621823181819086661737450523752122023926936423322830818564497766882774253010813328877019084285737509485457730026280204382250212817608719936173247588114356299450890096777498377744208455986876650857206031323064661852789736136050456799010627912458966191767635010852721088598248585939415870829994608032169136028143693977998040385137909160309669192182401884474033764391696778074615539807693521214213139913145236;
R[316]<=2560'd404413529589931660681153341462121827185061796024770072398936659000629969094484870217245482116916839127568920174112160645243664609048268820276378026849757937983240807293048600774666637599040350154898055299663093376195362802633086577109499460894835153367592564536168319377087537377624311717682735771643934632044634905481065652906064632345496543449961382145385033902918956043428158319171798598348799483685757626548952980316418504922615497481807602218642691005360642817284443922254156205167105339976793284302220085086453832112259180084010735418308814792344701163555432982815332005618861641901514419676448461800001555929161099775570892629515263702903032908185478057376488766233672136066752768958959000685811208943389411478172906051863437432203706330212970437498810548184561521;
R[317]<=2560'd433300210274926779301235722995130523563559176473396597794481591035129169500099323929517723136182285162502096329866484160812527451337011599712092149760715004939288387712093087940495231132312223870148741971332835985604474502680108873760630159979910139015963637591348460756405824472552388577966140010442107876030975349135730762317010315241725053699913441611952847839293538285349846843617288321542930872882963154494063950126855438745928308648722665250910306709219054090071216608646464368580396170717885261272742680932612692339920264347658268941325936221610056360058218695147139690013470052985540534492994458221012664296595899995712879390150357215998323918004242660541317025263101393061308980452171706248094261995516460908883347006242380798256561637953593600164617062116966693;
R[318]<=2560'd317753487528640956892551930832204555597846079656674801854503038627670948137425102346775266764593919889881439196463828188569009415156449992055026111409179918129193292070290047246652767743838143641120156126220495202066788611444422203252148759968195151615068063270793035105727439671611945222186511189885028335094983780474130707679377286477215567416404086318905046371037656988629815706555024123081718781433786041377464058996450254394474917104432172980701567635004566952441292348845721692593123063773794163916320272677173538071098184515040124107099156477709750783618749884739421796634188491734412672250358687464094006888413905181596019549491099833695218970062338770652615795141162503290313933033636300745561320470797695384050839268631641632895154618000231517191094283369214840;
R[319]<=2560'd375413597081230582857346831035717323606014621746355866405339981407251057172005372460804974842727197084480530474266708636934391090156766453127377951635945976145970367372055955216571093313714004428295503381572485332940164859848030008368051020364590780758230594008288413724944343710124723809234884958625725980294811584965055592069662730157728778404107475034254253500177240892335111460551882273083713336707857725687318286941984276240140252306072741180074175735889320587868429254628572366403596001258264456533866379781835857952105451355334061309367284523169989624078340338183379260557351682256984019471129631157841478009913006988541473502588742079906435968617857062709960177028282627093885268353788032659750757799857682598899234024759868006008922400270320720124186764285146497;
R[320]<=2560'd433300210274926779301229606002561277805177390418715604256895368230825532602404728680887210441346039035044260345808895320896412922180909825623743111551747626493642125548271651736680456922490183723781949906467190077645259274783764180421810750283291421320480207428155737375132626619475370156652748794020737066844813989899766333024163011016530887560502685983564690564059801247429965343925316494628563140430074819702592285028019317164497227218233582889483207923813043059282630262902820949557523279690141046623468533709895680384890921497190544347637608085367561065695657796892375275564364052207306777408069712719849311964546357005726969942538034253270554924315261997683300485322773735605009704394857306304011601299705718780024737279501588532256418657404541616060207437469082021;
R[321]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435781088756880804280279923529145790718604549205254747513074568072283939335739006254484424971263740371889830938669363386336216259277288819111376472204431309589508049294954013528240141627611476064957959708577920238155587186774641304951942043411197260010688980930797275062441970370893991647265950591111515319048998863023670834804930375905101669067701114647583134832245506050880460561782853684697102747207852841245729632800553020038830415954321357532951421464701664954747092591697218761630657446136534165041159080940443405716857182462394703129492145049084857788498680674543740167370155580;
R[322]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844676230256356814121797090160771478476203783411205689585342738237236733847281189332292116696557170201411928063451682343754382614361736983243934457525582285813877424118882692197441833432945977977591114098346334725988351222500670390530248444907503436657170202865954295909086951073675598918130884960278905050930498781579795601353509813984059071195833627820920477091454283402556328598021099623050655865248402985442155412059739903807327660778834496841024040108893366511639520865437445803080282815197282836465593281219669361180579459002541118353159742438314786263891432269;
R[323]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844676230256356814121797090160771478476203783411205689585342738236416547811820651494317499585084651097163474719656728147482114369411885251926130637118315677630288869684722708618691755935655559047844656849999682519374482620340038182351769171003298699284489797428841724780679193982035394844578769470321916699678920898091105534216551339962891533730103228980609650753756358729286869348076652347034742308664589394490373383404804902441402993719647453269823973640100966950869153711774290479418118439174283856417977187907252791874312301339506869373325035763641844684300891172;
R[324]<=2560'd433293157862650169164853866944951571924229416956714629858109412911574428452357581147698874498672371781612625910044442468278646454369043048511802016590486675310993815989266793517876318014467727423542942026551479979241488980678095210502005116288850174684288081011110514707599265376504117621948428190105467124963507294445189025304977928501759177009081728845681652868504440009419965434965279436916830429519355545416058909640581420102075135127222215777686011958702137675438704128280387519957566911314019757473306431411311101321789080285849392895834485544209734551586970275384678268979786929519467000678646979942857635926066019644218379965655029227949324002341210003621182130059175033525386662533945794228058477238246599239480246131266216300772678022921386751857021485399737959;
R[325]<=2560'd433299769499159491167711856991994344301688017602532382750661244444877454234461360265723679064092422650743719544979755000462015507105105988628958542809835193048230816212292720658925537712837469175434404640007914687039442826569721111583822345721498768966541224091977579151484308602565284149978143570089132494063307272327845766506530090876693863827658601028390516187633355938789869743237198519711591268102409509209528965144842023373107386521683794035492315036925606804395137575433202323951928532855951652940786093577553304941349361003562667799348982235013527747793603121773229301764042365793611052471696315632636277752138251546937989213231391590120038685696210766011822901881351386734244097761946172319329142025436306680204791208798171073121551520992526513287328985958128632;
R[326]<=2560'd431494792732114584387480574149317485255490041294285843084011235853151415720129661044952032704418535377955157207639433714402264110159923336645226884927689850782529755326214611152488560057897970909065111166401239371018535685781308503610491652312494924716289418145608641564997215128402364017759026202885841523535605982263142281204537187461813863178694965890085178921907757493233899644594694902699658274407781653441854535675669752616965724361475257905714581923073874249175329668910693463982344989292622335143599821197798185210112589169645007999945387846464794753253096948521008139888352961123179681756684441091016502730063362240320126364696175964941316416936183907833036645667601255845084405038962264586864934652575304531222046751514135671250846030009096571842595378949208825;
R[327]<=2560'd433300210274926779301235722995107741553777928745607802858984053485979536310116059254498349561236083454375312419469374466026939394958948285918738379828006836337920358634704735229903905102515909142671425242865458276769724983450076238905592143125877398299086793049108004784535997388217522051856029370276247348463165011035225557159015918584822849725971376838685423051840884836514170390340279023580854256047312744530303825751442650705870787519107908472402567870045629861455080108841985359166614404378871357870852082005866830563449590535115355204397567682801733050354340144484212330192399886947026129515173632460196850416725111470435168250544285803719695917427317994181063606112717358720176255169910606106731711970962728461250611486735475247684987538732032370024089249076334506;
R[328]<=2560'd346633117637056425584457773547598638740955659636760317999214078495307508755185739537016615801349336167167624635431561527572412018758998377300717209984330133638438167447416014164857755545574352134491051417548732356282462517301761596437137128490068629300463371217135465075530036193901624986239499706257176134535381004201649169291840327863378763242298568456821887036008486489332528644992805731210202923011814586600885683834358338440490982508834799900417374963675929329008744745541536844977933257958479945863539602855437354090969584839412637295592648602300171226151359620281182664177399264461744497688028135792635542482347077476446492212326679036028626303647897637228623807500801894456552106660132722006854193085377627093677665302358845836683321606586793021361771422672935607;
R[329]<=2560'd404300250325349881676099252256220749038061102658337381988131624134960799552582350829667743034241355011108365134803152003261052131281094648306590775475239958778992832510889377272800566300243252512793286475734726586530372887455498045765117668034854080166097891423394301800476745539947630909891272329210218527152365486115603927176813130176732215816647560249208999197049777028802221561675514320905990231403820344669521227040001006531531677087732921571207947048512073873998706788288060685546823399392261004939220781196859006021929094442199761185651112429603770640882433779653415223794901740219609241226133326634083783101718817861117976677867188059139696424327463736687729450318796269978408207841749585131096460792469776046497880581093796691061787422513873611063850214196005559;
R[330]<=2560'd404526368186357422863263038264985142427021913713392977891260533612329452237621557229627661075152904778704928643397413194404098324773048374310572934513860259541973991057769197030268535220083502275894109504197116097017128932315453966524343079616991968565875545965985561369061505947159942268968290633995033299003406730405246995734488278456053804541313673778444443495845244596005261484546370272567958275883378970261116157118699204472264839587269264702803908049374436715851220145915137640401635629012460793710190541251745418436150840883752516743596498592791597172330920859401025035240997092001687616162158864731752436671766098698283950380528872990674233995266435055324262100649564531131978486699956754251809047330552624418715528190574867213357974955642579021543647524372264879;
R[331]<=2560'd290785505486316415470037835398202284671782515390475246505358521014301627001719993215521777430072429861685989365446030565084872049594159725210695773449283756055331757479003589558066896629085444056775802647330529619597666905761601133694935334786619503668706795631430643272417754787921396730361606796439182279779656694170031787888096664461170008714395650488065022722414379521860058493249137209969609382938984540618921133977396150834120275210056202468602478444193694626144652645260150081829702260530562831243721627892495953776735121798834637117168420029037084208694903736239283039513094742843801703055962723188385607590148774769066412762809184413775639011220916147229103964593836705615731908456999454972636878874500704579548645483650022366630370779848052528451424992300623837;
R[332]<=2560'd317640678323124956900021618486922458200352481023900943273916685812111872287193094724120787269541878999841065511572321029808558266361611476126582137421668100020833020015596031277640273626451563535552275218791149969906998398148222759667253104562543734165596665098400557142628969247226153049122419114269526497195597457082733090386168358559298886449438422878740983992090814201865503982969067469692131450304319822198277513904041878695871501859116893657576897392457109345345355210234910182990856280529931210844376258722674526605156097864947374063547508169124476221138764187061768776438234506220325271973515771072942815033464223626662928018096794579070199198998195970903270376007176516109198607411191625816968327780255531164383242870605687807101527274597504708975043594058833615;
R[333]<=2560'd288866806850399463467726103192287374466697981464853208674740201937540775869884007675146556869822565364305878895709958181817760636290311378209793481012373222343186767959929838068296256258626848052641524197045224947625433037473236885093791913133920511476395276081667597833362774240064161912184987892953703095705216766501196802618235971978479137553512411785100917993331139337464083624053544397089720984367179660086856148827470240622706844826061707225095232431391813541717152594878442257934807251964166101911700695754532203830913366495810279611802699124005507265552010371599388040506259368779903213854931141481155129814565232977844587042097136705658474655644266130224059118510642889890935658019404775163008658754742516926687152650012618168741834142274399465921132306522168063;
R[334]<=2560'd260093403822096123426765630247844189281134270777768526159257553257896958867218650895763881315600523574864283395024668976891861388357379077026601999692080826489696662859456579353475128368153939861533018529781919447849820841959485312309102312454707346552887459017405871711440750112998901228005864380423046834942417942131050494563843516295526308376186081773252784929190455108510798467716928423748416038115473069355914574395373073090611551288102978855465782684192692043194881317911902500753740176727222564146707057742508266017491568994876481309935085958416166310614844364930346799289820492013297253536393392290149913261327979994160507790133255138127905964651312718547411538812678702895645865698813169330004067422357562522831125437562463430391747487878828255240217826976307965;
R[335]<=2560'd288754409036018423449219204706583623081419355215888099173056554009991689451921694151949152253947628383924743426385907892931393712739648496387270321484383995062727617095431984210361923806863870728983103107620405282645466776255146025184273118034239009091624724800708885112313344338706466716527413263683906335097540291951960737389046912540326917706069999148855497136588294219596000054641152839357480801721022378666447460455958879397171608886337709346832606482866851230146100760820299987225005533666470285128703940330366280377807837499826331467249577166208097561167567742450583797687304278041579714188688084703047857916646937094241790622193554130217706817969201822347854863879606671475761113136855289818682022120824857343648066818357450331560609883549527050425775458032258494;
R[336]<=2560'd259980153713467897998325343683154614318625539291822060800258100328369894236466437075483257669647425588945233608829916564358337407779912116714301128389929957933039248374731146392144603694922320930884199897335158568683335054811681980508448420554430056243973216332258413862091341879561781338081096391918315288356775730706790043302318079302670217432617743079043976242577199794115247228826588345386140533647719200938422446173259604238318493427872592408308697909869409977146246386727473135738180802000931678331383579138761331686719903870146848668541854565187848955490565531719753908631294155389330913114656409349404893262262008656159643746836054557889975704644269022767951973024544882612129053345238748049881129176372869987408362803063364445264054846506260391403362821004378086;
R[337]<=2560'd259973514535172450036360634841930539436535949338713415576736251562922241288387574787557096792719197327813969708543695869229604233984118761523826483202934971927995121941033294318571189588143376364422003852385537021369752604827171665940380225897023397160179900580481757711134558262703072274469831773690724275615148073266940153608226036275958820457697603033147408777194022267697691171424966124765060066301345272997123769965345884505709286716040109858993875152081122779653625485267465116805149121336802212761441763766096556249900232266431597897098595262357944404699878124959568268327523238595721011973567798413312587366285869657137071120643468069205580792967894144545778643578748651349029835937011910210992050720033360834544148201135790156218496488647081107257843486779505143;
R[338]<=2560'd232898863029500490347449143702295660766718213075307989304571907620178717968721413006862097667362099000486504160063170780004734270411241772651284431607345934137115471501546733157842482522445793840702264100243907539435764173160108520177734765879481613577421279451563490030810503096954133003714069884305135827403395738162133205887108336476064548560587963504542046520787302057876877984683186119803875260282105772230856262335922448471843521154471127167526846184105657852561907107644324719834957978318636686241660694486185782553571823859617206048000446865754167936962935988637701715999841491863629534397163175954027003620399679846618404804177319664546947002131821371286220200966028050222152070246968704739263532071400139952031045055738493176208335729853991378126231914024008111;
R[339]<=2560'd259867728344325507431996863011170381769443598006806237404419437838238401031893336509151502788923019394442898937433483375846379113496707447092368502640747668273746054070290394608814163744748222054454082372822806671318944463474638097965374149668218657107909224114312618430982957461357642283864790127467994913651648079884207566400199075542726157095337181961484489794020290392154110146488017350941150553968167022897241140353290091286729599706844440958353575314049466747746816617568926967522776460170436899007762329726260316854507257894261197583607893450209406967729351534013902535709245644208663979109146912896035039240864189768018164756176991791168838561447800960481307406564141558489937806389674286533912376502472444811254869227147201241588645094938261410882348688242154447;
R[340]<=2560'd204117970338287737194651345491710339553356400652397168817675059860073059502727126619360854184715202046196542309021369742474238839827875013972192238476913700885366996409855551509659826843078136987694945200801485979718886574737802866795285467115341198239828852404326308395580294911162554084047689013969203760807550855162892649409912179502166434188616473856609519451494969545033414760165657604592391393594375181544072220376645564424589285382687163910356902356162462097178654097976628129329561581629282373176067320996833099662047844229550055558468149291405715003623872118659235711942775858806015217095840979590248157239775000973393399536302772226537743056825806417758126890462699444851952135253934193388087368937173886595261470443567257522239060951942839487866895326632607595;
R[341]<=2560'd286948989771425881125445867288783282356096571927165994798579090108828987102778461818987380986714960616871496602846836737845706378469120129202391167183506810220697614983690148546474972668138211800010701348637827913021836308046321715879009268769772288477931112051564208978723425426844650257693804980465138994102649858809002129733060392870014643120959382581665117700563931473397432250034186825208367279196399513981958099816141405371786033142921768489346416229673627345750499221727936795117988507509427503017805777950722207708992451955739740602678125308969466126468330551395969817645946481282182303529380390319855788190678395578062962152747616284323022441754470204681416677545664001896764072536750665514926025409674482880107906974248461749768266701965101502082584233951358890;
R[342]<=2560'd205929970260374510419790256314965470537329742921112206748586067058316465496242435629322036930471595604751637568910153733373565944611271139775728020263613348014891494483727936075183429158702263047103154390545396905060927176606175222649504912277514229438321698266702270824860668616489753597067664127929440546748620078442213704991577829941608219113854194768919442453731286596958776342628602716288403218313472438474913985187339240940215182545192783827911775737106391777777748361132734179348287302556817410495984036856681443027211186457395891770065975982244383444783662185081353019433470301100519993871727117901960186375630339217986147322103383803866955131623433844499345869366880070071369884141952856050803516295434497983577486776286860285232383391690410707275581041543937976;
R[343]<=2560'd150326718018552426306521993418130752892178764133379066002736153074331546964847293620299066757736753079035432245652916172024584729076936590860395661302454573514482156166637666651052380832228008738236707486834684192515046888442421370299377442912647414283296998292722084379855543429179567976082568554229337372211416321138571420085714543936842362635603277898377313439601893473196186986540085158277625231118638095298257378803181076612605889919348189794889742883868408497464324592752296518702138687950480351070709601030513031831030127490734287889948325390700995828360250832342473788803856038749730604744814527735436935964547967278818041776761218837724415795618282698886778404454860786079651022512266115740835871610657743109795884590442077419976306678885805123702189517631211;
R[344]<=2560'd121923596667169676294134752798367944622349575864731413946524682695792054026606958245036083315470579380851136334436796503224518191758071348909317934231211454581950351174363924050147296802746047941804936273071360821177840782591843810015060847416297791880886602355693100958896567100030126692749796479277641347696872425818687199463438953053368600337608304478764436528882538207429474269825362413774705564938702196191855850787405982756584274283251615877939048663016184828951185481801952092512439204168014757356296954594680253914988770323431118239125953197370483396474151410437912359730817625247700383348118863827860430314703182175337273677444797538702402624138899179621940279063001862786080772103530233902494691132745167496211316927970830119019079689664232606195073861578;
R[345]<=2560'd105793905257971206008549659007166801740410365779760926759815880805736673310563983523959714590906496315108523129381797560699087396712681600283321562502120989121255685528237129570451626998711020095080305480190139736480064839200667258415403644685546475425724373264195072399168780706683253283748863945923002542399573876544322190505461834774051334961433790602504394754948719543049208129152131342389963968071386912793097206644402818042367188008254194532427040467997034029675346313337716759804394415230518373538651059412622779367174073607996594519567638850355317628435444662042472677156545144545026154828017550507893447010326171683413278947579942069313368646386502057271281869747560197049293141271886021949777113294619598598250951920769760111688408896604815131439299949090158;
R[346]<=2560'd27081296589112829943597442389342596363143422228314674255051421046265733304763889582351055786178196464799564804695240966871862658634740541764212263140518892711866705319165451685451773605387814098082655255986929963519539799951746143348991242007385502358143889887603442057507313447221532312779345336971050554394949094073578225376112389846530207060533740598015642846161478578342873604647487974879993476614046637242334028535702614360829258334450459631579497418640333077034439276799189713835553793800838438362699252505285258507838375059632406959435587414477398402988354131827765795177938974635420884827734117328225086568025780696152537386730138071027896403698032949934521126582358909029084601318654005749672559102664852754255818190781429235137148937960501015701019853510561017;
R[347]<=2560'd112407155962532525955949135630592314026079563088828566222804073560207152941579972977704623110106087903863677400258494528635702927381978334228071899234973568451870099941931277922761803719202730310825743045735663668702075520885910932399272825400508448742059236896601617052259568074721360919814159539132757953920493285768298741572282198921069510988001784504105730617176897028704889409491364188570984983629583637596322478951566991038394832780703667482215232405196743042097213427648488100091236101585107867956038595627155055918021531678861657389548798126532600380799265013725735058994923526797812185090410813408551011918469951609367872037669063531522717635782776030136921902237370837655720038720951084897874751519128833930278293735867547499446815193872844420914884861382601;
R[348]<=2560'd1692999895198974024582285182675216451853470162127153238392739948774396004441260349495150492881494428127993793894014548039177669474885185195527883098588506605391280686650780234493292803655414092480686513055273683690462604406896691886907575094702144388530394459039382515260882920794360881678631151979930218693810155293436353883466315871297103028723494117892325402234615253208343673367843304516375832708358322904001472254787174077206019410702321528281710110078829236020501316774123056794046411194777280619277895239899543626110084662681700371815358162900315632898890141712672846285114180377805748698844547900150686132058732724594917360042772820673205635872547001842085508400751948482360492843226730317126156521489773933734532333555655165312442442448368094994753196038441167;
R[349]<=2560'd1693030570715009888017321101032297625663912598853154232497189174803026698255680171823479133095638557460044714190301224621745465452839472710367658795851430593019241045278092689726822046979691208647950100499090539952534708318002869766228017193732797028535813025221159738061474948224905745894501442745321248806039112214655265003424229514378949965211552785067740169551785886294214402260945070054430685431084336615713922124683773555100141667217137399174092116044346606178560348852636115951831185194220537613825543845526699766096225470721260548175096412978606422928348125340424935635713891142692788232887816542835456375556232715155858341642690217766361207212055131795518993329084826061561297935834802948588889262250508945192460337780361715696479713906679833832813994702198175;
R[350]<=2560'd2728813343598131202768395789201858794592203856432392742334877607836741914047880082289382250000241653722214710388048069927274561104482750597799115826022796387383655302064600364179702717947932365043965606676264058704998256376876501136289892712552011972467593283768868766364466061972313530463562633587945761064623675782330077107670115699686386926029178270570142122185562196239642239090296373153945137886495569146361432668732341953711771597537394599089057388360432456098397645966590086106075112243897657014238223032857906591327896691638399587578447821989095620787111442883183081240236250591687916132631225368271079064972713452107656144401327212796953762221030110447844455642664695331048036665229794726512567275363108276027484752101188627116874118173909901652045847787902;
R[351]<=2560'd12333113002719420867311148689805955433277406011584327649923974803810419353893496966109616116807410543280069855712838669120222928735306714623817553762237985758985528558987382953912836898684257415386114097449739437745927249233633755261186076190675955155228157598757497571538096796351333318020083285458607558829380742356226195460759706082307206702475648095751807863744263696863628687065923191783911838982001905034657752166931160914551023089972415577780137888870461202515815545738780713473139045777356709210727729288915065292497759136742380968623016123877529981458350616277854380636809475200583928128278285656046954720316947474702252930639515606787053724253393560381903051291047642656192215191684320453689044859929281329942285389171129643730055359736498459449932374538207;
R[352]<=2560'd3552133755258743967657990599909009815418084399283931847415206028293911493857005480281605188050810709147479860956688611946968873880802730525511572959780051731882170261191252447917544744726946858491021056551589145515712500469415849648204404506707905739358591634042019230040105109940678527489635432957425234698898587932290531789704786527659226231435910565698406810622481673850469825796445487320132778926030222592399411695284286870304572905368412841214706688432844746609284360386427489603223387689604721946423729658563366822474184530443161266902624950116543234903457226542128090889019337691326295479632305647679399938954134075042040662430275641842925484847759669921427797557017458265581886066228680454656016892912713516191985445837281349198447975366389736627827032903116;
R[353]<=2560'd3991086856639054551689892069072562890404150853676608834715350237876460187928713091748839426486610699227357923313795181845602609266546859954021689791375073741451458508802571549906687649203099420141461779431851416670360648781362287763209791942853925946209217513837747074675983429531511614501895605482428305461143705753167837114057510370789666237371696169106477350976291015580210962092345752202788599894283809577381053495869413434206234058381377951398292508137511845363534397160521636187897591838519602918968951269800876711309866793178606533468522030696925945175281028868134156660088254001749651409497012966792438057848624196878625813692734087536995745650352919268260631576246042647509086398263332781738788480072080124754532712347961711087481471854229174282471670135703;
R[354]<=2560'd3991093554435624772174268834097402044400750834298084221335477856287645773781682497286360707118748081758765690266778746916881785020284247994579657335826260232133788871881406891260494134018476965492923962934478283107740480207832668700476765512037504502555861568583321623121808790318655008951331828852593525172703821293548197883884546043043355962666944426873458995046078461344974359565091892560109130352921020106169806349219557695809893244217145272868499191008466869084461636355775975704566378540933337427179783630197561360764700229068883656514810431734138142287144501093700500745988618254443855859577048006988896189213519382482825573238615364661617580944434848670301207376653858976107195910283942653954285681348655770516278619595576670242440491236952033352969598269340;
R[355]<=2560'd3991093135721113904874989031694802555432236361543005264328962763681257021469890977180375116384283851084116126292781659514106758795506504167478869443854842473089950877234066495288537179719461331228343283747333193952328021111507457821555532563205013702370077048257036123169275774727313396378159593395334283140676528606971498289909908266434665588167762213804758708674002295351378975356440544635099344208776788746826283663507443249079985337900537320825544512280012977849456341008982470511245137935355184847210138590100272774553056906653446012279788013048847028987644616511214993283930691865329853946797824971189314707648718633939158806976994403237060542258256176341333114380499870043791506260463494558347061894186378991204609924051956166147784960274400730242901105626266;
R[356]<=2560'd3552032843419607264592048733527003984696903187957225618596092569868990384444659438539224198841467401255776387351755051721104938945531910162701247654605865245717774628608583244287971122699756584194134576470890709582356920874708134906117516995772110301089533568737328198178637718942389825974350825672801487887051562281075840106174488736121530435834983509282843296689989001702000145625376546149899817227854350528842827033634047432958455479418956911496798748715609484426039966817232186308459146443372707687531157964217981421942027287791979771156210228687397128615613543458023003563790983971734736411328235785147266490616057846760716249060539593880250184058945775164509731905932763850647697937195298154285211673080156561383822762090059225634875955040180566446162403749219;
R[357]<=2560'd10575282465504576609102472217361843482831562499149049785835343314671257320094710523831893176866457229421240600153374347519950230740965696050800136076542920692251924724388338129695510033453929570629616555345269981474862892215663550849420107263090452960757926948488597431195004356764271539904164541346439049037109871864004665151447905727995042028515844059101486840771572215925039919332731230468883322960180188482379401254836313122316285083380446235458763378415298200227570138906813840712917070886850691256479727812654062133120189060532396042804131242307355447112267048847446141596708767037564902777918046945781068083173027431821299178524799283592701965858723650075076430995489520607468904201385266391561422764890045822119347665671589788783820267234908191748531788482609;
R[358]<=2560'd11015950621521399553494875255119206882997895760082377196389239781316313535654072772286279616809591544096861818343335591811937295907441567545521375556271195554917874838820925322262193414246882090280019542290940644478909899884280619830470321148409008803748431364653228340272888185009025392827697118145176539792537476068842755921258009330789029408694248750780197547667802413158443311197256074239534474222553894208682294286991591498858269491557095007328996076239906520468054067411061438952055841131465888769419933563095628248560105834195302469757000658081717122076244589187841780324872216723407516407282417905575977594607170036497965229115864636967461348807854660498212753256356631104691331344792415835735258823421341593787494774121761859237105291115723919209654005346852;
R[359]<=2560'd27085252614844220819152009135992921462709273855885601210847826175405970846285970291921076609328020450685225419592886915154072447234832377475807269751335703132050180290488375032488184771013700502553179889283896041239430115154219552605134503085084901526145778550640467060564290832472820657254183077783831090796129987090407004516845172010311424283435594441237816953629552775220560375988282880727124811785801989438866369034741260990916860887765217004629663812266702925725218326623286429351321707169028747396257448554011685470796408181390385357654330043644231505986833164814501301013507410356695391447240228797172710716293941708283966642325460884806668176294199009328178204486452213245649127798402143395526585929502973944295357590555260998263295787886568881842207820499587874;
R[360]<=2560'd1696130979229865920388337671782779100982685860168081108294293922615235986252124766609714697958163293252141045976428474901926030563411376556517017771396390757760517291193169260506017052715061163708229876925871913109891963017907109008067984912977126374145665108746908789599688889339442742225441885627878838899695810859482087049499098598520092887737790486540357796375663200161298820904730673715038060052213543804276489301711889175055420767883678744616384039046487514381452782720369128428321003491432417228187324283854673646382995356435219675758282794068037236707578452201056404015533237812001946531022704206512719440612001348814810488616640185436519354995433884491716631690287113574707687615547474226607391719862352640424520594508042744634015964129168628237476356064097057;
R[361]<=2560'd1697396582020772435414631719023780925733831184081051268360904331849888164764798514516994023875423385620872113832487905633464489215469907573001047297839990127345871068751790740782631645214720227381445636190905220081736978413312994604438104583448356147133377223714071638954887635805025534314560331483686034538438038224771718037086518091559569925070721598157653421961624831193966377459846578515390329672475431982794037040574622863535824397461177098760659216189733258524111574345821364477563035375811356496855205935138962795447428548664977898110523384979220648991729602602866915017311463914483311784248423612213703995375272484356261978586764316486858466794329117862583168652622290471701819621273664435932797088531211759204223626554848051632171574663812062485097578457215490;
R[362]<=2560'd27099250696153734975544971261351739081224006951389935491667522640594009020505444347768333015185021366445626570121629606238536921520263619556489269725474568865739636303646844524812862910833152606095583152329656497821682004676628631939996215377508891892010241388691716927541176151325780272696370018105288718854566161238888331241812876664662284601494826180801470500645456436136456845754330514519299081280785904876831865941274920199442942653888740942926541256017400810241810412920088380906124688234572364149301679514197838122263617889370571965009082490043719758056225016411811321847235464432635815615434199566785625819832992683040799240912340045078060166722047665177669681786215687665721216705635809402895229939294531786441193435629073772188134341349067041240546656694378769;
R[363]<=2560'd28897229850891864504677625664416174121045756967373023518626907929436926240375470720627237812686335383666366722668238739722129762222202459002828444563112781381486465192118798575818083514396303685671779950194597586765685524086683717792825564886886000265574564091659631173756051058619405607992913462291817509683494046315052750987989948537437170840711030138774108386591498122481528976580197203145975064537694580365917330549340132510906702722434336636024633545936710494953136290354753673249630443787704176820460096718171240255821371822038183954988143555571333826334857773127981346024512062683684836262076557095943224277486078192067113902732467268309648039916783741916847061388585273390689853763673745044392131287790728462367790733440032233473766104105354529604160119665402128;
R[364]<=2560'd28785192685863981096640024393222193783890901479067945053108968737868753406465801739360140318938472068559524128108512973403807054181188370140784052425862154766170224981646832807103758064550721305448109806521994317529597815781354810675664617000553406812144860755752473555381461714828198076297526477993554888080853265451785633735260579110133668694865317989421324189412531589297775241977784594672403054887110750033816283941097387536636008590766309633678227666295371147571914950889642286427592558421880976906477577834994881870744622521329650394261248560735940745700984974739968370818691721043799865340471552647397790940018151480663157507484033802113504712518906923992847211699433132371866450990176299044605759984746865231821765388556585209556819036208031580805749469526115089;
R[365]<=2560'd122593517817379262293667314481948975122203673457545125478520527764951318122419504759913074111587743632310493257981722184687858801584659757971370083711596485579161892634544764662799472616044047034337891742305581741904512554168930685266858643522971268864252309356058228497860038225771836553955041893255392044136055239383923751503016991853015475639061276585747693827422636176883008140050368288152373571598685738224230731676840157782742063423894641258664152565867835102452745957873595995677249965100124090671595869569298581308279984110190650197524679214281872519675340133675016792712156030293370188966320605073263044494189326840098595667917803996157209631466311580519492026163291397970217955175290586613094799693603723072187286166476534079259329273545394340163951752459059;
R[366]<=2560'd1718463761589019285729091327524580892852963064205456388991918068840748961118244534278610868731934350131519342836504682111513315950961257308052527576119685100073579550034784771293202810283605544365149270200158474018158052457426252296087643249698315899811734864078380029508099610337391722426152499201626714360023432033149698019237079863928035122465741951557218853442403995055684765708171872505675878750436052789867318989773651351776101379947038255654904953703328638462162509341353122486605256660956002431239897815196836186743024107370208710207173827548763168222130098752935087527133896869112218176829280141112185597653132198195487845163170718566670272175521715494128845477476035430061707828261648991571696723873818477155783915005099907884827814799035875712735935271674436;
R[367]<=2560'd27110602279193046108731751700734888637263113953131959430871538148483242442973003303839845075855862778598180406313650679607040373545712426738293722368353382301164547341374936834598932207091712404299665987374168042191176937957988581233129770144409332909359013594879389430399956348301664645771536130170199731127898629833023045002175143017918393234250561076669939830758990627065069797909543373245157422201081011589021367066610219511673102268858789996049021951951716471065446148435728638524072914336488850387243898245110243949313731567846038312891149110399679328001005213183651481408804703061232651202194709010746570668344037000383770454390486770182586250141472994201172442372756795847370870392049405124239977437675776538592612500698865884900014233944011906066228437923734052;
R[368]<=2560'd94207886959121087612490858808409470463415229070019286885506377404589579189276117698990446946118091919106683551081599138653899664378751677461399955760454573429903431786915642470743222672141900989395004350388173430145968759475440641973486809448458232431889774731663801303322491626907871087033372854971407461344011944703823601039313664367989595332007024372255389029398432262968525624635748325508395051002166327015627495038395366791401232183874922474281471828253669058062852897691234771535060253457197969665647715609430629595499993480776127302677121558742581693665503744504310626141244759833793643935818453172121205179655787687435824156103265544208173922694292324247197119915555393397500534004289198107859871820771619332221905247573066727955;
R[369]<=2560'd5563451585595209175435383911122505377340840879980891704263285051385445040237878840918547365722310176808195909369303320235739285325123582671947654049980668718972307103695274465441780528360902633123466210737150901657679156200796948958747573141567670382746192128175966099020802640793304365646526822803090142296118922223617076332087143958122585037619015712800844632901773786894354077592017674107008225440165242641760944326955840787819798508522591056400830977908448619926103500257890317940000821831778142471218248785412380557486840775699929622114579672747202305270659976324062457604590174035757640604423429154428573020717853968208254748496715219130947309526477609308810197622191238977788690938596978950622249338207319503081365171121062827041;
R[370]<=2560'd1363860345048262215088241904927565987517441519791352188830089625535351440106251729818539483336794563664506017960506187224398933614358741730090217646793946695726161517755547449866853335010736794378881882009399394687886686478009974882680148152696471432111219745404474174390525725761118680081833816163983994324792030758681292226132684574337126125322266973211249796002732639751509738774670967162113959602467076828531105568735917519847921310503292287319453237543115557744693742047673686076276651227268719753565197052831508302470626126007843530001254935120811861244428721319530038242327861375541928434023457772673862171633745986848903922967731854737318577256299085219066788545490822745547001637916168133199862789465611458854759469877961234;
R[371]<=2560'd5349594597284138893475397197186395555973361110600450335076854512773477344679645313987519771398332244921052194331467701814153627970976630438902478140780131912142564876930163183781502326076060100834419364422159857317109320478125319429182964222731586101129291927114046549836758134299420457629018257672362209628247710745704347047102201916911202607360024943000500001216127714210025272676747469141733574589688633707073381383996516784131798886537289380496611216307069570159547562220796411152626746969955657420965413200196388519072512870193554936664531525508371469752320000146509084162671974980990986212184228709837027459799358161813046546241062346432418850578298834183125732690434762831722086341751861414830244170024115068555717037409041;
R[372]<=2560'd3961827782650652179889815946075605491022814887794528312924726310355645306566555434015034027404315357383913740762945270014543983499219206422241742974407426566418802632261314387074311549488309921985303195877718528090698343784612095161133069469634312268772733375650935399126461817696847398743668579895631440419235517341090281186938289140283827481683041001395794671262067695287389612379054589189557069800259230886241186222843457396162547295135271490456519406703500159158215012252758536713017874643922642134337413039642688054757179502442892373817515583211844318799952391261075460205807451069617025614298905265018537328603047547904131086414630075205470503317141894978643470165601955468955481224944990317179440368703116388362327573298;
R[373]<=2560'd91709760534535030514494256056830719852714058692657605663430971258296945741964085205583275306251942846787840649253468771893543538884370494485157372716096516653721929472774860499002539334227515551957087697163704973610612739509871963813161622256206675520821382439325080150684029006646743580017201922299738995369356893956934592801664859645481614000619709717687682556161187966852043626403887980804391584722836001544739044797007099225516636298188092989108365396036383320586141241340249032375446468273896449758092074154921801296470172517827369960326893593695315330143902686618540193353305608217530733033481428396090596406290208457068373826482554692502342908927972125211579513601872042645175868936779251338705343751598526371893289283;
R[374]<=2560'd40842962414425793178489861213563373199150557815541608692936472885052228388569126184507675075825549732779869605947264957489667885927482456189515787102638794543840418025588025873706627725919335038363396104988112882656168811278458550518243260996176613295164397319820317141532587058930148956546240163799853232670729919468963215646480040377811016598538374244697098309738559394194777697670199945770263320704633273465523525580166960699585047553971733532461796619480930520347123199779622896303213561709731624217427446225197822403198584267528639445724719728139510916043336707979049107551736435435592386844318478833276811229686664247082574374931025804068057201829304027005580148473443646313298465127440389289469537052631778479723553;
R[375]<=2560'd82335526130275352263614557147058148533723407360169169932865026235971525594679385954020681535080298945902562814651469200998008206536276055197043406139450075480577859793957530731363946605083756462385771589590398562613640020832159700344846926539538351415364366528728350295598219608144659746708859220800527139816371184713245698282950350190151638531011662943549267081421085857249506084600899276641741984911816922055303824999771749257663239741183134442787057676809919718849872073964015716501391140707207776976067751514798455631434060940538369872647631929889195821412361849917757714527889997720249210249749372456402346935355691196527099945994688510335144909964759757008223777585980205103417050767324888607396248719809636824598;
R[376]<=2560'd2498551612493125614601359651403483896246055022017652562287075779514148421498012378984664288631714968753668874655584918182644573339180446314776485358760457803285402363226191540673643483998395234351341754929038339409632189972104844754064084639075854983442952794566239833083015205124555592251746851218349248496221137721388155305335652467785418228801754358984614534159392655774903895683192179937177459171704782402626613423704809916143481363272393528225734654621631970451514119307462345202431968560000281531024357653086379608612530174462090918780012562478972524033247726994476107727080583576979246039231410857461530723920501469103784072096613935915369771480977686080986978271040688989122958091771745335381331125338198820;
R[377]<=2560'd82834446935425952956021935490075385003572388016321394957728654721455827533536407861031502691714001362725991976769138766795952834467334052828676647239878562170886844926974219098855024498890685380240099522576067633756318929147767976824820025814449299732139428835748490889620756031164721605980735317390369522627099010067046655143901514073693818927014938428464643225538583761920947587634323774519615601193249429217913068059542443264625159076032858942918373455002781472119670791994858586521110420640503862703901720111100413397906125252657566467424184697749664205011361625020479379063761425183924616533683487182652632386835822999578857579071653539403052599735915286999576300041395787962935285169043558548594439703577106;
R[378]<=2560'd13804617961815594851711014422846975149431661813725970009524827363918054724839657823352773314970181042135024513402737592098135298381621867629666946506351001126525955687150623805040307706666688949492988493236478211718681295687010959175775026372731854385507819029204394248453950266411529331620520580647337575107188769061653274163708707867970543797043451174100932901885817211289344003093446717176105495687909947742179366123752994032702763229069567324870868615803965858663349292943507633535900054112011585841729196284380488084915591023799427377308370584365609756005351007420047270529502544120297494221696656432632868152547500490676118702072689244857588198032155611123526970308334254634414238467051257203353188305019153;
R[379]<=2560'd306789551544134128376179870511872544839712287498930687371273659833604631214074030887140863737099472831959634831383389491244189134494729067213346909160848834228142108067419626592216768890743219558492651830642827283136940668817624077713706301971428375246785552270633250783528024567853385285198322802958526690858656876512504760333280328802063769377490674488561950919654531022180806794581977673922787430455348899035621030274069447686715358142680500276171584573733643706228921959433299522855386284066622330343402974991420671470733755925111231660433689613035616485667782941066623987809653265787931873406381981562903168500898168857656794728531854456308768601187128213448509987767784168891152504238967647240792289837073;
R[380]<=2560'd19170232540008487334980743797639608646966933268054318885744736013243385545150267180281705588529782649560046735853255911660257501531194181520520809008320504879197995657814554995477678768449510958974774462213208839418018028990696066613746231806997800535610180764434781350108036539176285058868795625191091443484633540027919985262110649178108224059761787299416339591755928355615713266173943875724328724725091783007794095620738844679097033237211277005512074996936719194047503136906471861595280308041882339545308557718471190906409218133547450017055631026668793265923729859081542057919300603984677737520342137130116269774194286490918766286018451554326306989329224438621745523805805317112856402877417041678105379340304;
R[381]<=2560'd4314298805738624375384353714984128297022971238399432523585413023510232134662943240093027401492130279932567363536682429498271044334570081340949845154143612903629045667507449211561485814058595635092332794543339805338505582803963730680125360824437819037468224392661156239412602714701348058949160998915613089634499116643974130986573201483879302144930630531381455778255731559315190809799509496861438665701972557255891109526578796302077319647120090328214718710030046652731969080932884968492687269736361177289664016320888651359024742193876607438795256597236014351309320818789957355718019449867761877308147762277386282561950409768495042031399924803438019177517129671926895209147908894389256971143167447784378571154259984;
R[382]<=2560'd3214660180265199683942863227724612352812027439309913366863429565282644614055111148738735183287824461331287101249620239899115708420123412900466975926237721776795897989672644617778005284557487697996074336652667646205785845086332243728438011416214092530227396298732343381162590504275522754915097853589546136270047570874162221445902077674629888232419179348803470141524083564527353205935120763514819212737868939604480992580165709574071926584052622068857649683760205852845663455019357745601308380381225447823143711703421718112033014462514640928446420333020688272523303375791919848164450692319973225579502139136731513084822243148137591405954115772648432134920581203018846702210098894334313379981546808705814528;
R[383]<=2560'd4806606856755855836031652021462024729766552838455343717960176765150119940817917220967891254182338477040435319325892709523289962687663981566089902704372625750864358873703607420679952687388194676380146861127304331426530584073670208508665160244761483182732950692498836253470448071414040057147947913523569236832556858852879895717845251542290066599722248691598715448460415418405765894065267057268938102032904929901364920667543436503658305962052409801449840538216049580392033143625687580837868920067867779323417407118570701992414169669492592153519616278258545829677246406367972384700349348414569576482813042533077316475213178831083824950676510004811760968926745185099853434075351539746196521516987568250132305089529796100096;
R[384]<=2560'd24630265345133851684592839489774321983011982656094776659580810676134317120630757126922464337393195083771347477871669559170065977946530026190729056053583745413337322597566514967134315451336490925012066512295580573712385970094756990757983002982131592206668138635543237685589114019073817189961247297596245511322310985361323271922712839619936854038594363490225020395533397008822907767735569011066006704709814920286665635391251075601294063069613156460021122199655597263251684712746378603476494167122472326267555417187644293048756186036899448661932471918244320169655802012659695482674829346685203089351643969443920698356634327989861039724245287717519426138990001667585783099726841965245218877141604981543964595341847837595426877036081990342155323751142576164438016;
R[385]<=2560'd279026978889740021175034252447841360769933350756339039675642147474412079941011156945839486219141801349000467911720244841805384832603022901703601097550459815023997025153712571377097684305189929517755903854717461858697578987882106734056431582840898518742276540637679531342880924969109987104107775885930621726535484166120841605256798421979955768790425111808800843281184016497399412311104056456958352706831089164093836549142473475249129843208850367368169447685182843160913039153994666853488737729091129898875851948288670712761668554450441668504108990584698350655908088730804440456051668456454749307355972001718666125899965833016912884153165282666452404660848687495740045023464013928033171249541534449664;
R[386]<=2560'd23489251465925075230210151185774156554233534484953667317186290388030343354516627258288386761202685744061840848039003501143386996222094433729614747770654120170775727249462034054381434259201992264517972882605176717825714646454999907926888695787576658860618023380054261939908734877287558893015710077458515034355865171322025601518433942722552043197182108751657368265313598727613830628199103814786643941568975440579950756786708546644649796728013552696923548922814039276875858246382129362512681913845016639199755613096464817882145581185367376268218375908000815789261853428251026622897639850369745650033331791867931409366186401276251950685650510862860790425935785654252953472163060080539949331404659226789857834271971470648292520894212682540578830965687713792;
R[387]<=2560'd1635603558075294838429993247367826069184389473256293762549991815096569328450350072700812131654348324725781875806806606016262040819261070973349527915252573930261119332768147461760123255068895278659784785525184122607848229849693896619606936637642811461773176272226182997177689158152694834959064271159807238400467575218496618487977343151339727248960700748594313190464062819022845731242210689406846397083347518918466485294807423471516168781792616454875311629669550813884623582670594809822714205143139031760911448349148290551736441927676691372442452846857587235849237516105861606836659795530445692734760467299107411041173621425494668289603880960539757266697911160099175986189795316420843427217476175974607018896649712921838003340120422585140294552182189805535232;
R[388]<=2560'd1539391584070865730287052468110895123938248916005923541223521647764652063202442912823694578702582639360052793702873417721666200745689061724075961408386008509324890582306957034595621446479549127325686859562583079616327493881997738770669671372178810540447040008018031065210498849687322326721202377254371727286163776208992933929881325607555046561280813049257375941001302303127808740571584855974865025313853908115401464356511521349287083350887654736148820978901599300253155775016700576242156525053810961848478918351684005401645570232717448041082625791356508483687833784840280107266141959711066487036973218349459476403443163828546496254126532340894401724459496500300599504514373001859960667225508235450034745588101841548980548106440404422210946897116788477132800;
R[389]<=2560'd400877108025885365940578713010340976505649656893603798842761879947784953318807136546739696439973422672254228801221841912582381771385705937706316671636594493784934245280466202412304486714616591754843792501393463336470757204638944226096112111100743226896588923819753474454666129511947096424156551994128004253024847775418830670286191612593840438967237197304467159208853712225245271021179206804218994118438582569604773745486194747932848311847275863346972657520567760205952264127554720206749096325338999611983060293335696287725162425730615490972380928375367407841047535627539751536107205657109999060269823798922446012884231956881529943225802891486549313473439710094490961528623226595708619069924954074774482653190892806419383647914949957502701782523399110656;
R[390]<=2560'd12828159211716870479923636824733980678479828995339403413231333377965392602570632879112481943558852024578335035761536534278655355822061708991314485877163540465962606460062375901904140239619639110929455472687041757876698122688104732467216790540563212432620839622645672402518116996369839237308095190164415941001630370393218148944503035083373772923200052696730224933287921000971965932646529420612885706852938045153806453124256538717667245975381221252126754569102660499530414517436453199138554809905876769582740490575018502410636488271292435704913782270454599318205557426966697653289280965889198909444885334658529713837361745173298732973831956543502739004007204792247465309603646862949671362362767623343971484831409777070694238217368460232424585056021066547200;
R[391]<=2560'd12804767449820017847632614557476467791618325434020036711819688469167638325137724914983293076976662464497311728235654519401837777034398591633013667660254350530768239919063457757671716985810800004144366327440469693539400421699665349840834639945845655196787229467239469540166162618236069012107851552331837040909772703651601340473212755083026028174045055572423361538680234456328242839963397171154483825757389625685747009086913031555478103499840020709327095396809769030257087901526025745790126479269398182208412735690022056777226370636553577929319310881775613937494068246836968062420615029333109953806004429565639077328331527756014844634560777292271848538860133494985702420073189384461574849248358922399611765654597898500128942336056294463391798157773109198848;
R[392]<=2560'd109016741454249125990573393814407413037758882684390258038289791453418680385164906408454536446923713893169002161254291717505139997631423025915763689967991506043798023588892491056936097975685243233743461009925274478744007477856735556372894547110631535701063348288845621038183598472641465736649126125566848738447588635296032006011307147858844380229676241548111360694394943965946090400212782310570218281787551445771184210196026849764441330743665064718356845309773400266205695462042638766257532720843767019038822014282080170732395782870904458068837185199611242101057991518295203915653425388669031782734364802530614883399056096078011039142116592494788374483062777103900949200926235825336273826470086505147434979868372724515535527453039458963122433169764768546816;
R[393]<=2560'd103026982330438231806869805262035003116429331390727072872701442756889362787260865072318596875531930564472179625991520834011346412588262461766095758435821258577116925479467254242424669104344709190232608948172328207804724808323501395909139482038531545558580527935415112293257856213453520487623678298174523786773991292739336917671829606693309044352854053164597458082920673557387107185164933459248998318172827136196159829637950993435742401637118836877534778640032275626503442708007360422232629469102330197378154007639095555105084995743272318621694462592931359635826332872068806782188361820132467684016730207815474885306031446189801633134988119083314342973781474362173768031418570005231906700368924095286720570416920991142404063929552284360804222813600902807552;
R[394]<=2560'd400877108025885365940578713010340976505649656893603798842761878908342338019578395599171169943001261154364073090857214126229440830838361839267171135134143895173650757410363776319085779921838852367009585124128112942077242709985907134021134956435485831233170104723064208088126563185675100825491036670264617463370543961490609241803105294061725325232438451150133444509899222492226438202127833524082552837204382296691626478935632809788448687478004996951140872641732469791281743417398165031951107874335393308654796891081825354507665290877591211394159536350417870896940692074666615544571325355457038380134247900578463917043965060279880524903601312268034948494864704093558579778573573653166516012627800145903485109628451121081519260560308829910928070006001369088;
R[395]<=2560'd889962143836803409860214085938336937524937632439794418615816774725056656318775198274332608440852525886236077086598050936074074419370044632552842147519377349269533053100930934812664946312670843904282324566598407020381678205532965132548808417147267835192084815490355307508287501585440057935185916805168009454441619698909114070436023297143264985422254325855561079772390854903858287706165823533928489790682217936796940739474496965258036967301095893871571832956893652905456563863887838579097198296702581224302945317388214298016538631746451592678548340248083588036655800874639366125404774276910344943930746518214877085763103578139280690267172695884663608029519129330281742223995305984;
R[396]<=2560'd3691999855047665944681715133635658367279348177316645925203759316108454721287977937375765065357731741479875239491876424521667663861264409663985883626442970852268330900051242641934934771527843969312262084645835916140317163241544066951092728012246497248530278496628883934217768894427354325889977499977859351643372280773110253590492807351095489506271765124000299013551660308479491114954784982318736856960234311954907601686225218716286055022515251901508054900500002436492473714851013415162611560703452554279420894110828016399940822402736691511092235537216396387883380552105355171427157311093082084052363764245668712311830686051000296459932802855337105978513939253176170486643556352;
R[397]<=2560'd1493041787808189526630419137355951764459199019333429443015935368902126370368334481384194930503113682293592218094954706463693390243200598200473840473763043808188974951247761901407991991418980598606605664084166742841020104185890570271520658114889047983179962053326186097296200548425492480945175684761678070910009508198118348716442233277303853387030339626162590007727950257717188996632396659238433879878760217779517010591564193697637704051713131663442031574496232157054070891104757114699605982816815042359826092213259135009509921239560311829880111396123519059227023370665638957144654205638995799347967820974734673546300481968343853137969457427286562316590674144413097151517862173027641673160814685086836053090878675823577629364588001736737635172352;
R[398]<=2560'd1493041787808189526630419137355951764459199019333429443015935368915420787724144570726446297527503732743316380166432582085205754088147784150913365327659140111593708659078172841215659883886774776425902668156280046165390279502624733830993464747575991993680916893739075628148551641743913689173545402257623407543481277382719120275136217429105135090642596103902953589422858561285121251586103023373844150957912563442542937598559943235513585704015517284861301646100177582165848367334059188351219388514647971174372852912785559771027588329980890647567169062752639597462057995442473121023944723496853427327682067181725313224570660581744142263006094323361921261289522934516955521537729425413093332190893499600336494986340304709969704921275519941719017652224;
R[399]<=2560'd54454047507783025985260790972171027364175609815406330882763344710881619338936320206682374542595760444940873714988481614793592072482787972865565433942356001302813512880390111042513568996730519186474195380961310303521862514361688259409650977636969818764173289242949196420071657831768923236053579460026710703151940728267153153840321984210533302680561306762446518157630928179122167976048276744492891480075407788217056300658459716534112776261687620246882677255440061647355094981939690728568233620403334332740020770641687606910190386924582657762019247954407854685698756506915234581252937107572799037195149462594327309247527318232130269439822177525847187742463025700491609126791902052483072;
R[400]<=2560'd862759507807732459914819944468806323091541822498361678160148720473875179169591372640270118711054116335522799055929933104777825257482763595817077514405379589594422965713550846949705214144378810702260907338636827241089128948007745669877946238543862482951241689687796920247775855192157142378430051597069072666111452155788404007556627219388847256847343604728702358579760346386722521406713792616645865461446781710003516847543751717113529280482966553755686205914893916696907659576289162632296825412938304628887111685466545221937366337532551369276503103593490808046200984651274273928963779428242484930952370486910640189330958783685543132334981913110424357603083197324722176;
R[401]<=2560'd50785961068496665862285318833381157918816222405146543552500652370625313065206815915662253840157389576511623787100448378497509971940721310108915728621989669538718723051922537189716677802487694600899029449677382583974142226021381988780750550098454563665663574162726827602924255946698104656117907762551978084500716674684859957290773508417988651372758850101492623825160274966459430752902559391084328214352635182316126022696712878571240325236389994369622094295164000403136312560381433180793863110172708951179494454915996914712538948479124733345794135865597278512721570559830685010972206477541257311206203418638120384171967983254747969242340659192760945091693511092207616;
R[402]<=2560'd418191306422039143057782542486874579629101109224944392151352007812340413620777106036532495766203927556898522360586624696936826454884478998599596606311774307678612981477121254878418924882689198249877580274322024215874057931606171899492640520084642508844321532916652329632419601499339464958888692720491031311234700079208321749252798802065819175604773797365483715003375697738535682461027957035233995718259409492164680850377824983660653022311768064802417194590004293495423122664250289641107686776039917800796391594621252981005042325041641528216527394950700393345093728542594935056680459702222480711474080110167917807640222709921502196640205060216204398362147694837760;
R[403]<=2560'd13888349039301993794746527822613710493286943598119521299381781665099834314419013698852104199200754388545497678739107913911793757783460774037928208893379529357130343673298337478018316395196330634375285990621893872540179646080753424106420697014672505967998641199719161067404506613838514805265506828882098251982926786072784907687995883869225995367644320430461801065548778175806665203258196856322322129545037509263481835850378351035354147091113831801786056820727015578902842036799036147250173955087157171031423909898164163052632018845418216349137502246201867548226336670202184149890108545892868535868930074743566559569992157937418724665395884703206014252001926316032;
R[404]<=2560'd13470981613970287946777546274048680870179544693219978897365995780840469016992491223689955797689402617172820017365990198222965796828149111871482919757932782227759396964227241540983889826529819125992779852457756249816831210504612148504074266679074675640940936864907615489330760398691342931746547812435160478735885381732704737443429898064793480204674316061817894132741935360776312543127632174195142977244977174035475254104887932135421474553436643666241226606388862818147174267721721430196611493417365524337815982706241800745830937563547451141679652825051230832955608431270736164871266434367344279372843823829942179482837962025520621302849631123451477753344338859523467793924096;
R[405]<=2560'd200922828540406531708023638636155799731906055247861143214265263602899144235869690960584990312468273432138450134900234478171217254505431413034431120707351984320590816323906398131522610393906461905316591332989494397988275198051106438361421969166706358456723698079677499762404833095480373839910348196528677748670096527088244531069299811296980349131070203331823853960910419647870216912915426945314471351177661518915209311044537963344103279586969647770997279133656939696043421819013999412719944282876299311230583878843066689845253596881946046695268403324513669790959108619477176932910709423527070396931520964628645205032390488224428099637862670397206074354565120;
R[406]<=2560'd802933073877986029794809829903275455291981564479579891214313998630976590205899010302523618630724225830425178299472034270304542302236196679386551079829287533633392229716598261063093274102580786585760331253599802816676486837952775814670956868644686606144208858679091508607347503306534800224763701116317416696486164088572140812417929325451196432087051376197852111353664135899245693176432557328114454972723203967683056064828698647313090815416019159965775736703906030157265327335308984653106132509301054888008472419937844482958360575366410132577013477540225190390757163136600657041951909120133817126148903810715898080221983090011510597167471571556581696881681579968036864;
R[407]<=2560'd841936350873139605322074738748897311010086061938602061180165296926450545129318685815930257953638342795963536461510736728375899923053680205862519440487072696252716854557095306970634889269169748651696245021783327097338764182959660289947072582144502056930645168847140859807282823398579376749828353658537777775163902907105070489216912972642449819044991522417158826784348654986557925903345192161052356915870852782036123901662098003037499650917604519561987321745452883545796345653148586289511329066896715107994942653996970626847728327926124923532916310199661972742930603117883933434193837089565637541463798349707964097042603712326937948737810225593230678551992211581617165041664;
R[408]<=2560'd84558727106507213883799924563964108508929340679810295926805267374410489302158343503925779238882858406087686080609727924217147394000910682969520538194262284016478194769056234162648664909647894470815951513675658958690432275784916180932736239132211311870047008630195409987625074926418772854040599512077000669117433600246928129840158824063045852965050869650091386844284063728901174729436601968403316003469623749823201527237797581419611977513588993651729144840971679653266456632900004382657758041412891385847123750891815655076030202038164434261597044950515775576661133254601423307265842485281585775702686938421842479589263675257666873110623855129939936258650552031662120863041431186683329087668817587279053776636648149277362818553741312;
R[409]<=2560'd84558797964279528688573979438436999816447336957011071081169898418083663619122001332653743163522442145546993792206617518320029541597480900435410689587019447680659428629987530202224754078110118777479660077897691847017924768310123430585604951172068304866228994074532415400654119250850254195409003123267756103500651174090183339259026797842570467700787056169759561367165550775297997916566880788447074160057317870474956172271870912039761518571430130993154947322422672832511035886694690495461692094194288154872079197392118520208456821209203469053692123259021005504390109521217350255093944388497381192810762793110205394353913882338709794165690135138261561713857127392167390106054320248551709293767000618131165724200840917317346095846653952;
R[410]<=2560'd331597771775338103801301767564449254427565619614151679007094689846189324020044666722814337666795324616983220019045094694719164781994775592256315503583526745633181435665379098409622494907072938522165138498397149606425090747165560187051286979103621599184814185527968348861897202131276138374622545516201652028148667008040546340415626799875892491049721109233788417815230167992214595186491044634554143224377301838991006384776065145522588405735641022269713734615661717907923581926539891988285812342806668421117598836388048099915404050002926949002946323081765875928222481187179360980278371103423431201415265033758032035967678716938075443673798628895899085289123807085476972208672350193729287515298072574495007830377979499574764301713408;
R[411]<=2560'd331521873910431869398966839258758146793226510980685404875941772773667879908344038505959572156456198945798954632102234114489879118747165966689797643815972108664282179362444285289514636231816012981540443815121201000006687676938459155914997657258013482368187634638593718065276531170890437854650961726294476459776696591333132732597652448454915132705025507380543310628927647392172434214724947572392356924904670916354904839200948376679668063390407826592544103779116494690442077377334039624341058117451360758399228403184788078871091533864415001638516267445827768447305243763454282143854909492330300886782743722674324947256854256393164605014137852016544089843869670460269890003760724909061453839982865665133679258383138994212888878514176;
R[412]<=2560'd47208209521469483066006922156132956292907315117999206838903648761181888818001820156124314677916569984432460551879544012439629021079282215503144657502739898986253746163250053902228920503499695699696628249984989843478709745754435933876100357742792649839108212859029389668910283012062973959022172706304904593618715774863454545635860631349448713125354066196548458701951279477164945653184254159597642533438261752842353764157185683887751927858493414345853640270344843258170417513421549152732566319754213466378549415474039602802906876335906922984764050320946460692687562061329005652981296435594312684105964695405185270597572940781229465081454002176;
R[413]<=2560'd336423515957514694676592972830334627781251583854633120954712829221390308448031326253513382987593393590096022240712920959244759783895891161329187414110195423380450735059401767125956196850645217017279813256794657185928081933778563450013353388428215165434188419214263106485067947836268797606029617765653996863205390346587332961625675055167250299097731919176887801650585186718822470268662620696765681387153888148290071537819560237016436983195711990096887521425443108723244212465156412409018840186882079244941891622751725856572872206087832792097548357687255710918053802533790885933021148355795906430001318766594910188345736834905747016237711360;
R[414]<=2560'd310877654655936111963866340110776870252988962677858841202348329047835081525773164313268852057665717712940947192670611006326723001336189939600066686090719677669203965902603179247932260641272710482112228427727299167315433150974884719941595383066936189041804202475661291518460500725929295721698917932119268595153118573351828647122506920173751974873204887777011165422598925770951702754608944685257388333765296837204656019852047541632424344821849069764967539749516947271929059568514127265136922328566199462178278553847877689143497863344775176039418981985270064975095257796833818644779056575051850512579163919623201922649918237393487647095688216747548034357731407426917659513179372504254457120526080654461673524044403907752713332457472;
R[415]<=2560'd330307508071932118961607986367700424643800772845225018777495099613324774121133987082848155299784281478585075085924414553926531319170398469407275405298939374572672560776468160776823315853077615096693925611149726744270189330970511263406050615664217677063490183384940429812731771850906183571357156405962848797971882368705732356965631484044565976936900988503117733260131967570554820867298003715835437443650112650270113067414939538152075065335839718665183326553216266362029764476180243485658644540211148748706586059770242956014978815439651070267119639722349662455029512111006564353524028792148191249759343284720599527122868262042652397679074822680701426061780471982379485080315020251495132231061528288554260139272377824610224823074816;
R[416]<=2560'd16071998050459114315688786864282501165077657772274693713005243883014820949941526882057136816027612695602869299714286425220131995398093613470582610047558877166971970174724115216551943161194663713388961942141701818079035970502906389590215771236112803323359471257512298036792448828221064860443484231929871643466455162987996672591317460568236441504257811192398269408713560942319409903353041673276579134677470651560177506670258679828954580942655293443660368166364503262353207179468709379111501486887605094548580845431721095672247168238495995825863736995864985046010256903837395276439050936635753854930309847867275735783242635091351997832348201533852612758808411630221862534818412804928470656362469788175302656;
R[417]<=2560'd16345290347096838832583423010815392501898857101168451397308824882146827428620176752916887510550373103707908740165257566824007232276896602549611278643507074655326724308017422375604081840849930875995539321857394396045229353097437551388564910264611407687062747709809964869408571233738422060967424897948566394700663000559354070591208918055116030652687936379730030478168307085058134259312502499110273610348119688235752237324991230269503015529793502003745745101659264351866980741202870160055784849235957302760299304952472154644818550839856255014346261698050076679657043121822386217585366046372042073150594683339954059853761960086228293593984176693388189055410590771575459455826153755869550701783365451776;
R[418]<=2560'd59872858414274134917887996376613159347614861176441213909556135099441307005238951653136895245318122529193843673040021706779645859137980032463698600502206997579100651506126037553191641058898011373031203514736876201842661167219402374861841124100984648647320509056851947281294314425847112505731177458639144282594812944320678997273140539963599420018586420965783424726418776333068766266033195115513595872976785129878936137115043114878035884349768599849066060142379677691675054850621857131340261114684087784754341684818519423368388297501015910640444666654864850588675435483521883240373532565295953530221594746669898742424754202310183023640088315925199266812167628027279722263000589684590778501228920832;
R[419]<=2560'd59872858414274134917887996376613159347614861176441213909556135099436430481702590687526449038116444880857168602675445754823650977185710191719441711553404402968391136716339302024343668506223304461963385430878821578168015523359758813178123531449519505113664432217341863525982853427905755573364572412007874639571709892324902514617078317344902871726710991928025533355131648115832805973682177739590241471279975318046207119841066078760976176326509178467025306400459701288786390391252439505727659446749816244255210795544715598546748868334968300951320127227295344779165720190021648033986554473269265864214967571699443818665870020073905976287357333293620289855206695166533987885058153512891247855742746624;
R[420]<=2560'd16071998050459114315688786864282501165077657772274693713005243883014820764945281141765842320406578973054717942106649910419172432595607506398836762085183809371125231235185131186073771523836770408103280109769513220420841682443278539861706656503252399016171317238555394771061876794942238691253626270886949940039921812526736934471007217960470382986877573542478557285543811259323027326727335923305508052285931047901357255543961161784689190929134100859749474621407949310349906690157032172538404910188909473449771715043378634252603047312207856771993953733351013510853098580839837505675103065245739197407973669941823345341960736154479680204310783439181219596000654247209371638450696646729321875616521062478512128;
R[421]<=2560'd16071998050459114315688786864282501165077657772274693713005243883014820764945280527435683359596305367503631343239905708448794749203169689577467684058839098951914913361799369748843055701269542261278804104765399975435546959816440386777338344233165811184874341801750146700345917759010055656649129325246771368039142483780544386092799182409392217796683793431368952724634955586833975931115347926970468683589336802251564707145267272808305241180631431567800775686370228655490024956754755575528303204675748352344447065908034970476921839269035571805614703209164897351120231130141936320985011515153452468170306706147215028372003493673598470502890700690974085374979561823130969757925403080307889883890624751770533888;
R[422]<=2560'd145542856500637466779511011192686848224711866683983984643117033499555184573191688545554602978920383508211220974875009745231956849071118134330649515759408934888172249457035630528694974670080119758381736391148421248863456243277193659294855630176902692150260362914540907867592790071239794660351664319960920925679377306754240779089574745013999058810117891316738095201216318191203923328427456729311330822961110882948811144588698751820886183648646974651148810710862366772092183506017620728780268470659697683276285502323059575828060015649197178100569414015256294642247247054754343242315738870113950325361149394554462947049101012783092203520;
R[423]<=2560'd542189430255173537666686639498907034953504264642844394716798749643052202035333585570241279680073581186260040910044056309812101596783202764054633192431838058102034393314055866459364330812662496340566600161157211410976973017594748787633044295264091979716605662684778578889747713385118631699469819744619705658602765818427511386817446375952367050616385083690861657450445690552179448278680972863413327485358022923204701620469763478253617098663724949154650005040003111492023009137266025651153293517192529133212338392487860900143338795733335620286402278094091042540178460606527278898940361281366722923808880148528477268120168300544;
R[424]<=2560'd2298095889994821023518975698609509503666522255464822801260920562110446064383806023305340954630224186704253909881889299075023958284747055175681640271379098919349929483382133423160723206024177040682559573563893724631447200751510276164132325723740011858260858783137818445005686564709561775676331911933143619952339309902600784323597363866075604514180919876303522667837808205591680091305423370609248920457009428052676805890020959943720740595674207556747314269498012412629565742859235243473664491881886229020004270563585039592792658822429367381430624914491320523109469081149359993117306015469910483780386207429493981708288;
R[425]<=2560'd135182367475692618321699195834733942352959747211207853694184203089600239935124591976640809728319968141196742232337766456230489186840698351583826057770218625633651201632551660194624638498257128270566283699359307953130802273151298081143946327738142564460038456570466829514017085188941248197821592256217470194764011244020200029437904101202020794782479055444256881305470917693783460741296225006183499039088266234776949326971402910237406628457168064306737796094644518006226285996610891207009226398921163992050486228349947254742222027402655462521759648217817288646922906304424103212577978809276313949659356675291087896576;
R[426]<=2560'd792410683174719618142403921016562069266002468049343401034418902823387987167004328920977190408554508563198793968545959099855777589639191708059158262344484735000249456609466385828133250581140515440190962228310087932612688501859038552843397147551670156386803987248857059541509165621632133849287375055469161315861468051164295180883135375448301335191110883514132997832910059538697916933913708676139302547177374850941012286444521919557900887550520161419887645778451533284046320485224609037337853209297860723744980286671651893803628308441664659199123807527390992501552316600242445959612154726747709449118290008613457285598031211122596043262305367473772230220517151694959706898432;
R[427]<=2560'd13470981613970233508420866657281555177522041956838837817585120754073501529818791348098189281650840292950418274060416403775919222499242430312238916909483172738930411128726891369873047926967142215942691465412841089456815099070077286837564939435662315223778821604021767908735666344470513094597255279340926332162287956470967326953058284800357632132017748832670175981930096414494537640368158348718725131635672448340516000027061360799980250157723420059445878984296923377306806513978095397033923789310451178992851798046820661253201334887294475580440346820639609714982565426978645416973112264439737892487107033728917805441989700371936185814186195968554745192778068677726368329367552;
R[428]<=2560'd269643382844131460043002966000030207080283123902662509776847888948396696354802652541803917760512822515226341965591835322086722575665868969906939372041570233681998804225943775057706310253806585715823463928567469266300837170341847539771855666579081377453006875519145811545731332485700951557919226009537560955372538085968683335378130455113847080547028931827079520196405424605765532799351246840402296810067289688822231475916491933606831174386651650195008512242656555208322260565906573525784575883390792509905831528107290509257037750410610854824409178657047694880416967666337737719340958079577852090058020710618659820029106775028132462032300954075641673100056384026455897660054847359363754761540021836711838921785344;
R[429]<=2560'd269643382844131460043002966000030207080283330209231138754104428175186588095072227297161447849651313570095332160372751562941020078143663646028273248144057947910346470742965251520584908226802695471887817063040393183802577542699764562870689156292541126021848630712100264416777569895846095797756925564761807781503869334414598641358181059093949248569667522172956679396243493357557546215773416179671123774644634935560813151122947972507567662226370815280435513868657345994233139597394808599480626457194239991522482685355018262316518053862752282640637760627469470817640248133475605213382774881129894089935293747777225368266040157230143055142915210064898526749253648270700762083368934449001852512012394929027331498442752;
R[430]<=2560'd287549388736124564811483631710969713018310329665215642316088126448179996087146943673301862095333745446546114612296804948281926091530992900564944573243546318658635876471944444183951485043709821750916568995831055483387766408933386434394080415486861557470507978663924631765324367176372312458320445058312901664185474867648684638304452425271159384890036541267785509722341247488039447474322218525725419669539175846841315716083499177506780529595436226647805335923985760071476443660272563059701312856054638673485049511560884405876644925814159776689339331743663297885680141632251419604216098396624831166214096459774074539032521427761851108198029560809433513573277797160600744767055307280741276798445647045446039890821120;
R[431]<=2560'd845238058904277106894979680903215812043988261786891851059284605293500833442464071419492430486060081575812714298691219121994109708623891866335028618582642643291843496781449798896824425410914251584485542597863047106432436613061362537803329320647200698919890385096038783805497470532319132803385806093893150114794704312209912919587775111322505842547963065275235787987029637439812511582062217748710802224810924311118937732468799283934721387941727835116592576772247427743205964912200698511368351282967505586019850295398921195767637306768880882163025620422143884421159678556443505430573219863563682699095235710232248393277055179026422322339501991038605902190558818692015214034944;
R[432]<=2560'd14811500922130502915847482749949290231794744616576855868049323002173864180226355985930687664885644589159528574400112275443094521205481237006393782470350018009214302243023691257460706076205933516236253553322936977327539905433957053904278728074551055137429672785242192322104810418163353839208303047340138546785994957040314879114051014115621075665099557316093427017774855694612814336488496091598104302945106484341362112366937922781372503703488597144412072502072676696557769155036629735849444226314646502952133842057479156695842249184805122698772473365033651769856163826645097339715742039124891737287097732597826081220722934866862935839148656686590428944124457741359800179724080623795568640;
R[433]<=2560'd13523808992836248317003575416723618493616963940239526826442972261613706096872451237251463753410753074703569888073901347384156198374218970109298669354006957698634119150014301098479482392107707330131062058531815857535057347723364682332251461031408109109895566911913669414083730986086595894489857004242213207263764587634958587537040118118778895075135414319681026172439282564477321626644963694051421842284857924308033545511655874589673303090156914215795430135607460310038501456205168697415422922456917132100142166584701656444396174147999054166191351241774910196875294685533396173237362746360784225398649303564358334988683499989586371047190018926309371833045928130858860542951424;
R[434]<=2560'd845238062052265519812723463545226155851060246264970426652685766350856631054527746102095360824341926389297223771870273459989375984412795246065280717852687321417117059782204304802513656124910527798388225993850804838511065405445058974535924700195572371219631870938385074221679474214818157684388687725605645471890247595171659563629517020226065515155662729123060197530528977397865242234440526752375265343466254359377627929315903825355085143355299254621319395415437942715351399968741829992937676922898474858277208152143191101334627863508036096329676770158939787477690955106937621734955184282450719443740728241077496410262784153061317401818751988249615461924984583040953739116544;
R[435]<=2560'd3148709106235719456584922891962705471654012201640927122861627170309996890353343090866778271942482053757967208956365808865024130678500485192746342902231511644035496747853738914027925953917060645516218783725305022444119990064358149519039996750280710646867070748183887501171850639793294340488552633023766395499171962663142995524275704071478674925124206857776635769922273497008177434898928752015743152729513841535631272548560241970016610228553698918980370016649148998480458457860490901316308269024476615849140066367959431571458671432797266805162278207023172697336584749176812541378790130958077312084079378613765530451322590217109774101554217957403736004462150066110464;
R[436]<=2560'd3148709106235719456584922891962705471654012201640927122861627170309996890346380038953307812758021087509528483335326729113042308413305887686824836021451658213002559886519874514875897706164905821897239749917560317859655554169639291964610525396054101617735068629956822093071797162978414851141052394412750453278041796877966521506690128493344799165693303935790162692483682858025008543458146494586854299608728879685077023190363353589875490830419416839546969369580054326058342505178285642787409547517758562369020149907244955376696743220437941095075349355418903533410511743279908127276055326048468703346527557897921081047538588167780968986888074524197237941097115345223680;
R[437]<=2560'd14811500922116979106857795255782587865282111016134933694843642746086981352182119752018729370255528157829775705314366535878601279590024121230826133401780304939805510706610007970683113629837000680225970245951769534309369604343434247092782571872018579447588497492920033123655326516417826033842877029320750365005660131047470180826467823480933440595832699850393385777781753174541486184063160006616644860085275619007768353205752806056777076021362184792220066777414300926712643237721374995432495790984799119406984335681178524264210634875995120155707787091958501854527796377086488002874747341885533731582121221002649479965764449248513765654321926065494829467072891822614475213511933798513639424;
R[438]<=2560'd3148756965509482246566357553836023677868551730286892365665770119963860527571112951569419897661169166596714319126496440173528437272906176281899476042367689196519579112872419531838897858037146165091865732047714400030088461275394216281887402237449102228469612174424407713251165381133503952060292452309342396530114447718044479107135105338446267002213201134108746112363232395561351856820707742260355796083611090076797039536835089688856499042989260107125922132075421577181115106732494845252656199392534787799688508821876291002056792980336353060101010342210503807365982784782683048748905209699103260468075973393364606767051290220231390642079732022010209364924373143650304;
R[439]<=2560'd196797135081121776396560308361260205244419439620552815370227687006829426090551116870897779926909895076934756412239176000716318188533719925614687090983289874189395896752859828800020735334962979557569452569014352411598495059485856213215877463047607579221789691569813512083248567856854522655384565241157676559331587204779769372499535206894584966421213936008406508014068961536058209375130908855752770290497316866672148643536798187134692195351424510382129723409675051144595402771714717676799728265626643939496432667126151346586751070393567245426513209243362429708818279556737305927132203636133028946015562796282998795845004586735941202246351887316737651545730755592192;
R[440]<=2560'd54454047507783011422259729797097033270194882714617155610913379283177909869002360116005362771992929250036090431105125287666753933946809449647894872753471683791623621027906278272440682525714654385429321432918167307422162324203753898853618032961672820064268470706113069281216850782456711487388430585837422018336114766407637604822872864808259576986182424698010513717822800035155363967234739079916366634541408864227279482077839560903302889346339938160778487158024643387788351536877604146299753770257160822721802708690725878948104067471343308994998378400966867309880560562503820866724291383895643422968973614703715724507502370435880385720144998774541937918228583328873394222413629716692992;
R[441]<=2560'd730263376568940700859625258789615749768712687965711991346677261175811729158954226168239895881274863774638020774561234630385542615154831147760018432740970275360326733515286120856698198619252633784829269122475159130506419178563416225917993890243057486367603571158105228807768895904065573675523887786808417700400229383236545702859655869682524395613164460274019422080079820682596313914915041098487506008998595051847697009534161306452021141827009977360652246848687829960175596834285381509635927511458608802770781426697988680813067082700451379013832071312691587806196223245771540459033119989825407794997750399254307497362163130921092044267143020862713484017664;
R[442]<=2560'd45809260524660112898593220507712568861870074405937356074826032238280469223436234072531722698406858741051918717045216060025340105887264435852193487873932951820849591688736750924252191645112849916267249315786691880602728258604338016909905550478741916461545386250246482640652132968716526189915061786668090522289093898146626212190225397059519936489255415853225660231195241305992741306248078362897260838988721406326803013177723093518747483404548158540616247810047170377718186795235474645237424874796083899946834421203367379039596915258805244955175683574364274217623018126463808377962248015036486468342383709378293265259365178749893819636448969901976101847040;
R[443]<=2560'd45809263085077121890888979581226871864563270901472757691595680351228265749225082063741073629744023580395871775550268981650993336254378003354241978691654443304624138883951824625483812313093294151568514309073135610387369281467670219283971098533696511311913465128346015752536983147859868764564148473406247759143544149090356823164196443128253877524095539617989281492753957121118435000502787897024779315543341714571401309387751478155307331216837112692739382899041050818105395101639834791345594648199340853767392188962853717035357598481537850174037088668130472728356110489930623215564747763119741027740811314548671763988511836881406603104592153827286167060480;
R[444]<=2560'd45809263085077121890888979581226871864563270901472757691595680357754639375096570542457361198040451633845090036594938142707926810475817488830501551293462029389434936286190828425014525948855819981737756187648050237097694952137612797439083029020667539179044726243193455026616662219448007340467466683954252654617252167239135170161074106442516195538302511626281959766971403476094192543250137641771478502237468650925245365028216294830671056011080702485074010642113381340680674032334830981647410911808791908829259617623279603373135779915204249412487198032439138435103691826154960580292540623373606367497999673031049299645613372768311937565867203529513478651904;
R[445]<=2560'd733115970444080134464653929030276989293939918398613455429644867339819748097647530281667495186866876517085167224342681094375006218187326521271771833955869193399902567587186311072706857764636638210200677115278341502068287832819503634309135838262319247390497755952754701145765196066744463730167738091948182616336894037010504117775536921198722727619110460672515519049452856220145745349720930459535464771857616208755486407426535190824639636623303610023546256693212395397652940053152558186293961004946592614993223661021325213932620821958556442500598270697742370156723352927844494094131983785805076177426840654860963926507632451512009468237279912840224330219520;
R[446]<=2560'd733127110818486259943501657891009354012037870473145889994383805000918290657889725360900188829268286001019690770150791938514331628740252630516050527976230451370889760142951602695896763602923750503015238390782061719771302782712388600426974877699841001209901578533081110389226990855996971710983706674099422864269069763860008422181604048562013769533011301930695379882793735293077183219537955887290840749315119557381907022241762487399238044303993249795893747956784919028618771894963525658815798410680357467717562591126369285339649687398244781527616470316138313521224234528341679778623481728455954871150807545912766796732195919883095260577101666507601355997184;
R[447]<=2560'd54454047507783011422259729786143093150095513178042938039359956983721643539158251693961996465407827650893396553715278557315235857398858263772153808847941932164807140347402738301989141812200293693241669450028441499794938129871519697425601545278958371531493126100416129330686152760136580920251565403182738590120386677828373408546424241340860886020284409803429415745894552840678700983038836121803392267491106840247476339952691974012169976599784862661302039530543376826243465613652864757311780759354121689770626169902136195116151974643648707423030833687148529349592661085475097867498540265924646644270874966618621370910101929478495622794787758573179033943628374829849418803432839127760896;
R[448]<=2560'd6613030781228709494345677548871862230391902859855834286189875385946889970147418863843378937639127808320203918191267461212734660798972334263574329132439242458557321985092634264192249172378434196639715274698269277854234574133727049888866744375449994196704090442916061743414279016760767639908978961737481326435522560678761227776614366352108848964613002883370448598529478436466239018254640083276022201769876210222880721911618790379501668600570368676068409539558002257905640313715245227741590638214347747779976947064752649116892277537434578427726868253377283024616785456634033647606824960;
R[449]<=2560'd3742053650892133432367999773538322459225928823527575869347258443714776254479140165467924450143929014376701328044210206508077474988048249115724382795449561804101395202715992313387002230914292414059919513091074291001085655127805431501636336560296045569746324243978906254446466591849730349755870956762936177892782851939643713181740966787046383467430613283629097749174178949040940972825632789533260831929958383570589789904893954262698957215539182337793190391741090833398321104932837941439383124864410410169059865552096602981336053283190008904738843449629376937574265244739303342293716693242787314983121133868443337025544869584683842845704958839918288197694183624029882344176950644163128895865880576;
R[450]<=2560'd63614912065166268350255996150151481806840789999968789778903393543151196326145382812954715652446793244403922576744547165432261570959077952571638153982433111289420534943709725973530190478632002348363667765628640519045622188548733550467879397419270917704869042279905901497514177990680038142438357617337825038059022165288544133831191571040662143605103607622073471930237432906188686528532652635376502133718381446644727642616911834846640083471404715357699185518184895695169730852456060740262213354288703994740980366281772884771041343431643898979817989455582673551300690651390214467256515866789884599870046539273261241666652112102117637283520267890012514113754397755242168196244403003542176238139342848;
R[451]<=2560'd20457887961217337850711660704216106603052382081189284396601488260045146429118212912885467223834120398278215254834494797878096153042887635028461531582375768235145639305911252688342071658403807887864460823865411988760323089076260661199054717223543417949865103470034786887653762198635835677854647570532545651722355004533373752959608405315144793750248255861290040655857452661670504719406408628512230906810771210419725412796816579695424767133605630967580667887303060649470069817518394244695633760844047127831435817281359916125720906586493578435155214729216;
R[452]<=2560'd5237139422742051275910067458563335677476390497642818255658004925335665628343701443101850267757763208003488906016656851207957351656083537981232274796287226688644920531267598182178853338997359545296310920265094654649833710421359191951343567903744436229332548880177747842486083576618505431030836708604923242698658960306178629654578754968424101961188604194627382498277180632776202857356547201573318305034671885219769939003875370099402213834348218326234971600030181838130790800007987849114825472964479550286473906940374225301134698173133062583821548585484288;
R[453]<=2560'd5216761448334513262235020346059532842953857036693831205524260891982235708253796029917131147504958483837639445957739536261910902336491977752584629942583919580782420142466788902460823397436657399954371592590300465083947279102379702362060990670002460583038443839035913057287457313757631196311001126112267844073065954881194546357058028711262818899518847523958911566563201580163467480419324753689252601819321006458995052945814473170221082364693783027833926008435461719299681459485641530102318830755841575872063155342675833891408287281757020986573133984038912;
R[454]<=2560'd5398484928428591658019859315901837254618609460557424960467397595046241867785799819536236261791255857160682828825132898019097135628719052624908726699150013771315308705254311093661850922121851123725498404611126069617840386482507754816797494876919632356427745061425565758646124548671477452321278862327560523404452788008025977509203457669108034616296976370068951527211100740003651069173991535648229865337948932657183670902573147483919328652386308875271194386945472031734122083819108400229912585720301554190645419736908403731720845132237547998731363836189593440446578688;
R[455]<=2560'd1519538322892631660972446247418949219296324005660624011595222751201040299131284998613764783832311835811999056684859548384956917558180437956864974463709618965461634658861980317112507147254549864374039163530415261674945667518581402894270108644200067468890728103521908246228279066125851830914483933740306494475993677541626231874788776218921387681002544624195771852882182800933841321029244363237022221245935281789525239476747159167314675535749548420193024960067143414092081706653914066406732881759537968025847962808305794624779588126810668834771327495557348248582291300001807794700288;
R[456]<=2560'd5660807748171842889009917883595394469475052619920480256643646453270818409482158895416280567894408857367596058491783797983844982474676383739238657903329025183868226914645658194951307391548130659026099072512557787083557891156602318211275084377723144683922830171766050915247007733710267800324575872075878754322866446652638550264105884047004347919772489998410199527645356931176221833249657641478650058701328979042683180822610328327848812407694795436119432985926452630212480064293949232598460562040392617062227834803941387206382992302966499906565623879124525446343456347652096;
R[457]<=2560'd5490282102021674462536968404635136178847218716396725159413405606031980972945914678736740169760034912030830659299187467384220946240814570715391257490816324287608305937025179421088364635214578296428037761966142146143073735204106320559737588779061850394222976611973857961752115422857106061546141221704415068022311392212012582424011107790576877171450008099281930411781277418460306188702997392994166403526587343394494528844531030463504442031938352453641324069947746706459346207782334520956241397098426178335658237397905081340382679588747039531102501425272911298560;
R[458]<=2560'd2250297766757528060363378293585466094909643757097628584211675966172632078907267056294086240674665098970649373303513462755685013357007775537918393306611932825408415628470160305351803125831300962704603533713495202526872855605106208030681511048955926840676736176545671896108157136372877329031250631075239401076619354906914337843634079002429616026912533061368350411797158040366140162477045348324533244592219306643816665325778936019821221051122011380319768027747496477190900088338993274945612594431847987885120756999385317254336771073608852169406984015919770661094668954916388769339961131540354022900891779849203318125141950464;
R[459]<=2560'd38255062034877977026177430990952923613463943876989646440678099775994602510038551423119701779575718676984194365267817533231549432406789619084650439829914154418713400444724739365331524259382491775918665237315064254109312406660655299032966018720680329248427685900396388997026733809617123856947905221947181276808947331306338526751243739140965932059961702094349265754481316214940765147301843203330178256584602295420210816539586041976615346818006031354450972888879652532529996288959933067391119494710394486956753332543854836832638533117484583340186988903897721340107336921758517010309501944496897188683752808854560907752430895104;
R[460]<=2560'd578194155599816621627484493316547994268548466535886801176320088913447313106701098213049063879180391798402051474652513085989015020705677592789148856756327054470737723348809567937812926546815316185587961904667592583608689740667260304054630754335686386736081823942911032109910206852139738960650753394623378324808600484502488015895437664788908203684980568105243887923890418114632410152978585623156162825315256450325623104488023230167779089805249812089557498919393664942994641327640278121381573442343398027983207981344502842639834776033688365284474122768354816888916412097899281211652931155056804375145486278614167519469733150720;
R[461]<=2560'd17892249913945973697835124540432957712749807493348620904754986542039218993891706609560285426472804379965466008021994293174202941615430272135291187402319850069655139320871501257572324637687591284113044777748162693504483476077720032294002383164913104444002110515540030781087076557176158583325438210528444172106844431720395360109638612474623555729459854848788837252018018100061281023378716907909091717425697387304828755326728416684675605852704428203494889965224677210388369505122202034206744475963664444534881851550403341878981721253189082045628407263026993316172811172319494453604631096388010351481352573838490384612892170256384;
R[462]<=2560'd156692734094860193899222757338943175120748314120155527613847053562246184551250611169549460061154468721401509664083974031162840689360289044304193143953849793477964812166946265323158620707921666761939354103983836313814480250733172709496247687761281139165835891455481906688131749916275057612042452466976390699197810546547891694736316711534726912235137481831300730920962225446950878735036357129878551472595263453021061026668532209781692593358490611580222001201185321325021217550427808815144318208560368202029632107220880543637177616657404417235384696070951962281879358936168732777346075626845475257253011596683019676844306677628928;
R[463]<=2560'd60667907776991146471202347000463109132192141788440003476571522293024134674821788543153332786714036411597384955107640624667015965497163518457753120166687084966038891051036030899525518925008266059648539075454935686599784276954881293741098629449712440606109117237868112921716547602933654239733337464411436182741283062860674452579045255278728084468649995446826734620340834657252203304599971784893025529029566865432481841898107217155813049042396272662342574995515405286127559271476642985512589485940586399609544804393683315937101521346965113018688554648404667332415268500360033998370981592069995234784397718881892862317494281257301175934944308155564892071439317553814412331582345941940272365568;
R[464]<=2560'd24630265345133851684592839489774321983011982656112682665468339468736876812293776615626336789837756771381025545554249238817396088481162607203904074540374710073187058030365424918776072078960827719730111103066613019197237055434859360553938933599812973275675194277508905792302237133514130005620068615063513743242625082776242047098868497762964845721084061956342699458428489195231726181927950808839655440687527847444944435084549397079421367059992050711959963668029887855660723824271575163886775884396181173354924770079581644152060909518402816675368971414843847200141886745871426022597767704252359846713797350933562741702378688913474523239589281745969072329504704821151767510049944404519843506435439266284176401187533772715342591808077507142339005182594886308724736;
R[465]<=2560'd1715054636911677635422294878265538158479251037731161574604089646357207061648773964739148946377290719056712207783378194615087604282713267166306510433937976679728933964081744934245786436302452855399267922755402903509021479320002053230906432788496913884452536643081508813220089208832929207185119145772670991066577295069252236224846353071219263697892661391303924579547270048003276510222067136063783205666736062510859104071438372273986590905084263392618387288025493973988087922676971162274458519687246574744613022301430884707806780592745698472137708387031969021062232140515302738256580057475272650285803145943081308726820846868635127252255490298570420416699983602736041145438654898944252877191698187220821285149137534237677319518561341313182589896842816340923420508160;
R[466]<=2560'd6437614734768992877050454372098012541450403863866512650673381132833836909457710653322613378993222334465712912365466799916740955700903491030805658781416604528758135584696801772397016732875570804966201064936314343498618605615823955162552917128122509172483867787234332892294528956917968342440134036047555551875643096825340721698373233350735690569465173368363444510743648483807714358229529591013234325769256955136139937390835380075062394883213752700205571863459328537400660072388661241287979538167202502253891769134154486337948788438490454927118435073347517425556159387237854165943943584257776067359600108290686064107382871065599524528943089971144684396923326144140828153628555737670344479944974455702991219775195882392864345077785461833285621484137111093248;
R[467]<=2560'd6414034110726200009033546941810886386503025053126107906715922020755233929037325479446792272561786227410607590692534063418427631467251867074652040237666576814569932094398112335004343581006768566745830930315030583054887973788485239888976939000657692430289478623605239757295111174100908735433944002302293880570511069577237083529830457103943351556094438316863156455067219421567228713988335319848189767166649863439483498105136083108411887273869651738450293734833846069521029942046778775480265369584901901925897087846259965644765076804737272444422799096115682195261174671014092424259237369285567342119434210466523015486304295415229178656024736616039051176167462601771298431388253131035735674526119389735446371907416429564166359207847394609814372716841097232384;
R[468]<=2560'd6116899231352010588692912491002517341701099968160183252840080180177279449304537884595888951017519723646296354700704913414084395890029279507549927613850179013232576632648908906998869401600065813521492912413895295269913092727682544552863974753057284840451419829278963747589457155721839283898756522407557331196429983396511036164907962668438981329680838126433939947137004054299425546383690506800483309481694913748680000257544476650119304716924293921065040968801108820345228473270722031583437665467040789389720986408229978270343758293839956545331578777228912443949036512109092911518616962456932498232133954354488397388165144419112648965942153369006645857708184891332534114342716178547260628090587074352404137636995961414971441583222632960859507697647616;
R[469]<=2560'd24630290400333921931617441007146556724093598996443819707875036586452786944245089467559389312042984220644044664278154460785157655936202529997837358099552723706667216399826050990129857442895023165563629998371285947587932997544452787518471491450571071646732560609889777508141004543032422877358859967176415205670768369549574745546759910442249861797389816987940576082481623383700931805563689991645705249082432531924346346911923201555974196640867190386597079705271790245433942868552829517181735195372102627984918489897392234868786118493977311989213447243371722434491695121789177305332708722824255612531894163818807150535710299516893950958192410888893053893006988635057529363590466045099033644807953335106811245185514063637901684706954475762059942894789406935220224;
R[470]<=2560'd6725704456905100107436900048333174295956510044095245913092935644490609821169984166730443696721226607314087231341373825808163820981348237059640632169127380006585638223782849229547380632617666341091297725076324192180052336512473551727834603751385132263963903830927989680207445848450350481085788942349654412957584513067072602493314876576519717483175538419370688723570464671163377520069712141440789454535441605642907366891232111629722049754136025920923623039896843156546804519556214811202853774952204499044338488344041904874894309714977962044832070254821684730526042111381258811994215263807617649748931421511793599945805421065194471812682152282803657868640255255048313793542600949505342901734989777517449547047673999563826963452960140237243510624209408143636037632;
R[471]<=2560'd440775767288133425994122028163678371364413113796015048124354045077851382237722743186369036681088688340366260901455331400850778455819776507138528380803825553741459834298741631413872845597456129419568202523364049556906705431596386572475208895603729247323028325507855042048390460261992831662491892015942478012714006083923072668711414492951424761946911657049320727744825805003683990200509123636364314438524875472297113618101999280794051147647392168650640564197002245630790573134205710505464650598173737929150741689414668458869204246458743227704812990451218979426807447021059649361016875786945845043321459351185388692484143766403995220212235739955562980465264384363411338075036348057692920582515313157986089411775875023493207364226509239520813317203414505646824538243072;
R[472]<=2560'd1918256132487621974193347895151314843459405821322660565899360273056784924517511088016561893061021147572716138203353921277904629118532150107389287887027297523088344172692926464883900265426508337945714580423564174061471447844190756904388541075193532632683029700448582628715493699051368240506317064656454454350442590178225433687267033162458867969160774279165254602886044336158483431400162907587820894621706663014942150394744042181029264407019298386670032057593326187897854244832760115836963258610666964704805549506477670881547210008737217161778491380041625789855988605143895785473159356288947371824546164985284153613131548979340230941700457764762602469670905361652887083864260013117466970378721807205720625742396402500058442635535533335106998825172390103619284110996930560;
R[473]<=2560'd59571724885910220160013548916082617318737527699823358414219598071889496175694824584486939478462670779234645508087110321805507538873878766369989439569198156512526757456959807955997459484895445504016006057667148534895339505038231842007500862490508206355685973976085634445805990383526156961070298230349612156211291431170248355649325163574410033298336524897161135897859679336171127365160357877920948925605452243787899907579682019343769457692910941027262803471478153510079070490958451451810618912328753824349501502785432142968313266861175725355887455764108145755137998111381239587760893344452642660621406241964796402411381312418525961459636414924173336451950052097016814377254845012779171347691077791994868095499901032289648187793365596227668689115942431569017638426691764224;
R[474]<=2560'd59459328672721287006973309852862471023149810363886454379565684593635507698543432729841994612555561869509104972700598772578688470190405595195284230533708124695341403555769418183450005993743298969360093301896839802070376769147870507781459049902910988753223466901112219454381416911382111763456480434685321957262736505989535384726812653290136372377438075192795541919774519653629979250746805543873040994112673662315696524567290397553956874809729787974649214418827847638305228768254416986930608770050708587037651744516085352740576151508477603754554096696841090237534664700673097567199276533123929856943991841367598401925372726369652013028968248646479477379818534486963058866040822693118696320339858813779511153211358652903636105275254279221380822597319209722165983723007246336;
R[475]<=2560'd59465940316376669995299468068298596700190956245367989826207244611483704768514375491316762861887787918220560611252636690886127377334695404629887871741498007373453442570544406768228742823682652491534178129580193400804038525294315410856829095487140970205845265790640969865902642598025174019397062724492415442192708673837771232843888907692185775669429371105832481330424332491164642761196124107800337008944026662517757261064222612163151871928421541057527111858039791083115039531569372149768072438027901071395823116123897587973488659506198636344837800228688434860226762104312480244814767239536128041381746386801273348330427323509893363879862072845196676502657182176821335096505305855358655409032504892278465415181374157029762473395175718184050202306964629786841874415273115648;
R[476]<=2560'd59465940316797026500361049184805033395877581029460197483811053876762743697326421862718406040384442648857655488147782153934191911742901737272612351006608976684302730525163421680789441596328505296464883432826534058029218156791449981837642933205120399379822286275220301859034879673872352103513238572524000455497477499511935276792833138718125334840759954189731141886847952980846992181346698992880278118503468223496804008562770620948053335371612175271039007648777210257330798735497010115618128632093309561136045544027922645221930107327099870641827728492792052948782650043506677191703403640924374476578149654431451575868628617306434232727556228830709403211518901921074918869885699893239616168485519042917789647817562270360791842841220691157163188164145100803657692521741418496;
R[477]<=2560'd7052513162176988490277952070353265252879260512207169097889679421607081811548535214358234060440298694150441374056364309242659718578059297926831136661898702340503093247917063057007253787460953830734586994406687748883831798322389646048995762832787905149008883978423527681301208688713540488763977535954422819614350003811266875075459771159949390147757124512468053971620755509570541148566092611319664299004061614510417293054545336017363728907508982136914052850521075159872977182577879409221794942026636470755029472765009959160145883305982750330134597845193913047515706975869333491425618464414039110605706107411380664763400731513416133209147702573469691881352088728595171408655281494885773408625431436940950739850888558530445955584620811078778994880208253671236137501336080;
R[478]<=2560'd27548459183624633824190032542395180272364721256983231403337180728595118654465986728926427866374383047584223445444697526888289541200313659799140353096725545957508657394722554852030326003058108124151706077272870734204812426356344387624135459026824924105593909747830087190433896550555756788255105245231187149641896999948274677982054736148912810132572970107513539197697589332897203298209708085905168132619833985093111767383935817063382088710711140096121082612332345138657777101848701735806258987368881778193097075107710598038169993850003202198206136038344665885082079229972231943731631291929808606286515315373926298629205260088971939697517643294066229259125177843641576234421829754885446669287186126175465119490988995000254827450774799424989706676880669931122418857011;
R[479]<=2560'd59571285724758533885579757649699876520710639178279911664822497227327025832116481664776412656440048766755748121333071609499013298611007842233260442066271742993528641451653458582339006193868318219393197362052252481366887087652043593076861487645186316323342142320278552204881183175945402841703826313078600041816934660313014947711579911029986736156276993243839835392731556029354372089127681575112036292983651807390292637006218260502708856995517606484115189811681524123968782578934146940402755873161584812836870455563936848547240621377041383844580579904085078210227099438544085092599728038695687567486590054190256177932086705189855277451857295521170889896128984040558614248553146847896892100870022554539898284366930246943889666324145842127047839390112636972241283693796135168;
G[0]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496925171969057735033576824097598527785085168107277894831459066049712703896700389723584085603123985382312747032700348759204055392658519515229479066063683907478940621675446335499808634277658221467868366515898746321489526821436448892255234809771423692784338485709772541257076253027811387434301350638550706041630006625795290237392112172169576127108230397325819288199629445391225648884147093433265605986003367626965419536710250218152876774111707016774453848881614230668348562743377910263259548821187040338890302397901142705369758211051793;
G[1]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495885461657362351616942036405055437279889255336241864930055677314763570635458205460184561168312520156065598085578249936891055439719644307377843714653052538577238992161495635718356023918652072140449425214836217326681169233260179695441785720782357967849083623124172994134169194449004694799156564575237554956710998632650193559704098691081187344565085469517502692623892716423545311837400316086299168328558858480524127677460733402436907697755660067445968265274833241942808996787320990971207470182632938529830568454848362249792833255969041;
G[2]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495820479762882398559865912591538877406035824982230441511140989020827003877267741823680994220707377504979258509145243480211848514957438343362174504069686286684287087628569789063096980278065220625429911958738540217069392911932024032125534843934686796045393786140092152894097634177089132858878168719236652613450328411617905812052451970550171320323050384150441000198291779612154739007152919791708171024672790767976023290138649831773079193021441232896799127071525401227622309808810175823632077653727579802877913693746488661453081647583505;
G[3]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256726886656705387690838569640404804394626512985613087085960452164785960795291266319037962900116132588746050923464576825700744542036273482094243137271001010089245241820453418220997674569053607256181953753285570649572828097942504885970199450666676683975310783238291934575770465838185639335359281671756863032553981619559000483819473308010066557841226250002629058919028782902281420294913984258058312856291270601534375372507601463919685131983536837093847640709794298025258153684301057787653311033492737303665729225868530351418688409183162564787376401;
G[4]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256726886656705387690838569640420194963281239716087637041200627760103781157626234004806148409984126522044126952283568265301873440184812202346569955815731691494918970356662483163400759294258229057714293356378539646479793181016196327703169990897127168260792598417911843609369873714859998689164439005213811376889946501104323485125085755934693831842693215633228477532296503569499133214681634548287116594591274422452172970673755502351720666788058483960182828434134651724244427220886870000839484185519616381088687239017345664915448118739697490978738449;
G[5]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495820479762882398806118766760188213488882907009426975330970778124830502226705311902217392435893665946331253446190595833678970912370688344728648091941833772057052841937091872099113891255436085123824248517206272948131656443452209881379967151994189788881622867753003753715737666487200678329162273607104951110109256884055796026167656297860116747897392188645869519721427350813764064918483830722705529918771947583778851179621536172255758268926033782435710003157923575238516382618512471159016192401793462295974159028330529103380258190594321;
G[6]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495885461657363360268696530396299207188186238172881597180641662343106683607128635195158635697312025023809598136801353534241117579032189092335795411645343863927481433242331619788403346597894500368782879405603530663416042926441487009908669585397200280314324125140578532406810380530514160179210812785471943337327355083250348880507740642580512601583095817449562936549120150996437436242766034758473034544408255381911978823492833444076955216323434117915629489310930414194381740647038770559276759749257626450864458660625343720038146611679505;
G[7]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232174775508864414498583591238394676864329801250749821657960681663053792874854331674239364769347564989278121697808723623247414884307259839149748138519185562796709650272958305193381230690867545617997430837546165766691846433380862908816443447627273175498082666424595776097119707838646635500041869234534408306705228390332475736263432494583630298298538626969906645598807346954182475990105269900851890990688777414388928458460528446606840442134755814723535440110016148220251049841341839590052412566911031089664518527962264259108564621149170708234215457662422001700097288961478191682918284700533108033614217509296880351041546618999898250351191830033404194;
G[8]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824479185114775756264140920112177946826528997419765327024832409990686240335086425151017697486436881360672773801842456451597907402859781510036368043915875205791845801045224586715812989092781906160010313088204609119718955690084657501611537069657454038552830705552216803840850533031384886277818278787849814812453705865727468658060876631490742143539785929006209689167098589919961131946873299293168109032963488613832920560280378433068839632507820262837309113960058357706133329521208480495528382018724083952579453694336253944955742761656586513;
G[9]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496860190074577781962072055128020061979153237400715533274288478437115035947630506740662372593898067522099442182006598829395905702486904276181033664979058753280946664190140600264144499797915722566165997333415784777043111961461108575472954733554261363729712354954164174580819788697740893184708697648521354346113524763382285291670343930633408378578612811824072410798626240074239810779614894274798037888424558757717278815628390727941030307961549382643688230608148435171119536611385154867030468203613840627906109342847369558189729121374481;
G[10]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165752099751766101640786769962842950346001115369995052370117765347295950928206182138885618529781207238163983522805609939357283967308935513766291572919747014356350704958805121167926797383742231445870559655171328841302133082994700264278280462662192838272075849193270154071410341381005210754296977744290275270995796637396952631724874897544220266798713426312157572017468888739914133943713430846458797812481258805823655600713267878194188855223461028719300907644453800617421399636501449375925798581608545448092774243702065804429557745907424891153;
G[11]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165752099816747996121748232540606586457763739814874628963720449047397930673645693713060477132288873458851549425038699749094357512771993754841550221498267294618734162375515463974617730259194936983063380868959448406592228731475827698195346332880565255913785640189924274968730226190772802693202267667176822956123053195499858106394703048475881099351269328303312154934921902463886363392576328864416440824174595450011264996453166789351197115675943192246196866226785461423663427362358862781577610951253047085724100565242815590735491807764372660753;
G[12]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496925171969058743669940763248319605247811647831208998478245048954304944774812336908191093642114928597947762282723841945006852363762401016934149844366208162244397587490307694224896533326661830146614344443050609899904529197636303155082763269419809784598827211875078839026117090063850319572270775276472159067826121516177835579796049282368171278180425764857377030610283024550702824830761753949502475907358273060331460062017099032329546200063987517975813646162735403211290386129021326238513380694599920218899159955533523468744566517146129;
G[13]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496925171969058743669940763248319605247811647038631921939535921258113103399082276035033175254302574097306998481543209594715726453015284369938152363888381485617531031747758616690112506485080849871329884441080199680636875860095409960354609757679866521061560496663917682074739390395854368910010024537115686564855836042824324352632085895347116883435133077556432211716711890696114657549021387506309545433509961236441648819976422513834514797650878953327558938899849194637187537303145740393065013223109490646349410370802757617223278466834961;
G[14]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727148381052448431195533254752820664014040582327444120566723142423263118500510035428475023267948820970722888799175270115820619338529905994308520179963183020310180787108877809683007715897640323485781188181656250109405573347309540194513398033450429042808355744510464193492942052038258109108455177871166449223389255281080447366700160502169911411161773027632272196429401625334243109557002966062167722554201105742867170297308022136687988886684846431670648505216143576380678631505191261147420634866045278103192495851632293100149303123009306526622225;
G[15]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460499385428544099517477423912863812697892456033388195120701513307999921234819540801856518882708811584204518243440689353744255171077952232898711232252945866510976987722063786812391367579142184571658788883753850855331041295810952665052543579831758419299263812291705061779049163698384053016224901615473728968019293265833077973010066710222313317817166305663410455828093631270919359177042570328046642588827601400958375106918334951906898595415995314424010781747408802253234804759498634328072151690975491412942927558223461424215362915807540817255099184328889274571460083260610879591383057955394518880134989964795952854896127601885075384791716204737231284443188875947638191349296670315881327756579099976209;
G[16]<=2560'd57773361470875804093833019566109674433695879417384223129608387403904402167250072637131979281911674448251581307236049970217993113520392092419472139540270357944122757113418820042135829294691517870570749300734767382744626488491777737536128148077755423536549651649782530533872630290384839686995866474746025453236905989775139621028806743450100933830312605902440972457822481872386172213131051713486456915969643903323961612588817025473855540583788159869984360660624870260581637277244282038226747660906391688159889165140051682871927764419536164447759634334870074950522544212552938198520530110500268695368886692961196390277476760469828313834039092403769145736761052901152951483646185812064761543797291106027735165304277436884655729148261132361475230091804974303192798411823915554;
G[17]<=2560'd57773361470875804093833019566109674433695879417384223129608387403904402167250072637131979281911674448251581307236049970217993113561902796670891146474083859820929647618772269115388313439615823221975419955944216016650585033401614194353125674989006753564381396031016308298716779700295703679500700976605838151877239685530420852926696169524400842333304543368084051305730376503645337498878820038491537959712558842238699921721976640734809033265835556195553419076933894481711648579441374738998766782663001023641115086324034735500341617617205367453917696533720749768509951064124072539492224902547398107791096452529077852150340811597580651342272739066681310652059339773569332113931804234353711011642717462285972996180062999105376826696120586868295671097138261404053427406961254946;
G[18]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085625552810549758839157686887192360015491853557651277330748104484302423664279556299905852019446416191810018355786979441072188829115311002917149362909851742472052929785152139006889259540650455088369330148547988560186530171027156553674747488575126707458967617234550212269992491986739733661067668058036416603709194961922489111354052819532385178583556984773629414806620404397006949689063891365721008552914493814068663801978845138365429046420517091187096705546896235074699788892843241781506913491699562380285618047124191606248605591485231664362787006934088737748288173785749740168574303926587142214111969830710153966188224359033858699930807575409006616386700714530;
G[19]<=2560'd59571753941400006215303823886749080183769045374841949891406173018625100446153867436854295960766780898685394711409067000301951138731849584122492530585391867031803119572913471766899532298840111389689226517124398200723414578740156212415759534376212567114273561688044199701202385905430144646443193796663847656849702981783053598854030390287601970870710499637838316274395999258316145507335996046742967312960055186519337541123898484065440457752522993729562037675546633654336725655479461066160046878813526609323658930134355558758866854938911646550543605007033650385402147980498429394172063423791216185821640460708777336745665846910527003330303291637644903474029648072921431773902018377111382081045427556284202092459194576000483111000011683461222653610180979370440799707283460370;
G[20]<=2560'd59571753941400006215303823886750415393128849802575100091670664018299990268994817805160564504158454275751080196444786205875766185985070833675799610507736463523651693118080352080271112120203711693751448024068793232936698057988978925603266284134506627048994196881821938626944893648157220247390839218478907182147065315337570840073941977051302332673817570110471934852685022250359055310692698345379510387771878492474022893039543983900814620684605813915958166129802285117512771533747150937659549436849436468487804547120718716017997180381126065922558081845499207117569298372260297895872591289214753409575537227109984193851137505920070301527399118343818392081528546433359808549950238525857819381598521896172656479675682443807852383826773148217828953759725248097406822403197243666;
G[21]<=2560'd57773388810864421437930531091114993515029669712413163117307995960202087713925947334107454179807402365928693577530566870122788559589242283487533487565738670107163762852042262104702100212243712423793892887281944815269082035043932591322461618076972439855147251437940225701575486993684735127369902047898115163710815434945552165609070348916392793844746966427403106676307998707516516024966495782605320629673856638571953796587219014740757375599196234353820735090333481256813182301743573008411453892970942972963908043186565769404360315222500307985846523148536328016739753329605078958826463789782426168487996694081738877802777038065447674753553213460601633729638676342195192961421322178600164545649364680582665311312750595430294642342629311854948169712054975829408117480736563746;
G[22]<=2560'd84855037739454993595159871597420124053919749070307207440273862488030192032212558413749210696905526655134379140441401731810246931774570251068240566710100896357759619930115459236647146989955767563035482776101039070529497731319759295847732994793395185194520008397464116819651354300578739534910213143935457022733633870639634601442055786309642875524886690755122044680094501693754267159500297314091930905011619451322914261047218020987990115659831389841355587651022773229533376099462041761134654321177672244669739769954215189673762591054469887324133509373330120671715320044156017868387643696575394442452916531770215080461310406798148710783645197151113221814638773449062869817111535808615403643858762978149602260263860409449864442476250453121906632222408032474849032393191465506;
G[23]<=2560'd84861649375964315973845885099264100136387801537513608548830186779299941401213838028006693028521728066952732277283717555851361467363909521179296184455927202482001987750497632315579928703118046611367538394692936803167299286428805606412658034701768743509314817590660924812224508407579536734776619211640236769979676998251562995202363574953005908729647980011515448060601399645642359458400124370790060710406651183845025981317767160321277582181453683371820543257341946458266591025846962527216951817767964113066560941004345788104127111549566591979747407523366798148974751320732712117642494983319304844752574741030797035481266680871101640268099812630170204929232326187672096792478223549668912664308143559077376551928945226172843895610333255526866607338085989022354895218269102626;
G[24]<=2560'd57773800423978826422008855176583123029277642765628285803201997566742748536679599198696973622106724829573889808031343835210624691112881081946153909559303887450973857100125453180148253299953714414097598507500294136557970380575469219513589418965649349858373190334820032812994859638980011515400011790318492188673083021888523781935872932284095880926471488320210078903155786556919851978122509421948854253108485449872715265251877329411323900401549679906635839605653735100236338475586066496342902255509003592073608070773817473146293722316127612917724205510636958216003006840623823674791750896939652148540243122395472308112499432603146343286418397436244511692694870125014424622689543047222304831010334641178633632153930014919363111204780600814695872802207421825094822847347565073;
G[25]<=2560'd86660014513223962792591522700344256656394165043566295334803139317412879706684667599858316908390012711808695590204706273281849749653704577103150234771230295437487456415111005215582377716285036997971729521655269959104895697520761295826603887312639993012247370159909956635151139085638832988557267321700436006179170209875981370833836602055527302266316599222840538486466300351843249809430058180607798096494616475867909772606827100514831964197184459933428889413114589280782888579798570999388814604548822033486631586190444310771638085185353982190497311172510527519998300552400962132437263779713097701544468750720520229458678818554532486736509316397430854306484932683337122853721923093159118019104673313718257537442470293835171829972846065434507551694202925494223314402144297505;
G[26]<=2560'd86660040339904447088341606940214871905057057788614051303714740170003409999004904548831534089820594493104659516864472504236929727330933463854983911684658439985754458796364559798969202574183289589357352392494493857816283282416832763272056726441079477312579557217452365686733395302623232897266941826687497822742593213165737500646486315658185382546184816698369803621128904908089789625610709444128705357996941756739383423747633121650388834094131673002518425449625073611147444280912029021025574829990306943542762510433838041930192634908687019392018106150361972585946698235718653516797411079687220164598646597358068292180948376156492133292569001462412445456219189454061265903245499529969661992607086357749446333194446933520870076840170604112392314206821047321405445801151439394;
G[27]<=2560'd86547644233906531695676106026161156479019208583566578239607352809486450216677615669516001570929543478177497901335076358174579187033260228160700169875188466113270107718212700105706625402079807133056700085445826897380974896620496467689823920064956900282532753057224835840687679776725543177713180534190585069232929923390163631021110464527397841792399040157021861302872076047230047329286133086823417158172256739972565890398770091725267703623355722541056133575462143959473312368451958068811119873578932523811603733505257039285898612448659298887274055764402361329228040492315085723967004304448666125833148496558280410099123211403822766100588887209380813989806941507509354190164845584450446845413159280419685652408381748467698641165369492874647102975551125882403184201282232866;
G[28]<=2560'd84854652053934553614824225744068398425576138286243924469359133910444881964043880193450730255912619995779529260226955235517058170709580779285044604250844259452139016929293360138414377969491272466231761764816328315653418620396174934592391654258862803586949879910372262027180037630616695497354326007694139411600314431491895677259171081897395421124119861430308459571171303817218337685474351649536545589222076796077767732146512921911998992560178609699942637148366948865566650807818831733112213802307554308859450844532503532434914574426150779348266450917564987891725964460805833766363786601695904506686177792805122687994885806342995595625548392149602303626145658448838271187680760123565779414086248391245065221971233434264110910762520356119361403581741477455645674775234355745;
G[29]<=2560'd86547203465285291722476897711523170322215662470489136199964365425258687618796678191890454241767842482254485900696087950633195676139425020183363796822585646957753994772561559322601017896453552951565056846357102701123343251697872808618949524291139285516304125834556986294941525794936939967933019849508836602219909593205812379781483528549500321976714782114344488452127648671166613301273689743610271155665938216156996942764577587117420717520379293383819629297856384922706141369936854336915652988724991918979841989761514408217020792420669820591546328078041871726725600817775990299042072179625444115601893932123158799431370802281554760383850181616604042407416453832512607223817843921184206762501101149985922119732926462649201790461988077059251509393662903090478818928292405793;
G[30]<=2560'd86660040339930616723249281478364409469494149684169156876183907180065310803612652682707429820522544802060219717174049260849377166333637832636740496601870303604881833727904251006499526246213438970770765580881942926698673929281690278951323288428312902768288359071074016326970065395701025897715405018028565826839317216524023778269385986277745167394513463098642504305076319007398379091297048966176490410932937991990799221850327129833932974574324726764998708434868740969447311800007938802840601357828389037315163352329964871613931332569709908165242890586414723097735761623238448198703347442762863190931327028395353976286424340267944254242241942933144481241993466446659963345537124336213731466964727284341293937948144492597175508642401845980199335334128984296173739887932088865;
G[31]<=2560'd57780413681355008640628930113182713118747241993654175804706541179228309369127573683999938698569696370497457919191008525309738713355954437446092296253488048015950072461499178519770094198472828747955556172552195319385416393636038336560417226815752650472389175339736506613057520632806957096675755367695869243251547227224463448019456243774915540885018416822863419255996455082625003472486060762262167339190149400213657869625192085703872641921115340893365940566305596723342529720698633662326534831363338813085334000811401643293780431883150105326523729919078231157666990626819444733238068056218527389562239945067441420883437153229134808970914586304085688681782559023526854160796150200587293939038236849230413914109056006735925216710428968042658839672225050217231019953394688545;
G[32]<=2560'd57886199865530329942500979468504725219262342551789626220586234433884994531359720903957987564301759284542441993091597089985542243633051169241798870794140110060464323935545682820563220851371760417112120254275065071192389442875877162959343946277945033712038650295618237360041749094450278904438694185100328189830107870039547044847311615817406939967606677012519743999345986633472814760966260554017577771477582212964688114449815403042413588596400265773897513874337488853541381155526932798951479789679057496543442746974849694243507004210082550434509737885365905240630491813613044925707157164854190859053948734208347143550475574254940524277625755635700828501877065435356060265949515935868046756277208794649761681666222814751042245035568391938795575992949067514249231137648026146;
G[33]<=2560'd57886198244661828510717820946167075054661744869106085268702554889590085950926884140769977040184220190139012940920188935375827133687972971161180844255580538655677880127167784186788911386627692921236718485460501909456197324405866695636816868275550904130651611465148449336819765636841790623804824991842553473189280410376348175148769800206246586893469748927590092426198579833753131282113218888915999195603334689077477667173091253546277507994270350770720351478216435103743304521535297579876460155617038482675715636854834764778299587159764509387870682236264552633617673952864527558085635061734829892710773319418557891109486627507071156635589183582207479679352539459990922440650724917862492781461391189887234322714568368312192591362479396334981862285614061863909836693067407906;
G[34]<=2560'd86547205173614332816597676854006876673828861112006029106104718338021488086319260357628662440212863533382706568147029747530161331968736551366646351126184278545318883029238817015117816716152439540122902751962647772891802673978839265326692502215233361755172495013520727430124014315080752769276098967533807870505236597722394816520752249939135766611637287785242935328908543901470626179201211130558378170088788281237966081469156827677123939718367790698186918717123622929182531830679162787537947182123278220320253269806216714293920028427937999227561660363970818641119141950695240124687560268842391446783164413865589513517134934515808041262028035705214877863983036584553683309786812124617710672155269784950114771993987457791036933796888248539025192891669312025041445112653160994;
G[35]<=2560'd57773361376689771640823383541146674820641875135557686375809918377490925896274175771886835779009119012445829897850514739139367697677230512565121001098651049848281158363423575448704338953596310138245550700175615095503221166721457764087001592668020377673164499299874225816933830584719210098801882536817742789336583997703670514839420452191368232884927213930549656626714118841855819495705489724435573353995723927971600353586470542664683069599005486081779756057562287286607922298551607642747641336647721244126282049401819907658339136627923403590071666370447904965607845456429671375057304781051754315152755700622566356438297372071129100002612500246357226579540685109458527151937167414079700153454076079320762181876950410262046527407330469767412667707042179615111526910932427298;
G[36]<=2560'd57886198251359823119006638081691267587542112734823965061610623037391202157803115475415536320492323613731423979182718487757005503734268283504487936919078104815512879911770451515375915885934213789432923363804072007271723107151171906513727288474496254330884483879377053165239157537327101064753763369702581193165903340590408446928324079180197919450013856715032160818635122045503640747795161991307662186581212037481291151228927537799176912203291843368146040406744232580418714678888970654688312112627363588453923143766115828822729031959401575910443405909660339793642719760284786049510400893492405064543859779738627237800281116598720888914767381959398841655297947726699818122847513534869788353168845885579406593484043487771918654972327693103028851851909066264206671779610108450;
G[37]<=2560'd57886198251361362884956388865772942505349142361011568304536944642532825608609275863530084300564537482524051045954764722440046020388115257587816074135857998118935803149384679391100187492299487974666972874027731499098130286355031379774450606356847085229600928905367566439929203963276667129702297619643090131997664219909891562888183374723271533173847777381691614987168625654978850143770126262442900454123067883181113784275584675987997273177098527214706310398953347579764506129741476605982000763834511910519819896277018530589043427737994592330564976826171245288845736986015834338315999576084657672524570582069144797650123697203622341891479716776735094324488684274768408590278011902297271992909335513766118439418053524861196237018582435903010529513927821236328914538484343330;
G[38]<=2560'd86660042048680007930424800345681004176341087990407829576227206209746178345307483002399604700197562652106164500963212526023189340038649793980339930972580352679432083332034460513087123591385148125419820973153328485619738159549173698594888409282211571877357583547142898306015112072350205247174317127936755770312411411693586027040434386623466388350397529896710233456477533158749789138680995652610818576500451437259063655345821948860294348868394977506958075541074921727366642595922609965583749203239356406210815096373212591342724953449309696679918901494839009115077701494686084580568767530838380572751595092140650073784987852400515678063033849267804834436483895136116412217472711588333051971371393409306361690400103150870117496165980206234248045291160861965942148633712534050;
G[39]<=2560'd86660042048679905706670498856373919482003898794175655597186442797913916598133336510808291049470179530826091433244407161837483689279714717458983399068705608718463423982668844191285205820308961360787975730947033228784205554511973870570595400115001404958024409040150363471546836510546252112220254743349592469762208251818544966223966506781345018860860372657316735475663700807050157946346010571009956211765691703288836572059946548020617996322140705043368266956776873543059031412491587328380629822282492372629303267348342173169253345297480883465722242117419301415402591205043151548128163893523847739584571124184305104389616741040570007023986978585829369486409042765540664523465812738604160994690648323235147015429313378754547376378805199160782277901230400651992247384439661090;
G[40]<=2560'd86660042048680007930424800350808207770364210028497301754987863923357610205641372752935678039550091572522003041783745934312988038327359585206407063320275194926839170651772835255610135691602168551775290829420238200378779123079554976408936152257332781996038037123362327117539134741957429672217060409240041804235564137101809056731910526844491126094189188948461662103521570928142203358143002428570163069986949953749997869139193198907139767167871204222884272790428141546375064702285455706607297118214720164359224411534404674296895339816798018614397846225868141849272260561843913359327038154053219650426720632769714494197370102395743588084854312171857729955167229401443802955303810997731640855566890389625240489582995154463878181999214972803938474639502074081012871465137218082;
G[41]<=2560'd86660042048680007931892520149873807400491986871039771509184460038271334125267982493978923024194940154785157601869620972194770800722035832975423122078395569578541867574848383078727147606562615679522385202966964639204835346694710913062255413787572672283866051988072156467524611715182674362647441642006513833187208440702160149722989265282912175633806154421244849949726360240496799968087194066513426619308970144848505337070367936072532594147783053654717921663249152773176171907412744127310608627792249177502451229167428495730872454357984598449845549430027421692292552886711230882632306017804662922059916082752788015874164581842542824957708070717125036599105414948250606094621404683868124026831987692944991524704476683897398499820063823090774584083342223360698587011382125090;
G[42]<=2560'd86660042048680007931892497743330318551888086268535203559603953441769403432097744057686600165799285004693908652298606441974580378356132249784747880817894661406182914340337612737321449103395255548634327765664635831759587097516789695604292684211039876843469739824805876449568267560585422605835535729535030097423010863997659361251958923996503899152082566960006768428910889079586332119143005152560948804893238292324046962336948643652418446714296728377833536365639073129899532850513254608675801332265714400247117818624953783022994023433915934818755110935423999759147391730381806265382610545136879302785342101605266695462556862976531700785182944195522406297053197556783027464192301303883549169431263102333241514726988110648354672251150807312009905258073014901885142495056241186;
G[43]<=2560'd86660042054985355860246763780396916595139182190559466635839068717620643410983751612470973283878043979682038317225596061411597801122422374198740999968555018281259349058096889367285539329803776264017294556388629227213048382211949399230713651452609736672323414140581408963617265023746837550025679202405152140389164706442121713283826430504891216959352374160376029740971943662039106710608550413415630605525773289228953698323561448539950494931644464335216647986688347306402714011952472905140060776675150709962334424321591111899227655998383061642129229624306436430986721559692071109299575757639739600840157008186915862496780206541075407246397818893784681180175316913578849787488901905584619042841620919470650133159830882409910802025923429163225524339952125024767402361628008994;
G[44]<=2560'd86660042054985355860246763780396916269160334582353078132005935403743489602691486280209604110762075032424719011073747437388053381021371005483095637757542075924062003385256723917034785986875967151561658751595043770639837459476679911982232481628379789530947174738997808872157510708946636806088920525165957039325218561570934317108747938136780249097782592875767254241488565205067232586220883402529424569300572553643268529189590555465755051011317267163035256224075468125950843040081584207287923207580087792820889801474417518264917943724673615212991298988540099568322964824683497540272962938309202119133293683989582941709871084086885098482064614193897428738618652714274482302680832113905815511393128946997365474103712990967494320292947876922398638606109883492192402488804123170;
G[45]<=2560'd86660042054985355858778685563434785797141114242058606618279755029643986252503841159238337982373373522297453321708239130508181193587222639643175785141262499175365150930215420476322445313099140979056554663258885464376960180253595363327869146774646048293348241851738589776482382411546458591260279200652678111827201917596216500602425825785734506640757584716654700261918021446821983830852542954649983826490495095138826222757346412631606641200969722826912266526057138326855753032592553269327441363632816523213364267098067020947763252537789432485641421847507823980697786264267176201037859119947553721497384684460383506658502280708795646486055367638096250286245814750100233639831026197252572770639983663269917990114237885335568394672320313948658686073541491198935783307410022946;
G[46]<=2560'd86660042054985355858779066382405788623482250413339828470726677404109926983401609525569057367837882879673716659670988501639059061533190796507301330288715979317615683978991923161455227764577183962619778907542542109472554094303208349837277898053186647821512372423648282563326024547826524863117877759415844814019055182358143940423187333920642170143876799721844601413204186161691363458288353772713795744104982268007109471638230998766390143070893203122554730045298802080564234751843798225994759853235839194095432386979750447943741384743658650779508547077193013475970813944475127315017307654525089682180161533648972774299163254859081500767493269254686087768828885241591199416773498659247008239352651124664780893748817581582716583512186618823542017140265328915116482299724702242;
G[47]<=2560'd86660042054985355858779066382405788623482250413339828470726677404109926983401609525569057368668773025623400662470388244366892743885762918170070295927483656670800818907337668544186404805592140459291021099327367686731256291952018066407275993315670813347494785577955399276487194650408226703891566795138771333928359675354783538047558374066115593308217645274858075484253240317136155771767416228797557410093885220710958160720553639777988533137201727653730245843775918844517972731772271242985837118417244787913808585553420709014784645638265834807526002793998618722358228203581774568486172236176320791425354577624918312860363721252349022437596724463935482603154106675173606972682848715322131912701256410406167811418028175130148382228617059462605469627935968313951974811806868002;
G[48]<=2560'd86660041953681068106635190087510969713440941542676464483039772789571657224392012532835602736332189700746550521647143070512378250592769974059210208225936506010129890717310579264561821424693774201934009037606695145169579412924506485936819184245897881768761893399790443063072619005679457830464831728868427028195338488299870666971059537571240997379793854034426032495661859584850481965099782141472667977266300874312394229603973180882537427451472360673258426457664712771275056267509506865999871746669068012206726090742205757068453733365517719733107360775319570590314469875004886307885756955132495717927761215427428718502887981193603519249144464508381707651751396031120029497271158946974718152538989190001623374725226670535215814444508814492992410851889150492436499064615477794;
G[49]<=2560'd86660042054985355858779042580899650700482866746678704041470904833733252705770564303813670944804758412697358339856341522116479376847005978313110320331129082551712200291654589377646395484314385839419833649330714915836425648482795524352252297710274305800723421933711165455647250079204721682755532120936562128005649608726034722942843790817281561864971362223925547390106041092159671008922259389816604286851488889821051840777191447248525470367118465450615288674990520292540887701672221537125054542909406921081405933303903026407698916964516177325423005288070893354234844289146950189296943220095384495813269597692297316840121679319147110179317869518231106459751515772457473682988224202063375939039064015566192602833460870034510836296665604547330546357519043726408002409414664737;
G[50]<=2560'd86660042054985355858779043980968140366770481462086620545595401796867242285987613106704994512471427422609518420367343281228865439089590763145994576484637848798146797928429555580067697568787044605904722067256150036211992223016792815597543373529270477752378208115103125764767289351920362471162881962336062648556786164643667450349270245713163997721014453671779864593900645597745677344744607891290557220722794821489085569056788105393787687549248706951708757226395505280418501984089322261309101517215763782470241646217022226204352806139378669960440612452417474836242259436480489947332242617236069416926492520123053545384099127405148844865968382427437727048914443141877717066782492015465632299338373606007217998207839972801816214101341331188259394178043162720768420624554140194;
G[51]<=2560'd86660042054985355858779066382405788623482250413043352435936699269989113289295720328931914268360236876286703549620207161845743995848687972284182021581571963249461170347198537116720150521568196841670154613461642106724424343503426541990099238091052445956698245557683529622491838211463705697014712530800572071296489420018433822141071026207112230997636269996911769012252172717744846473496606832186446050599195978858900571801623932933941702494693701636250341205809441503305063956861696266668222810482624494016976815333944599894284133570902724027162659038813429950665570787946319376272068806772826657803399228027775516171968011000718870389947345510997219794280156784192631387646782193353033551463137019055180906303330128059904681487917990145720358641865343028013328464934478370;
G[52]<=2560'd86660042054985355860247144599026105824097029988979998940762276780325789130097412983589890060956835943811174128512144286711561552509151793218700130663381006090596347712456249535970544951382425260880999576103080253532286961330802656336551597258989204139046459794367867232059867562542042259195000808293139155549836330691145335769872881982597325860974691542243359892521873305329542028496531215507817167296821851009314637021303705301203311802510459399997698577826067418921123933090242315870125008614593761434473526081935722342557341645076228863805822445748326863370590851443957362959409675012813192663313938274266211410176697464011428840929611838192511579860650586063302923127187381674738472196365774868982457452673503020967358621030659055428043928563942684591420307260187170;
G[53]<=2560'd86660042054985355860247144599026105803723352013448569907098332314825916161197528325533736446466802263249853318558896444694473167967781433179911322579735004264415448757159607884486251350952810936618514875423816401020935806798414247633452655310136172884986605128864547303560169628199684359852190075294361673052454449545562569846867922934291145837093132908418921107393086182713271879202060377248661168042612721595942915594912041817455848479559102792822809333264612690868644068424994363203591589712725146368674504599885808200393699176748664471126639761023891752123537128100812932515685717003398818768846329897148320503360070075386091115658994810879691487893930201329435996319950187571744456848164786539646008310179080421345728263409910618014426229044018717371625854717796898;
G[54]<=2560'd86660042054985355860247143198957616157809415273275606401847801683054913857724015869745738009495520426496013595254019616276918252706559036730517567925473363244271953587105398395330906366393934964797975223198396016120608260661861769916522741701562430487704802565771171974121498748478756099811215555868397146141947629973775578296202785969350407834282082659824478794036290976727007458231432687636371322854234783724576756840168982645647592586325283399145531717890934896224245883118321463189347486181123411894310714608598622387317373797837423011868063478130433130658438155209134363490799289507124301229220315490872305174607888249832083008571358343548194415762936850371307920039557656814731410650870255416906436886636958771533394917216612650844630355500677524331504388270072354;
G[55]<=2560'd86660042054985355860247143198956280949722965719013170516182992918348259992078620245111975407102989111853916578911136083213718743485772775757865926940684976263945545095835835188288633478832728556506922216040835923396536415940403762396032571662521575280428911570127456279089384340186277286753913700687373968115321928218621365620025654220377864661426507486449019759142129249239478096336245356588196548407353030685718024443562275088829022202809914785289904365204312582236277314656335398274506109220768073106488716455041809752306896733531144310276814905618743558243836120827268793661427595130606121998647306549936409736935664975034252464923140002294332016259704076187707574689083790004804657815154570100538770143114324124284153631092209864453133829764091307207712097018454562;
G[56]<=2560'd86660042054985355858779043981309953962880414962069547848095075847775922625427489582415750862091967253328052725540206978325213666061739810634858717468967353304268472712834328044181562989527012538596253710812900954806040517669379490114845623771986123640801384449011394718498708721114687868235859816605125059345700993619764063046495890656224728498081090665336437849144552598671341643630041412567173661725035643574674330802730444146414903626867336233063307290384715540514927540493527168620502825629918147969105637112564149048525634140599476248418606541400736159309141458345063456857152494826856689973428975043227964087802898167014490378516400034064683444741894127522423793142833465796575689313408021018989621762729227017912525848528860760229580771970275881552674274953798178;
G[57]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653889653071580632085654872882052773954860466945031344557388528491751004815415037772754542432001558774931037760633855271045753308239093177283751596238697575492571877863587228649850810627442910149468310501082325262472746958994887076736180610419273367717968381675228900809217769254646675822531975137636038620897956612191230723601761079561482789884126472727012933821701461639816945634011358402017287160713397811586285965706088767883939722716158734901187625345536477908742564081081119999404687937241791681756677956692823387750957045160423229522328366853541774990458755201168200148209490223331170614846925008065789226289753329394830035797908724518890210448878089486856545510497383360217012571350376994;
G[58]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655774719271138450876403253247980525681756927955966313408893360426260923510851124225656679336182992485485582553762903069025764545301208114675219999682369604280730677280663085198483631923891355892708293046662423203514706204260985181959773672542115924493013880045541903868308888110937032782676668021161123182781339203518315111239342409093632303811738022643378105828812942801845280177714538499525275336523047318019422703179843371536885370287948675884308699991415931439016261119539117062677506538690338435646801560327307770818536964588420905074823861949394928438047705722746387671863216717295875754698440463367648245777249910330319181731115072248424154841342736256206543956355384186676383395750178;
G[59]<=2560'd86660042054985355860247143111453335554939794227014796182769643518569226213756921341259859584655847331927551925801083113722239420023735037221501403343888797101784485428091297633820555426628132444240443189637533982397144847074286545063728176258437372280520181472519077892055236811898975030208945229754974394771557861532894593339218546953074265959782279998383053459704937225139156610517274077379498937826253929464335646026284249469511805352044913585632132636556730659051006616145226591426780570264289309424192224557073134779761862353093720036827761563695692023726541237184707798368999946478445971640413873826589891622623607877163896854987379886470855753213378759358483658500020978676937666804110303889982458638106352172301500584091171059591696502376120599261557794747326754;
G[60]<=2560'd86660042054985355860247144511521825221227408942719188721684118615840101486130318455104011422578788422303091856281883711360084916977256211647218502040761647245051742863180649101461518057094087840151819189108974499674057614671235616422250522400472752448260249259811871545899956176160760290117877614210040413383699659879470926122939900051338539712209862023458245405854678800980242689599924078883354409708333679516001107317269852292268317850954089206035577539940725260913867976686933328380837615663909387119286253829702699469042640724440276197900248930779584646031149548226901857160232709144580209513902232730073611422576456572841936087366733901272610561546622627932260379133331353589838330387301273102999180562501618591856542526039496357707062027424395229927093319338435105;
G[61]<=2560'd86660042054985355860247144599026105824097029988979998940762276780325789130097412983589890060129178833448842981754766926594890001379147084396561766514151442423472671271577733176472177794863122290117229327991146330649779988599876270363413514204087290129857463895920198410407913527516136848088444896902525138266280326727798974060509784296848183943798204047143464899439906939430535322610359458495582398461804538122504965104670389639025874127542309375805503055588810948109769636623272370047194653534521086637647811481683316443839443005819800083587861183169439250281450333445303589191044020564224250397150975415711283255824104345418673478663530374775470013642209012515958914020476419772885412931890234560281190493717948886117424940064712916709621142325535805826320419707298337;
G[62]<=2560'd86660042054985355860247144593557088286338093993996778657407142111977074773564704401113994398020312181502375568673229299213298229086782089927547314589499022370200138585108553134264391182968735434152203212672921688901567165354811641616822544281512587480774526369703701706251433092417736083204054321384018794465260161047941010186812917382737087082984730047006516031777250047573064756337075046695917698846612860215428814265313819269540558557398439776460634922058612010320567848013805130933410846600838907792128411476653137423063234254767648774077996288412474606468611190359475636498202924225738676648212226453382000176794280785008176911571084945883687709541639425513238520573787005622755067570683021279389103337245457078656686386079229029317081083556429232540624452386431522;
G[63]<=2560'd86660042054985355860246786176023733696335048798140859661637572745133132077075407094941221655193685997491958710066308711411961925220130909958373031445522292385843115017774306012077355566114773688622847285383683582358559077329159837360381247724659056980258920352488570206225349141535596460106540733395603300599394190034753034850680128499067724535410393039934636073457212601735522974449253511152783567582168443389058870214523663659786863532614635066038869152188286885842290689064308722891679253317057604820768562795974105254950073688806397090219635756580492061551606914753115685502866408397124024130879769520727611290296888003994957005883977697732207336300379910097062204497652351508726415194368912322176652722470555414059290444593867646609145355676250843675969867774829090;
G[64]<=2560'd86660042054985355860247144593557088286338093993996778657407142111977074773564704401113936328769805573782886599260356634602809554320251888855117705326231601099455658690652688217618598901308434824433943915474864242467205044732768881459294144747317318127393209868176211744042545107818486254329886225881362754804420122997466889865379698418997204621840137374200345484093910976585121423400729312662713754018547441152143030815849273285047428102015827044190904933758651140459233590256543605767314173462727484340809640017929458352103275529290362106411955329236895162689862028410220062252259005897122191226141277063379468016527152272099392107451889430174137545550752082926851448367363116329287114974239064637951004550955224348074593717373293924037810464159181395398927198749598242;
G[65]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655774718399874576845311263545621133587374865287058419940707173994009136814956453350768510203102348981932650334168318863929303384803598438714880777773760653438309467308309674333580766875460944163258553664485399703350512389689746009152592891465470579617499246392134692305691882188906687901755226684312602276243870296708998556735964903520686379328169033984560048037094463059281215297534622478298795900231157184848021832456550484421748935713389747084723996705060202625306538106371830740489994778052864551373399262997900463051727027345947204393612565134831068945300460823215836937203120825596631300219200737609154155615517590363798456755702365997121177983711118824673426344802772334068935371661858;
G[66]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655774718454327790191084627349621299974825006574809757877462121585811598112810101427378909437936333388922662171105735217807267199793425598188658135183563724358032057353479316359114754616554325215643178941995856391230901090859599500630364463235959368824600394808655631443543432810959427618684036401442414844223442704537743259568172663689822152367607873679446798919686547135026592474419271324488057680884899658831462461733081526158376459253335403841000626453863934717473404934807137378114636605839740782529376394370848128524048014330580593944144835869571589381734225118077837757559349421951348300910035413251463717639437790513128612360105192064213447571513325311286738451712693242898172633817634;
G[67]<=2560'd86660042054985355836757893132759216999050300176990105433423042907694069227337621562829993585710125964775270602054329570312964848286606141500531370409080004217179229087876458524573909993767173353541741569983690097011452215581692943335157711625082337273452088155362138289609015979491151724013197270317567215016397895589488143744367408171640028233148403530609947223568923703591532337434080808995551208032112472717051380803676170184201384443075252129804075351945885496179914149724178321715988304098213391844187969658063265840143740972682405958357008644602236731043709338815233073262675242050602336722143889890945319882037542546079300604375657035822322658406853107738162463497108344086946922613949873220305811541439403656605271856895022581227425901414826423958301482927923746;
G[68]<=2560'd86660042054985355860247144598684292229260451362764261987656577392647736543370361488313710848856671873072791647228847401301233737022303104481537360942050656559379109093707203561310020078329455616609213664298073261692643884024823015191459955184622890351912106016648553401819722104181655546115603098605602283925052724782344142612161115776715102522772726678600693028614344343062763923568836896432823850079449204882648266403309308892407135748887072114713015499792289361892822207599883377413424244026019710030176048684613618462378857121689125996320360666288608862423331095099705296092543804564100124194321437686435841939382768673574851536518314568569887782433744239917473763412468844755838549484650598041515502392695080274323693426528701197443020246240241189182231408333169186;
G[69]<=2560'd86660042054985355860247144599026105825370384862450713255361959015294025087292967727262403019761437556893730939222285479208882657298300802037575160390820663446459910427025464988327289287183046129933888674557455821371193766728291409567502186905000693240486376757989222554571598683229120888859653263524696001017833907336707490699150744578210589003292255020429401758824390483464760261996791101039665210830411698043690738605065655946827548868455326266465220751831286515792054482699950551567349497745834860048513959155597774589812378136743362735191173696671071195226227253589540277172586531673396101711690290664997436114167944396052162106362849502501002874907669478497240864847453355389428257027314580058540716784625166937389844633065329991770550966658389420930642393390260770;
G[70]<=2560'd86660042054985355860247144506052807683468472947735968438328983947491387129597609872627186651582024600194769475967913546040582144638130874376358646389318118814786852448844864649616750418145221955943826192993427732227178816920656271276905585143533586373115519879198834973942479680809689136819032576647810312732595572241699987593350080061015163659514017086081785146239875106477794600524685253134995910988108331550005681068184799601299096865758881197042238117027682965568176184440972070007071685850278791236878233013284058261027277045670555915937338480331575087435511173575574829886103561003286505600594130697069131580070588727767626265269615924617269111125896874772906631908154138492523244743476934718646027340629865652900225244263688152028139895812604781531321130020905506;
G[71]<=2560'd59578778805611415146675009581581710277691063045551933687756480398422287305889417379810347486441127485821052919679468113542889452684809722395700140936045022572934856316740892564662612527775299204707218185663838635012072754076111058190931232646246903284622465844734391942262056614048354950998749653954621708730071231384805927464554913100265626297716474520693310320586703562023117512497681822088322064496627431618705816210851000079439549733964673296766382384830234107507829212973462685859580341388056333822408667819115709266929113949331942030765735241154336105484549413082790808164475594849201598380667340462756895651089301958848549135503799510269852440112386488122331536158859401750494586734685718641628289919093841766310500080242900024127710319686136400082430937478078754;
G[72]<=2560'd86660042054985355860247144511499126662105429321273068407277388151938834367485704448074122569444172098571526876043165783859971920836969264760530889986184214714476462825495155391096180828470557181509827704450606097509215211503688305040483176269022017505845808269496127703269358050071161707092074104791718970772952653536039658534041538746737519884610030312878945046362214805134711841492026238512161881333319600192118535568830711533085405163924568357858375656538450464542581387128911893507230738836122342122599229603225159031928116892112183813987831334078163660952121246700020305227035488720168916218950633486959406908687460877728095399553261757236528956866684643708270351675359414887359595433733068798101071801564818935401427557464124212599737527976729175141628625738146338;
G[73]<=2560'd86660042054985355860247144506030025673766809899539093146316106265538579527373894217208035140992228093770572926673644688048479952434091876761068352954624370313967179694144722519396115596716221149993677036153553749620405412492028321159047416322212101238817406986707224126155932813939280493474565106163243812093763248383289461620019636871619675083026048451029932647327890463018525846330569091012827951043961281840363813652720803421450634459595725809176904449959904946528405453617565759058238372018608034173761612594819174824643003666622470359816268396963607342574155887874068820379188517184069791924546505855719533630439298370134457181094281013101904021478007737640291588363532012684708463746009272487763618777157431999954573528906051437579347480856254041877843835921506850;
G[74]<=2560'd86660041954099789006487133204903260360956160549643489620338436618377637842576284359863362919106309704243689707478965570827087656974542979942899829084462849611710618939249259608651433216280325477624001316104317596466729371969140954012690077284070616491746351728564471749830002831560147671056706250114477967642600397569096089333639873237374815985680449617611473202653341468188389253981682060228151357854826269269897619172307658620798233705706620873171621459991834543602373480841465702572766633951399857104105277494966054984314146440101192436966681634547904932513426545098027989272415738681311799297143377554507886856890818249006286001241109250814775639853255995094349878596934873475517785221958114450158264812106537624759494253032273056539456887172795468571491207787717154;
G[75]<=2560'd86660041954099789006487133210372283094002980229243248581765007654265653577472194899509236465242444698557438206565622384997964166572406234100477574397674777977505156139830132600223453848556708268115839502061869003420388328807831387577338221680274160140737353483060194004219894535220492435436638099083021936946939639139967824451702131676013475962351090698562849120246157186119729566585232078263124535806048274395725373153488509753826952978246979174053340621456186806072963532835551810894771631448080623550609249689592193110569192389873730482553764511745817030083183665190218365690879571174825385991280416004869216602169328363378343889459927877136698575477417128475210924716016187864188984710543742423461974587831700593124739970235920631999071281594898656945873596513919522;
G[76]<=2560'd86660042054985355860247144599003407264900768742917205928978690163070087408492480637134593336424087829180468219361015914975598451995323508157199382690387690692398844843514928702170390815955241127201596505186844143653741703581129775648233164490994829785826559032053443722600385653813081705720571192837612192008789895713581204777036768429701283390029128714492492860866413535988313649888274937865120070894133677752082007591688015900113548459282696583556119301935464465004416053920016584001304036307935383388149030247634916924973060160457136266216231745761323108368693178494608562968755471783886477741817760726462323763538431370223079186111408194139425030021432821272200460005743589200945611397882829013036913810155655564988139486757628315312202194418455979459998879175549474;
G[77]<=2560'd86660042054985355860247144599004742474340157850242275773905930945813336110118196240539490019284497147557838267018715923327516985332458326214162622923935032900007250338680321292760895710080642733831080771132276743829180253147307432997290084635644489975363748648430396123195922767541394877112594560996448552795364929996576891672177881015439931564850225635004154449269300794129689966712991918235903256491757616054739473066684970639531734216110210497023947756414714550996636483927399207975705990206652969886904718360475734763919556982928349895482367292716115476342446774992956956151252498761107452974814663281784497534204432083595228598354775546782281615644757523107013408384213577019424866752638179442528218812136730985593652630334269396304630857438406952165630624722461218;
G[78]<=2560'd86660042054960725594902010747320149636123739696737298068478322537961717678834482520817700403422358152770703089804200239874430140542010196752272567030863787390542375799084797042880740305436258738701590595005273685970718092719258284346416099842744389568146106365680795020940108979300459124745005745541606269281975675153401601355861428425322813332853822314868282860085603518697367456251787738056850481336079477469278919551948737819618090357466945106174611703508873103241356755282912505867187682504286195515332334044507939923872067346420391291450201267737307196242266351701053576592209146137362958009141113321913274469153424631734344853704883456841716171248282511082540215444006217020418174976790118549107329200324022701764190600284643805639511798376487134797608217221407266;
G[79]<=2560'd86660042054960725594902010747340177776520806112734551072445687533085065021448737070947400136664116789823449632968933407100211141072534280403769520078569537007792782613308474635802174537698970690809478334163570631412643605553283048347016505856194742070928102753525115715195323556349282491460458912876425113469267946730167935278877587537012328036693322053917166377186328222421417452562140040373504779528146445317702735030594897981370553186876005592345917970632889970866951268394574120635906845248615646694132609550556497211472604097622090146301841019284956732129290307426459296785387053797423353574007693950943331632285563368237321343236561559080511485751047627371120384481280497045687940783478938756780680703394917024408763222317734320903198305034840010565975018362249762;
G[80]<=2560'd86660042054985355860247120704888478140837876365123543014150374342850668582094621300469630599648230045742933784209142216389575425264556457922311286053930068582254622325112018075397164352798510515175743577017133975096924825280536745183882775463013210531701767065164325694470222681879094027781227092124253891209974256562213127667449952245758611535158008384943523014702263896852972198345773215598825568241371935340033673140086260660029269570701662991495015670057665468054858190583839025745492539179496075518443982113647629562614224198611078900088975010185705946430345852047500388605612792166307171121399509420106747531104482716050218417932545935284048716286685620621872573041225179656281802941603212553170821511940296270997912335104981143764707985385150670693967840854286882;
G[81]<=2560'd57886199966415999422274459868880719125540374263590124869795440374651327475006935105024159671050131151629198127377876542703104025982922392775671051129536883522583656793447358129814165503768731187588849792514834040544807253935283789448867402026705581432365375058772472597764965932808718781213030096311926565294185957855310110042521569562205157534019507819107854355152510317494284522903983483964605963312489473798774998761307931619933542514693985202534158387607026119398615428324766398489587748219957943248718605013661819049738657691700116659963079334453258255115311280263377575270159758431180536737140130835363759448450906942390758515895892558919289980424573076460337180917149852867993710505728622602071866521405599262333943164274023264992321184253293518166190136775287330;
G[82]<=2560'd86660042054985355860247144598684292229255166442635034168043483571173619710347119691144225030345827783212616222410294779761664479303518996925898282846266761510152391272741003190926623569187827830321629584262815111917596656706924087217393595876587508488968085186850687018244869998586114352220825360249263999775994728817375979812312492335397673203863302790066154748820302833669594020234290070582495200494929173360892773760163848214934974637634110348177502057929162636868254278830623178642620108843250787630827113236425449731118530688061698145372752265186338644811567914707468253620627016699072244012274195258088502328593653161690728502743258132518369470836368284298865727335683902707471302377458690498583886192744776199938910473963751447473945313840479367679935282310947362;
G[83]<=2560'd86660042048680007931892878474455227177971028024371356884811529049464620789125649758454898234272000069661172069987269389899945767361027574550972953530686414156658146882063111746039616309348358824526389848093296029675936468034120445424222211600742719199081588357825713506969184080579763331048295605712708386042479337966354451986290223333162107928880627555641215916709142920994978626416705217902414635832264440558822987219714564201291986753954932486082169720587931507557958295163366806492875072812759787144098478572127948308523884977559396404699160526520479526138165521289185352674936636031862683817235010289653831282257759622960847192343479592912613726360950245590935504593119468479652345238828060076678734350136759719261592194605077595210590771535247821334747701596791330;
G[84]<=2560'd86660042054985355858779066382063975027367342790537400762351507145035035354631882491076581761791269452033454183249344953585965394076337935338929067937815323622118536437564297059738643985622505820504106233814091760776962499864597298059636168145275156380296688159904369128528449753683962911312799230433778806225091259387969225469171675201128841950542531180116230576449826367722593526857172521687380991124864003137484864476578707170847913234971151192728858579471574281800440108831643342639806729108253011705015817802300804819006806509556132826791595285218890642917261770516453191612904071342140210892697080297449383854621207259472932253846052618039414465244459335409020295559531631438526291491079580094505907840769648086836318006592823881355453236395659111836949496283144738;
G[85]<=2560'd86660042054985355860247144599026105825290800106942398952294747558040315764879639160853610891343641288103171800486690726035351073673038897420098791390589178677549463196067503209119942093911134633742650281137952907541928838736039120644646931213431112304087705918212662505290465616993101515620308726321822160039891944288240508538304355195681045858672879005331300378590385772671636360499077146404297835592209696539975963729580103811198511037593977261690843212160678790092497209149901299896578574417450022512314644223478594860607318104626614943274593030863303350193129768254716719146242445724555021203697150864406182823332110787462630238266984160936066412740342336739627906476212971555791033611251789021068735798176701954453565289380761074629664307338427911253556960591749666;
G[86]<=2560'd86660042054985355860247144506052807683468472947735968438328983947491387129597609933533007353684341990834195015035555132862800169749291769193498400956334536367377488232563817334060775311589028319499004636252388382801225987419238993976401404890105498706757207668415650809388003583954191261892980550012471897649945546194087881745460552090656867092022397398117193406979658263660999529979154606521646016363548806246759747276630646428830254854567210377701679472127092615248509550215121741755238221651842306972526149331062532715833584924367662404364017771944166046262895022778674661432141777272682723655851838789731391531005692757746195209800003240536714795470478775228159959576119964382052626711932844204986669243846253798022178028122705615451830431736486204494364140944630306;
G[87]<=2560'd86660042048680007930333045462269438292872062652782987313219768042637666786329122335958460617666226744102445578905364904221461546927122893717108422029525645388751312472799921351044500286877869119547669424756898689829950269766031585682350250802738512990086600498257138856310699958638986089000168219505650452112645792298125168043355099070288093785806974677681179875429651395058070130055538199697219290972676462000385767399321028894749768463796500316714247386234917935903966874879825735126556867490207321468054617049686778077196364220332825960605886426479480461424307056476950210290425255119077691922776496538179629287074916631800112674371952466862493794321215866845955683019940383199952142344488797901438377077613337058870934732589916097121038462490224294365744145232962082;
G[88]<=2560'd84861675209395134570513491296012588649149499105406319276736838570015987485756327961237633280414293741586731088976136143971972148940487030188143946429331268596433194112333477537741339933425127451231940167631068619325605887688332015316319583609062672603847286089448040649878095409164732735514694117834379512161136744289961940515034067303877205568319487864466326362184366844823824809603763216310873172285098423406636309344349882612942032817949443939487405824542659607168917833178514602112722803193492521142690442570845502604556226067924782481702160068820749451593355367918058027239620695017180092248959471178729969370265186115169532639379003653673051828582053830937560743687402763418693303907915927876440158786880604316169809002092108465290557910498115674775230925158621730;
G[89]<=2560'd84861676924448135477847698291933182969270109803559838263045818748479236104726770822156305517351321399152115381979039071787818598716118036135860369432465581798590108041026950802983592206926472677439521630309520808261520071964376876911173288838687824944292629663348023916598181663572056578293027286618106951985009644686038524100352294176314053080020437289159049437202541760441256743419125942677251318766454387953219030481403938808193893231465291978346670562009458062889225045766021703107876705393757635746182560538931793843005228315976760083046245520245688136632736542795252716739877679042209407899160438100649596451131403614287530317799995497836201197236581716823302975687026684611433470991825217419400763670120268007613444667507280889933167337023231189938669135715246626;
G[90]<=2560'd86660042054959186203317939881611136941187102524061743979684747305773603167949495082644218922157711575560708848268936227525968118935853211591921765680522137127820191149260207795389301406102020765633560123579243131498054351599170872984982647133513671634994692496740942454551662383337005529259762188189428878733662351435927880904894491560768552910911077507245816215113903432823048028335002012073412211247661151115357362557463804325973154012584687808645567279304741995775227059555612806569008844297274835442906291339343233052935512409877553532908582661020426893385277100762246654990829730243971258313374494390963976530657440076915392840845353560166659051761954419659216317579997726507014517839770197533900893059799519517117352681975597983690176737590772570711961795542786594;
G[91]<=2560'd86660042054985355860247144593193911341744314216542566567950625121514417320961545265830318831687035717921868537533708417470728628786172960835502560281150536811444322540321021624666280051158458527180083217040739972660683108646960734907174923438148809545509677057276475702326359921351356199716725897151800162569169902370034466580230268157191342897385056504582572198246638448441186085716310377152958640164700717121756407490338294946028988439924829548227277968666131301732078578232716388893368676572081268070892626593236852197383331223659582145924537383369215742952515268592973027742739965130823578369112589455882708724300530157063840593092846101088815575743137382783217277523949194824053843845730150941402027345955312396276242237790622227435788695200035768146667033872966178;
G[92]<=2560'd86660016228280241319705402358421350846742624107826118090937600629889003240141592941162634795809343845528595331948796376943280420059426728206225174983166026905954686969162301194931984869673934189588887336905977389447092857165515241705355888283109705347201233459613142005234012111974625599800771935083018002123941718459699998266559529779508543363828271916113812101992832598629957006715952383584774838566653855239296431294017539641105107417733543686412616418419657852779948152548770559799918658169235178764477808228146216818404018453660976131859432179900400456578002928432350073360801616209158185917082734048162681880639888469794787407731354453407252586086727000973075537746408607452424218360384551034471733566894734598966735313839546562530318185257352449484080428085289506;
G[93]<=2560'd59578365685520599527273209317268622070023453496135301177712986741341635673315141329042546278281588768226098689829256776952615299307373508319916431841088991861144884173920347275376591421642204513020731678329283323221134071872424550292060929125372273267239702001936393372232647442856865232732765958910024114724472843946724781073806920839557672830789699016533482169753115315835209410612555125427000915491568577291642802689898551384399112316736957662725821295865502386187508126826164420645561268783450306164099719291958171799979606633617462295216496813388461092598371906806125364472475770339535660341482661053731183081535575920465665746474223306474539741593848911353187558683653706304025041275219738960818756059694581554894703821979093868508043513628273768991527753050366498;
G[94]<=2560'd86653017184888847290607888860499116793301171011115448878627326734944596382599360131154941098967256317572945405638916113787806658507003343093032328610616243448175383590008784736674063062260771023140080532921183005235204347546320093412526250817370916490706489617900013663756741393982631401145874969955265691100697120391588651330718894869146150013699458939426576023837200578906138315525658080824218783059187077161043787456555229386529967448690631820918935253969924059486428940451687701725801934650259781560239744850315891204149294072157890623000546076020047442194170418033780199771495187730610911877115354789131579341469612130844786735220898547578744788951644320964256280188496879862710150821150183461613478586644227222815101456164501086837114136727300607356577347715342882;
G[95]<=2560'd86659628720512608453045997684268877554522436981137869990667778812834812671990664026512525963115700693400811458189923472768706489557104427707402848609635841029425622463354536924521054296828991062482676161379132402879075677623032776554689312060158055139305563396112543200348763700148975881292317137530077161554189469703575559170716972233934984998697908194612401563791075240431997702475321301617185051026974853497646358475438755762195631832201452267395487868782499796783576469437949165569391200489816803188434802137749133069211919741905418911266779575252159184047164775143732502543585929199976812200921575227889429623038538995561017013085720341203093600090225424262375739852575911017191455972907889320594018087406242507336228512974393853483183390029587583615565381687714338;
G[96]<=2560'd86554255971695601011258355623550115364785881895015729348477658261898988411763988058637255489790982563613273956254331608139476278349510695770746689239347307618022661182628740546318887950301788824771317138845423899527055407587740849250083501484625924489266259783071681167449671385959350429745684401329007963736056393556726724101413122411046683442012798464578771725889699809230426554142833133214217107252521314311918868145202167897835391539087267255167943154327172425148817525478299898584580066472738745151499381542318984991769318752527496618427325684601428323230675844822729984438812183347592621683373668246103882097021567910590170553539430679608862796861308746760936053963077365633309556338659268101057225217495611108216923909852090782490363361767496932859521981183304226;
G[97]<=2560'd86660042054959089991343935452503082992633242714398516883236922238997404852538955170768457869218011904834296788013324429273835373608776368953183717752638611392570234202549305848950797717692103387002492062145905723612861405436213919331624853227279001957876648458355649569849052600300714591545060117703648050020246347024814307544168478890979180428323929429202121562570654383892453506373338984264886044242753929183119484302479588674448721388673533382845160526611651236676778340592308594635662160448558304346470871774448062703799092567747718426319009338879306402555268148507359935035683745707580599046153149406325664180690538714384669431464263015129298979973112329470975255037595338111921181702755480919040356647032898303649266883992788258334668134784009662703216373822267938;
G[98]<=2560'd86660042054985355860247144598662928879503580519033858783424721397849499394200573087902534590125983009847885761199052743295786339410417145675947540670243424242185952893270762379425394223483331080337189350036778009575737659908474964089485145433064572712596553730591948375610023845093177914322936561740607913937958735409093987506730441751977527607300103560388349276401902118840081762375453360306113510550146578114423501712442751418917663555626932137353268358423297720792177136873542088617386465465439153023748140473945575311741387654916899680047246097623242789369383357766387040019028839612770575432249383738009892279308207807088873664450993990458888575161127945598983734601670023527837058119380385053655517705650734292308761150439133658551746105854185752914479152994853410;
G[99]<=2560'd86653017191194201232210530174020461615203946404805797402533605310811939325157651693098787039480532549375788446475899353142381063423834360829199483618737578742541979314957495021829235079925972558337686545952528725938401361992147402712017124918834262108385591353660303719483910705017777204887315741330100688627237945688881412149872996970343528222642707010805156132549640847476471890904934223358144403706119496791581715235355450151847364976407440159304802837961197452866409286860418363892000055663038445041327365655658590325571210534058728856125155725464528191427368468976265769829079406437035290936930508516651530877887575592043384621279585196499857018279015857039914752668370608302453899953697656397868065731280477296501686527073383456831151763245751387784426228556112418;
G[100]<=2560'd86653017191192661840626459308311537912492706353412262357849455382068952953697780132022856653801649120043014571473403339171948002318821178269118549736120031837358567315355481062664417623211795413611096659665244752267972530565984769631503924363184121228946517893202331780989908891838015149519190495491028261356651461485254097920064522046720481928872962622347284658797788827658375021590480610706555264513413934185699097295949741837295619558996490596403578334055340826405636650644245273842169050370932257502893749601966591563287922162088861973297830694097403655533653116513208966966266673664361158342693836676240404968647055194343413622931970947674405034503149247014012015607215324512336630374400578714310473500205013675649019033402591413284572013763519485397683984287277602;
G[101]<=2560'd59578778811915325908667584546007890152358405855393846154784101779059989466134168259530490133310863774475876248812450915130807339204008662063689826795174012548144582730092188068532659159010534020584039903446983714115523233876630797950085894409990532388987045342331138301824437462988099477234635280526431012834845898710065423546597152184126203525578595925025084729733561182611142715531025533638564068108751050132720577449616778808388993527916624910260097370490084071896726556272756119598436685178111939150513142448236610593263727916515285746153840820852407698059891120456175355516044856171229960421387935614101499970216269585457679510100513187480237621743364944926118638611963394320420594470864319049938650290071802680836435134106880147402641740237714439110970084685914658;
G[102]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531191671743777336545199199408972725121974067476787700932975915065310524634828185683019126850163311716577502326292494484635010015900944924282130622881883621451827640108219965661238684472495541569757446724817199708381302007678694941517379080823111704591075533418962211249851759250050413312004412204739137369688113956110401132480439661814035239509982133098146557014421426285618318058757427798596153002142793967094515071334475726070289968872588220601961592397108144280646509139759661504920612444035061718528461316160634404294258466099383454243151622385750925755239389396975227594161822293703202295043652868560682000645453040482165820066472421188353893980850152776028839101429313862860660045321541483897378;
G[103]<=2560'd86660042048680001542816121418274708133087735184218121714069309759070684200095528121131151229452618358424989144651244781249476201811325365763530691932360645948103441515413521526728724006714559851654784886348550217802339615546860490514727621003143368788581636201118420867407436792199238362886228157986302182827080889075070645751435640161008633004408806350119647167105101498606748311932226981893215389172688014645343007489325076417050892857209974073944895466807307814604156691105462408997701234236737923122557960891269118741313208623225968015517444427758015495407698015006754716656021007762071449482254245082819796025270672055588843838538620828806404688254174734602305173282201385031777930139348055970663055009810853620039501204547464719938955003477396050364228665432220194;
G[104]<=2560'd86660042054959186203317938481542736267124884929639370484879984008043132456172039682362200766207408574768244696095950217132994987792930293934877870418460833334887952689849087911095144844313777692529905864144415173086656085900327319089863740628222005189876886593675861025152301236300660471035028733498511063880233198761014139936520369798488425025931435221539193303349600462825359605337210880813865978179291685474045957611616411357425306730600387998899305227268075185348462181203705843465830126195284058407379190726369827952788953024668117839489272193540056126597941427784943117147830692833458468447883896467653342544537443070753418354343307170059629087988548003225023167070034424771222586410154011229506311120458614732775307837512381298122729102398736791154365380430012962;
G[105]<=2560'd86660042054985355860247144511520490011867604514986038521419627616166279205998182444861697463998358987853822776346843716112966914068847527346711602336585650717021411204835058777422320613287044925775558102739449877344826082577461742403712360128792639411979967174097852838403878490162384444630161525433676190145748292759542130805183788202814811640644751386953822749611260339977587171433683657436848873607521968768212346233653630822299217509479698169389854718687967384990157695105436037482218880949523542517806967156147050792742821483428334333566006508740169820700299407259315342604161447204505678566524499399286052508665064300973543077745718861877109193534529427765238381215709181802816473262897572959013813020954393270940816365081118121950606729131567706613616775853646370;
G[106]<=2560'd86660042054985355860247144593557088287611448867467492972011139694382357828526350881001422170328006352946738808627560341695352712217056082743129523426239495646348954592534136047416940292394810966226944843910833082683719317595857959901873693888897743886138824196926248342336633766899924865600486164442885449447300906959871761282120926102471798935511581371338443943374366339526674239587952813771423364698580963804213893549215754259347611721358770159825216063359056289493405253002437725128695941331026914240696192626889362767578392361557854683832419575809849010247301505483211969821673091405736086086811363951491129084549438962408628828612549361200691474582804402101596615077354176217779556033851432332009150115532801112221949271480306913700282778692679671777184889855681058;
G[107]<=2560'd86660042054985355860149655029953662886182500934189443562636301197143168485863342094738312080577243707953319893851588370792543370896574288963778115362270111613104282780710662141662175277559670548220191001411061928826163549123890050219712215268113219249049338071899793709974529922831131397469497749812697172054011149298335215279219503495837453231779150556466346203330093031023115862152924326385040606839801045191168797604254064189368559285212928647125886778757249984540128882575117932759243638195414328220129489401500599157698550722830622501728379287075279466730727995444278653312720139734792903997778363838953820261893592952803279252068722217568152271082894028593448730176774764925385809594671070282952157685388532386901578693920989386388355835850492758228298886132408866;
G[108]<=2560'd86660042054985259648273140169576149288481194431819015847103641316569059641215220702362129782350109669493742038905000801475775709483047968337069889665645636944751692851290677633497665775433706884580705425282207594267431225282320244883944801926958973506066443549392951552627029226967725579864037963109740410041735477779833157382391125514000711591725611911312906567241983597929653572179751054629738722084263672815253561543185532775740958628031336433681167157154421222213990970218797697194999248996494664514312945704825059369961568444134068394197570948233634203295397124341005163567029753198056193068728164510818635906955956718784123108507576766126019739906220105454558527787161053273248408900649022856057556793379442534924607255616598268536428255186569163133413974964576802;
G[109]<=2560'd86660042048680007931892877167360035653590610219408801888781839470541455566530072215186891493202050526535771182328503469000137235623913785574785169198965657953772138912855960449712120749846141733254927193518388407496012896947179628370234422669510361514178400579162703788940705286130801676298969509223236336847741999000163857317101768886140422389830559597136122457008639837160443934779853530137629836952005045198492666000392972738611740322960762387517230017218372805588431735696918271539267615503864178745721401607153120632386538856886345165992421141223015367955287607552600250679022664702166413688637731381294383336787141054637561676640577697201927562794878536578717713920298167668901896017062109286309047986737412120546095049400008232282265371596365099094710878013104674;
G[110]<=2560'd86660042054985355860247144599026105825449969542042632900029040998767072996059537952825393853687438563572255287907575485204458632165722500920842950802891374851772188166789829351591980014605638761421073032903080545541221407846875526056032049725738737927244409384568671261920670145435585640240253188736583699751528880983018681111693295156334520824849539907372779097521069498167054050948896250245492345191193514781560899231580673466836999595691539932145062192460568996851347982531443843902142459934669598500083793064663776610380829334275325463263551744165133078250964085072759162453009517008301091162117295875426300036911330233099698822087795186186756620453160391018498884376066473869381327403244207714809492948438488864934676175203993466672912197177669432509622892288418338;
G[111]<=2560'd86660042054985355860247144599026105825370715169958785187485252827799513318616949843969036653445638009022658368127969488863849987060137110702632434979307481492750888855974708281754858838279804618251520675084606124895045954479128287542543038216971282259545365902713489298011898136466020442714708925480911854474090388666856504964830000319452754869868837157424790006811865061859698121088961898519431503591286158106619232335949190574690605329483988937210840765463289156612266785879394128233309721677375104951032709453067189446590770894774869595893919269174824783387669179833748744325171608616549982554356617239250560300869160768813901391099880894952423646814236614301286607185781037676231300085429339317575399960139638454523524275198108493958985982151905223976366098492826146;
G[112]<=2560'd86660042054985355860247144599367919767832843946171458095363025144077893243547024673449360351809036885693006612255235701566186274850062756499714903464555666165837152970315673862821952288076905299595613667904778301205242335603976633875723371832484063146016433785842795064582190278057390199433837457521431972145197105389225393360197865308621339260531420861479117582290387894461454079392704008343925065748675050357862400898419413197845770929883998869396431202819396210363087703912996708288475019858759358357047058089411001255276579302581779026123515133313146381135177113074954854881822027706537047037536784672099765615233140140823180083210151529521766057349722520232493200135444763853807248124338142996266980924782601585033173166891709508072445751301374857300283563555562018;
G[113]<=2560'd86660042054985355860247144599026105826643739735921427569970269842902000185521934048317661086999095032192201833219546841405520278883887019582620768009236225959138367883592383347371593894760616255043437717480859755538593623906728298910492955964469527231365793684824784097312859347236756897726447547728272808106066423339547051918635098208980300760674930792778958187749088552027071520913767598509323781076256133884950321038343820122811803400552877513319402679712834864750181794462746365575970846207888555018278017151934135962601242635468845186206442850294446029782053421695447740062537678429051960751064500906909043890120472965540885941065620181624474772108502900803553047892327363501432631159307814561002219543610517633020437984613122989523966273342738807423982462673494562;
G[114]<=2560'd86660042054985355860247144599027524486588532016285764563985693930815780328138483249004206233050550659715898373886167124141832286160382210721927056250738607463729644045743511560742508903048220714172606173248847285115053645080855632482672533320646499540818886538288242355795749940509451185564184306643254580034780634827659370031089608987902660556922222157529951372474179196628126875546238316090085579471417882279012347266908165577908824872482364654497769293718926668378041175873291619863724568460881024041910823267518732284757385798552823279366718023973528140412565421073228744886959552310450725587228736782404686131141091603058648765715883553863883339517082597420459400646491105977567570352064211946972081320874608130445212959366263933772898374987333676049591850032570914;
G[115]<=2560'd86660042054985355860247144599027524486588531940387899657751309501893366630135617390547343470120377761445114141634442734379059990044064539289717787377506791370020954896260205584371090902488264762380955303516197732110070885681407178664832855712215546060350917919679041623129491692972266705213906356968667707927035252977300629708535915536776158851839669203110519966577729673930017807822328379860242206080242104430480983589748363730236270170713604184596920866693026098577230543810151331924740847167974060675886281995349529091501703299143404520530202168657822016840752413460173096150000995212878850719847692500850713708036266777697174051157340668518253028176215393420207255945846475930001425944259374039909758376244823544846271404092035967073777436773764768041958046810907170;
G[116]<=2560'd86660041954099789006578888098933835296901794869035775644270027082613954455392817303224710228263435492372239252497955172355130544379350719027006475636466526568620350637704022331144130887686662274145434226396951093172673534404446270879603451253506579460307505189056805207656279358528748417355080339749167857661818143667432844753424608667333620700346983167693600473285858962800151628337315448495189657188748443913796555553748690556744602543788809302522703315691136075828114234997270948761866883675907824574367915254772794593608661549459276362005186383653679467419594333066437927003847171883774427195759979581140368264587794166670893335128175356958638482308304241775664293961961587381220928670097858300635297755801110751714208566491294812365774512155811706486439226703487522;
G[117]<=2560'd86660042054985355860247144599367919769106529127150244342086001252994799012313212040176904645517326300018668991249838261928952505927735771224395760515003232941548297047653415932373474608124499147973475735143570649032690355234309605787969229606851140159781672913310161434433219760216905545230988565867588860964608018171597659211825151006878270333292826235603051246289946152468047226165932311285825641096830454856317813670492288966748803204430017048331066223807330981288010569487853194440345980425113551846700366199056171099088884822708579879692824125872664749636503936954823881858444725873789922168573998850175725670616346123226272308584248784774969460242609663442670650418144971938727060666847252930268783594398380184908367471094754785516980922697016165737697180771295778;
G[118]<=2560'd86660042155870922713915401099481642334036776174672583319018551416281300785033322120845453309270226465453160066596391513175548324475011625645673796497836810889695522576197054892788741794835222128143187760893181968123035025762556039571244575052163527021991789300858394324569172477241044319547513957882326529721850394738191152904886245715782041882993590149462192002413637428428981514796625538456107021050150024995832448621011471989257583161997538341527297766914539021336016574319003607120220145646797882843869255930184998185200180916036050436928040023216595874049420667582241793246197422422805304752796554591009973692031937532575876078502953144306951235647094479235845393489979814518650175311554506203248932848239565914785919035998302042981440718203176011776309701738897954;
G[119]<=2560'd86660042054985355860247144692364005135182539367195325444837164972273252261691372469817044057153640167439820893706339872661740617280549667106311944414980594193860448350187273514201884819403444570890780633275883322795859333121382760445387664718666558457943456029184633292647643781847512898889272535860729031913406575399085962951373175634456856448312367540881030052220993510222913557356293923621090326233356288919628502380266659795741991037643228882748137006950057873481796904403741300662815952167686996950811515698611546738302997171491802678017953343756565290985327707162190775807992225616356909405387991903514379920476386843087074926648297798580189995610895322411076474298398610925820805994371244181063032357106511764672750501310567478284587630167951433109767227692950050;
G[120]<=2560'd86660042054985355860247144604837025973196573356997563505555995059054939655459262649553745598831829568815277855397816544853095509416692489340062557487657352795028502477719666141954325284289825104303939820350239211206257681497981396223654889801442790898054577111210148902036456581949690801315309597925973795972818018983383339561155985028735182783822906579365585953835428793794644316486848410797909351105048266540062450073280243625015858982726015525328202907228094203150188328101427052380964895199495358952500124174313925564789822835444744391046476300038085081704737390767567132639569571910351441392237238605524455157943599693080798386848947172293316915646525751810722467869000881259724222195758772312373404184501758458775902260990952067292652138367008552056165117116686882;
G[121]<=2560'd113741305298053846421710712008767970354745252404148715328724415064242331614472287194116343533969700289096027230559528469149699554797668871602668277050004692586659637119633323923913104868157245633923963926395585119284553876542601337829353807167593140858965326538523587290223695877601920824970736218146014986893074729774893458663231752165467044494590882104266211146289676383903601937870102914352411642778456664079711765794502648165374758050398902335948105012104363108382681111463441044968080785449707312022361222496758784110446591736045021100967454427516735975940070774558331598679419026020224851561316474340455563919418983211555891526251498301729623951495103907103479966641181020661147884977181142160498176036955168184514459219681548845057620095849993290770917148695077410;
G[122]<=2560'd86660042061290703788601410636115491441695476270755969252378915257856653451976972113415319561529066905838571460457347265081034390201220655212173602862834683160113290360097209085955071294266057458932308982146310517199981441961929512779565312477989876227220098137125495487715490323954349907881287271635805469695503205226302911087158240264608616069376871267984017044465891003704237086725238095924078186527011552052644807351446727613218254227440472572387346737444698387063056542531425887045565206935235251741113363022636705523631022726226541431865455489884075355638866559611977044844974175911792161110749790574640526205765794680537423869633984135615236130660214126718758663205850933437104776995797916059590122989079827415510065044796314882963574513446247468675821236226499106;
G[123]<=2560'd59578778919107780082274201744615140160397745172935098203477919818923773953242782976623279258701979343768690115810812085746252791997164132388125526186779552262369312319257174289758137460348890681451681460955083097770147474257417425356025183691664637633085303598279517098726502698156505088320621480214538595982808944386012260854218781747590395561568311737102566462926326650216614260718458292204319399015355833117400409031196763806723825526636459393128787900536479841698414827049111518095635280593750729754219035279817809417491299681530561482036396026916917833841027027073794130515834337237042504564561311804425862904728167159447458518711203348652062992155598532312010724537809142586060849468819166521053567407645815063447390755822749610553033815010850298792864882670838306;
G[124]<=2560'd86772853203811229389245804881130417010254597758788168857200471096070390314800883340225316918822798947746347097220297314828869191408941793082022345259215277952079414153396286495222524283284728145265147281897431930338871540673741831370017256246362922932422981755389124879145874738843831916972943542586411246631862222196266219432306749666134087286424009862219602628367944637451943512405894761028094244961339666761607817225623271115776182533331900889770928963277835053808222028905479115329040388454943053524944432082425475679390220339404543166149480145323384211072335638783123297155401016651642992317761924518566895376915103867076264689408407953119439153009639821777428016539331711031053604917547479080880539801453526034441946945897426008666626292905790328026746150224798242;
G[125]<=2560'd115433884244440279176937170400711191292356436975518537097881303842390378790409998643517129098388973155256510335016879380647050606856756765720848911674684054150323434897489794670760665391277158602714941753015345634602982401952630386307537774198923942593259242840533039116840001333871331191856196538414014994304869048490457933371719123108295037190284648314329534429483337029594426024667051607903736596789801902350551651942745657911173803641822362601934660092059218976345614678689780866078844526118301851294372802825975431394384510396611235952637159813865738013960573397490894246123287241866579149424621121261208684312362362663160649250500802399865151479999128315337393853047617986496981917891123487082346203092337891113711449687672489593104517604119043682982172216451539490;
G[126]<=2560'd113741305197168279967359731916973413779272986003492927569896550740855482233812019528424827075622775610627851703025298144945068876407012248025808241980366279615944945617629855812170409669093839708884499870834994382676743210436662037520526338255085354363405868788596931428270585739746284556382511524379399509244718871352857235511288433807758515121888255614272860302903658215219253262896657603363159615288181934034132093387283553548770628678457632495345340235650230401495022252418643003224470815184347139077620065321837851943850926849454805815985434837997664452013201714062739625251900050270846503472323544813236649119420296512747207717687977118714725354886407337202825318481530526710719469681929557883124417394910130111087245668954961859549301874279537412200652037196751394;
G[127]<=2560'd86660482723141475309297140233402764849692836794158596186454115562150212685474971031912421787266663386950366732321538638630257769609627608015294412688120031701120034078707920893616087423798130862153958782341505432162885169250074828622206170083854900732324754875389598212084646792231308449813508682673396390748010550854804148082585111119449762875760228650391513726903299737148156639682133456985992087183292323007132370951955452951710585589038591407523822744622947652613961892973314465715796097064015714829547757099240136924315123495707676917362491285392673590704803249183762801688828181762326088986153493229194896840890463418013193946967295886138375931331463820086115688278540616536491498941953042259646507306220794268836403940781381792371709259396364459358889629540557346;
G[128]<=2560'd115433911691621446906621395344017774961608208765451948053988993542650720250031613364401252964871524442026342088693393035769071569242367343578106295586235676889843881374348681781564057982459406761779600439617628914904761416378132256935577688786411232409205294132588705820970248554102715505741044716572170166676624021605965909385058155489092254929566485546898139591242406065247266458449458763966424003700964792845753058184305456126091522180902349113961366758117778784239144470616150499364602789405338374118255948969260192924527777963823239282757345998535075058488483284034201054714739694338948843999334221524307627167772792372906767144330067493914141259296332069663754758245901298865406619233261725011878112607591686573951605150462756202402559805579234939802419734390120994;
G[129]<=2560'd86667092752207329484268638659699181250365130447820249983240489235938442052831601787983170352992237439836281018561242354846613385475545235504291821715352063122794224334257840738706457750233346302420122211054916083966887150171054697675424597500969651227941423855771768723154740040800290464006899810167422050277862484334478863226749798903525149159890752170683523375631149738953204817151606216150861582741416996261565299059815460614861367487794579722218086775824748002791772668651553778609550561757776760076640485407908212854085597976304638770419339010486342981305196226627951500875695427539080828687979308342679784535099462324506166414027631491267596360718405080808516165227731494249102768164153839924835540441475120656765499550547619882384737702346095881907666912326853154;
G[130]<=2560'd86772880651411118042259351832475164532032683832564565061173956304049869666511996078968543581134623465552832493001978093005390270560322586470451359310195249263172250582204868804701001371970468172891981426705690516066218060322139556458531670334158838000433741854986962436935200216767112597972921293183002961395743636452976506026980830718629412992011730618645807106734829039927435705033464632686320292804049929222549097652634924775763582689208856616071612836847145388775024346518124498072990781797024133432066585619675932761487288163380762642222172384276830197285667251854382803112546460433596729429686748048661943945763371192450535851817184164271777988513861430259552463610262736984709733738568740384777589484674837524266300678282802013798352334242254644108420304729154082;
G[131]<=2560'd115546722739980474480329526132057506326277188345202266293755563842614159020927418680845197180062235791576021463593660129469011825514441245747089045666831211795960504335549507766243687520403245963576653544956609720926634598360970211122331501928646137652111217839191671267080543628065778200394950378389071850839575328682537111388413421185695724670482829414605879050867715204622891582489057247351695482059784898475748030614464427667306359894568426382746677688112783654775417653766583321056503391116819219280675168650242571582913234640538358988182090954304055144867991012468518145079815979493146203720798819422948516628292656580594363313728024326604355419072318257622206048932748429706017416535341741934653080673367759515394200981211271722801369122577493037209155624105026082;
G[132]<=2560'd115546722840866041333997782632127078337649813967881559016773917877172545129559538400798818464379668576302661976516942306887767255159740657362400006406752161676358929933714450591660537091731539178817187021354497217260589605031265792445370006549610426756707469627246754091542081044312786293729645214925485686744949978415725257788770678217772773498950120966008653418527439917151797356158777889879121812486266188723249314833929041956330968301653842981966226173116298613113463952802367001954201722720855248471136159923051720904736768362648632308698262234803096274547531889256026888368694665846988146003530557398107652974765966318390520739252724813206918563476554650769668811584980222714646524558156297397302405539673745925195412868312734643717129648379455373060604512713187874;
G[133]<=2560'd117351699614610380288105473133013189704692727879975928932222075548945054987405629429136505774746338813056740161810019409871451359444624269190030622841573473994408515580004065317066159093295121006714438356789683402104803335366031064758180726473368066568444401761163577988965137727960206632933460183916592604449402275538647672487240957292070276152299457615914370501891211066229076429493458994393050821527857657209681790520307122023835358565780137390934776702556808396708358832922520325392585623776998494330264889350711077984951248442161603061622296773178961564548224294917518988824812475400671858893181540012511869083357637302587370108326113180403223092810130390425925080953210741849778358802893380376433240628983187632886434175917923653422861457772203163917654457948713506;
G[134]<=2560'd117352140276485679448040733356479861990426169536341598417618089476803698312274472108315541076051599581071171979968801940535183886808921791274480844008146703941978261152120235079846892882849952995429204175860118508455469948999936388350138819466063198268842250217370630383510282827238019705584060836429994359389096370141332769470159339326782914799993614251068421652879874344714854444338965353174802782566946849361829803626410338958040194302572562832902749697870609171826878614123976630867756911130494439689447998774678105550468204744179247204754364712622413027524340277922181804355880278238283335382771488042702166334777600502811498477797057411676855673234210913043627388294444652409610197423088155122053262794076442771685714984584442347312115024328639214054105621723226658;
G[135]<=2560'd115546724455455467521240720710147800655802196337676080328353206644191505466327218465292872810270508441029784160794638820969080852602877580923045270127255394613301755484311866723554696374622863923442264187057695011698286253892656056665536029939086349010191250566925309910022475789088755076343184091991088911081378924299810069586132289976111124981834114783571751899892802698469284828771524554937245118168217406821491564557615224658983120697708266968305168915525210490429943877826782489908108396319860995890810591972454299079645872055500695623566425706571022481689071865446262062857938829353348834178717790000782353888672653087321119261018405788922419387545188305557605496731993706447018690588204122841681295646005561875357572195776740975523265705178156756596446807279673890;
G[136]<=2560'd142628013430228503557081281218266479248212585769069144996683399245633662009596153772531916030154576050128715012382456842804735875577673674647149933444654388113354839339139602023687371982197939371199692097807650005123145747004004517161280097320387272558661224857750406343579106230107996745111220541296640508292004224008323160059589542606909462286967157117787201018125083934675997892051208732559938985109693359661822947860225571866937791727847720462857313390376491469228979688916558800366996940940041135414543890393789379379966242121555458530947618412308587318639494004996561259067052364607422023200924788975499021425647457784724348425777532187566093398822154305703844025217124042433252892525901662212779663543573936083099188802566226906654570203425719446124392000279159330;
G[137]<=2560'd142635038193554435080293935748684852685847368530203091056651966548940930371522730987522414312495251543955545980189530084710889258158098186243101934465013747983003364790447873387171773742648055933569980590461910492750556206941039327256712154666548845145759980239390569297427810037669098969129737377283362117480836753025514747428480371310242110307824603619230550145513333629118307423111640475319872035848943357384870893575627435436996299676683331238898043009918149744751003849227640833649163710448087805604974936095031511705213285632113165169763809048567542174404129447983755415975363259421935564022864018240503855095642401847085030314201446357075797900724272206727264968236092442285892589058590597386995366132330093160190085026290389888811059833445338308552656129227891234;
G[138]<=2560'd115553775051371517763048858957117660329690701752383389290083229214383843940670454416209368991877340973677102966579354923785116915690634065938696359541695609614053679807310959049691159235641335581081516482014820772295013425867742164125207122599747794282909184287520215583740993401366738901779501873703511149006307482413402106486008199178220130565032900379045038303019257279005814742000938934449341493750956569507301859779978346245520678026998739959749471741813863161264782904889133880132317154404787779167225716681502040734360580893992226465847674301206701209168537805800085148894748476662525924092983677301665216596238911694991845835915416651995443142724016700790055277810425065300988725616754988868343812156051437783329559285346994116855742517059496953850404729444770338;
G[139]<=2560'd142628013430254769472969110277928960657550910781411454645039951286106835109283106402469208982902919445754651827411248917198645566871629913884413988758740147722341170277961446331826121508737146806256666969088445203328897580932315784610115090570871824948192283375904537155509869995879153717881545989864945220983051313025586932921515338106175431146823539198494939542561743896561461289872648478478668557234321798261431005339514515641121863736922557685077166312179289876883858178663698574484247514787791748971183610736670009785049317862917820694878678125647977169299206250904107495977412376361554884174283801445368347036386253221614234959387141138220818111402541967389739678988914251763595084670168928855069132786403424727479790915921023487145171388779644260979670825169986082;
G[140]<=2560'd142627987603943738780099954543001557318226344960567346187235201862915381733807021941129528526297681605008410310971896306709923603008144289579932726074624877094322157815495792637110223994870840106107717000684795023636685299938423635826476073953993240725659643662708844197250824230861065775916338202709556162270971450966628582725558755653684853976322460246565384245835479017993025945287579423660793460056141766315847264154235417713825088079776740716189768167485310783076603786798438895972345934197024174768606278065854435195540952023472369719500081956490525275051722801899978451524056539760352323009975839387132729393564500236721527030227165175374804780111977621792256588868585050412050997080671858416190375072061896989049803551771976912763055476231702277591011036907053602;
G[141]<=2560'd115659148109124404037260598551147118601660598798483816134459947692508200326127097906668682319332541041387484196040097036121904001914479629116902993191775129330855201056774544065991921708423220504325278042099440735385595664592917688580456513388967881893713270907456891585637433577300365244146840720679577774504185407995048945599106167271307022024311863292763891084087795541677893010430751618665319508549552857105357902449992028539209428827396575003971729081626415891459451989985781575081270324215447883680474784142604034815695903331100628763360040474474597064828522832032598767019332075960156749551622151270457479142553031667607736260604084098413001857410811319419279776999155234226714278057952815800907823159049271852117699860290262864668334677585660431231110525550207522;
G[142]<=2560'd142740411245001979815233565212556027300465553640055745462782506843734964415186668376160815387863343418996413166431124869196622947314954016579837333787927166508124849341924668407599581220724197724023885593880850453100037898326815409020893954430923208104974045849916021825548143337023452015414703737642266451859670066509774153437402010568519732997659313285250746247174718040331185894760221857675531183179175502279158795175781148356802050683265159799988300125006053538116642348949330715867594291780169046815739132599489056171153243865915250247337883716998698114173847200663739410836294503894916581211045945091008790415431952997657112608333402257216246718333230017271743426190831908513758712201625203197364911572643296273831965553756169996610573221166072427095322518718915106;
G[143]<=2560'd142627987597638295391428446438176309383278691266693932275307565595716775136285768568741656110877034396084807908772510960130722768598234674215845331095969161552454130315744264760991676535610767522951783300212116686524003308133854499104828556563596912031169447347891561831504608052647423658701319451788346577918566359423336681542342034811663295019312863543876568834878374961397125066250512290896270307435573271362574724475747347813315368087864605989176192644892484177495857529157266394812677937399756628172094548028128388618840513943535913515530164252978228951480285133378589137627423250364552286622276006948445145839834298748959730445752932177105625909258912474927993237231921030251543341029987137603724660585331185986211462511189959966852396338048909061508025225538839074;
G[144]<=2560'd115546722847567115525661377850616914447663394563205472629566092856299003202915213009757342730339919271177687263183000497937250624568849295917183811229700509152715928629853557839167999028869986508737944555430973443121632877605046029980268921999267336237824541655979308609370347905517048157395015933999250207324863165408496718794754605248066229821203350160693794617157702057052602386195312301300928101708307801435910159336337561750032274812433220864413900293202934289840531027115250766702237631645906479367556583140316263875701824548671152854896747839279929259148648195153754777977395407714506278144582173596293752627354067025942025169123632066457295638342645085187549398308883636717166896366559512895849896271987832022931640371416237395358607173718835255609002577776227106;
G[145]<=2560'd144432964370988645936159619263482075605760031238280361861418489931734852553236449532135629081054743224715288152824884696475471025700104903823109319768893938684659427217211739444673980624638028490846764708572083568051553465974529923877002921719506562168009036555845340473344530211886005933180960297465594637089537575038594914653794479802340639834699253501476544695349613552527700085163875107753768048139083766380086130712356710640207537361960538249761135780687649357426737420161181660823928405107859413305531022296726611956163059176250763426322526554544745991920033014969886585757788959009809774584937996151143775843125885229017446224847505452002108410435993909804378218237498675472396237755514439162655853782068390420398331391513166507349515584113804524386569125288358690;
G[146]<=2560'd142627985888889102667148982273700462262924626197768430604900726135317488750968787611644443538881067636467688672046236397284922794569128138138528833043461479873888628375716529170742651963184267613939868209741942167674524110576038800352168942556479446777977832806498623004115814094054675359093416855151052817523869107272045804992893528486569841664767923154942481599879629827721336490908424463408319704465532803489722872638113711774995787499672642974628554464607847172543513423838978047665723126669143413621464474192912826376635617836234971399975416222838142676167328833867432106558111672636290126818425003693412015378026302880040071808069875785541202643457722696644175901805301228701704068075153678579535285442486586966397814238011475839134239358413230031924896210438201890;
G[147]<=2560'd115546722740400831010446310305944279254712553084346319214516267948232084959092997415696405733798435090907681704829284539214124160690450380250840407037892905608644569992501082650269571136101706010243523546897573036014513036226951616744795705854807621837236088159902874976416218794284556544107089764666053265445900033516409903615592146712406084248387962754011667702141118550566038865332562031838417636669667468621849160744647065566320340982122654148271971732787716540158447355968891674314768810845116813949774771898333999151395537925500675396523785086284363405100309478898929151095334030453332628208640242351749467028022704907771259814196349714782032463224240767961848367849327121428755488758523832075800727896884949386101282311395437793587903265790213664903257482593509923;
G[148]<=2560'd142627985882165040180857182943417696795404570648039823193039361563476295469117443158015965380570117786922091451964078313216705624027017057434102556528493999935530264173928891627038446436224898131306422280989380617028638091787270609610660868701040669620638628288627723365047875445084830562662658324496110665229551476398507595427626740266675649947849538742934195359690124450666715123000031210060170582902610821187361064292325189243423670055085585305583640601446876236798340845553996462346072614826299817860765579212854302806396950096333700996737733549066875057239999655661214488400999294561032346215634513780840923726015477368160736197853618780935557504107397647347094246316696374631720143879162643325545170954333751869279998476821955834628592354598376361783104145626178083;
G[149]<=2560'd142627985882165040179389104726797379573142758223675460181216702640107990090019787053360370948824196462846226945482515589157747772761876442398644189793869841064509865668507169576714796987654634815609092504922428178341527166850025139266334746159830405982810652065557306506486849569543116606659385081364252824116836575450455057324989401497587360339793803750829022513325685717399757769088664700258743955858851306862242368317885751106804410205992483058064136615534973961291152764329925777800729852496260068430145295529293674263848953573122177344916299587301356879482706167439967280362374443968444971336063227810251141094300763334685075111301255920350819152287440183063197862984884068186974973199726292693997547765604416353228485545524959945116455643894430927138026128539853347;
G[150]<=2560'd115546722739980474480427398013142828912679700492409715812931261214948687077476643410764615230881982208593579657478746189027867219490500397220981367124154655011105765173675197860632932595275939703306852949408934772258347804142784675424528495396861015625418462501559871215969389752361720199645796945084263969184692082567330985343380920153382471235904209730191341545355672631258588375167942385528937866358323842615882222426878489203382988312368936524725006711934646866232444380187442498176807141950215055327608829563488314564328834332596950792853650551175499408734029805898650172956784794318634859592676893263040084603138113283102277627351431176584255104655705176076682816785399684783815585760170384354682521744726073193993643652165869551423253819797807134295414275965133346;
G[151]<=2560'd115546722739980474480427397925638548308531439652549040366519478438834654444868392246416125294134944568058844212684724674525317405057630843853801692572657109569163962786637903340877505940433495603772752233046499028124746237022261328771305857933499832301001238386157593578917598001795739769838315884829403466346818846425781504141914206877417906853881083817949483590952866004639116819241422616032322576302203264190127196374889118006248413310871791582932685077064651798464149525172016815730934698663578493576336430119429469731413567799433803450780773902760145439566669468145179987284415014164798252440904001188634582414093542886428763769984928784503072535871193430703404078558466630145146978900113389338925347033391825897796556240458398237430907868017722398331885312612119074;
G[152]<=2560'd115539697882470037139474402743857410363892584359472314316925722115474212464212956018675945793864505184351152348820092921116865287662510504869064898697120625595469656923628676008856603383082780377639670828081901515972189579566054128536088358363732501728933553953215039843749033008262015764805676174939070891321687478961597517097828402155446146088311242145095299689564326776687624644506047406997520117992636652354334902977413952629059979213002726618982912026570124105164809431916959867590408794843917778161495702955918809664183115074078097835686477871863722972918601415269362884031189673331065147540018674678903092098672346306772893202798895846612751362590150196394259281176787621678711320926572102828496394178138392589933612947304314012218109097421056334970022856835080755;
G[153]<=2560'd88465459496493269409467143777781201790675810000144956849697205763661158676198350590498215134406858912178694433706536602277619284045209577850705170245573010748411411819408981189670590744238284451838403179418350355793914558559133070215999067848110197504582427484396748830210894048467927317147832412439146969024218925514340501143454363608163866742778123323894566649134312662156282375281662767631091228489661784914567510218391531497885474741912760117939676866516453045498422053895062256841539183754861433566447476599375017183023646059021009606517872223311701148622887858905780525441189315543030972003824236147796504075461044923713711607955600950384493215044258550372112404355435994301884377379794659389459086770974546165942728392398779883964812996339560881420574310098215458;
G[154]<=2560'd88465457882742914260173878620787944279274701902757956531911908073015477766881407593834260047377701477821415921048801958768908135575123796054242911198818241250330346178840822909446718181221875621464785538165299937549956601258266958763210729809379616243938118868697267008735755336865881808074073721347337606442723863572091811883084903969642469118352895644550741226358756580381908778422454127406091572891722436209524731834072768694301205017085338589646792536429370659114956096785313702537505295201808617069413300407167471432804864589996627703331344973342438671140856135585829548690448301507954606609355634531610389118638558201339197031109087665736616493450507344588416942983524094301251021429765874479596665546731966310642984512358761039120698882321765735814291691475771938;
G[155]<=2560'd115539697869883971922470567459517591622676940120312734509133384505303627294176414755425821157340427063879939193515370356166551383295220986624702991731492700197619425122582726063177158314817716302464870412103125648503486767647575119229660193295016000641380688172116868280218437990264069542586246787609045845021668688017893638813378065873996236010101078034776825009755620475925388050917646227716402796240547937646793043049918940163229884474564808333471484558323565697921014150669020618091497688638781037773655972964540009608080690841032329929254327289329937789599979896944438366323955250194753532803051705543321007021028497211562372113990769591494449838052431028313653010529902736563180494322300492170493957332579094521856703477215074810220636914634853327814093001294230323;
G[156]<=2560'd115539672042784773137874761808964209036897237077708390621441006648531858062773345472071859475079106971214627266123801224326743296295339291291993094586476767844785918665213984925945966520354105332350977146993336794645844783755569770688320396051070659586013743544663356992339406605149787585463246065115038318126670173755430830175338373939359511286686641696280837984733319755298612529969974724608347439833555413493721898684441496056195405974396430279594730568032412020654950334064337990013877528281127212258871283428415720867764577075655341858255751676906564740745308974909852159415926802775548040493909609747247368859910966262199912537380495969503598637974848607044403389649047650442953573698098846350383948866898587761089036944021085820662792145917966310214245322162647859;
G[157]<=2560'd115539697768998404670953114254977546069019197573880392485487884831846386064133347215039807707789198675842711996192754104001108794157534162564245418387072206921733292221617240926421756753730069659295266630148174755317343961684345522030513389897437259754880838334595638910510174629379022025263015950124804793360346302156659072440245356288247567105629656729184310780924002951762903981330638116181396542365640309249632700054634255685573345302992556099541101647503254399741605553600221031436521725396113195454135840641158937098821748599953141798638674108938596578615562578105679587300972653025799816708110994397221461540823517516487535429498268722424141120135166999705394678146008533848662274050723469364302973916057176603508244094815693453916315058282048083443282906849686322;
G[158]<=2560'd88458433018927122954226456252437156804967733885708061617607989569679458651499469861605752207716654612074528032077696707197882444283678031036094603340129412790421900238963360569081849792821571325863426234297496563973563981427236315199592275250058431506457877812537897719733478456005415315413820541948004080522106663275875725637469271777814573321589956321024457520553402812649631793768361487592483608608135745737354824244251972512148882928057293039038625744021407929847031298646352185568240751981990349338825421615511632072875175539927149867226388152509025881940827335099449134912210494900465426987765745353599159779230295354886684922299496224413896145561168688946439396277738267282440775311309592962433274126020015907839751022903194907174510095203814047568884963980030498;
G[159]<=2560'd115539697869463718019927466226268559405427677260419490029380233834677904170548738085168391858513504400504040853268418373669706543551198986492072276045440197063363383653965425764653000479605622325102823743053156778149036854596443648423796466399786027285746165372874146028458999646590726453877475409909306692482632572888239882555005580266277695159404230026754958553655129446851483944925713149136610148681846446272466703465022614340516499602694219430850324481009568740581583192384238353461372459863669139694241022384289829524100767072262536204755100170581636038304964836461768339684018443564538361502809054970613872717921889953361047214993166759133389792620106584986163712380068075029980923349768929538887764924644950566447878363960383276736891880515381558844058702030517043;
G[160]<=2560'd115546283679267829273206224454734348026439054486359117310285370833797594765700121225993030452593724296146801407664025558103210205963343817232383049428970087595597361889163279902268996067026852040018527893173232656797795331983377699383498924641282970354858092792257747960633416068773964851356713405629376627719760964865199035726622980597758480065452714818391666417643552171803946526500062553281830910666939024893929062977819133648141728574321882353646761652449391114235023829209218703212873108006931415201111086978163916317480178986740358452695354058681469066300286714289245665467041960871708640255145007595877829730461304337329087330671046212691518098521314612008291045665616110729189445259046271563712032974150199510286017325474018211055298682773416693842692681917211187;
G[161]<=2560'd88465432049312101679788652114917014341211474172827402852381276595888026718132566037135344582987074675928783412487339144758347654888120538258203969008373183970397042496673783562652515245597219644803400738725280769884338573630169574274259990755377423263401075534618645338664002558506442109226393568687206799260137193788587305110784980714011253486696788663257683349188550115547245078869953800105893193211240152022903871094643259295788783348251742356197236070759982756623698452348775320567771957345047112426445992548447422547393259246626593332919864300363640645372054581505677631631076737931712404525068077387559876887460960686646855081380339784509805873520852787898065937231317062104188211983626242243470707335019051304454514563087255581804848432080125080413283517159645731;
G[162]<=2560'd86772853103319753193665341698920771143646097995210854081609920496850576303964698753463797321347130400089286477798859057879915915162974693866399961612166210431982382448492300423442847953219572936991714719948408326360539523856216184799749291885592308792804113988815759235105897077112628718189120581785739439148718328341847513209400000605199651920327162031439244989446303681184104089055260087782871875382381498069359541734411066662459329884362274504732792322818931281350288673865444377269110275435338500991800257980741021549457594839540096141100953343704338138038397113689869220557470490195102139378969606685740363606953233279342784624714670640256648738598700208738834001310556400350896357780790614213034595864117741991451102661434780084168112548868250170485147647578677794;
G[163]<=2560'd113747916941287236877044712028095155134553165255421917791512490193721903066041546275285772485943073460696619647771077557934195970507491770429715897732674644762524387898043628507376892768358503450971389421505017670000233708131615821690373672595191057460405698517947139948397608930713741693315778035692397922109529300971681705946765585909495568913141132581061811111669696369275711053376674408849566453433878008173626230264461486500483257046350993143529690519619416203529493559529712323745060721006723432103647922188737891162688795966830080741293515895212042421395746759008513654433866004587520284994917093999861780997073167706166446695674809762473924317839292261620094378548308708634963211280785344878593429696538564691797973447401880796824393045721253792965124183197688354;
G[164]<=2560'd113741305298474202549390532644703535508520675597197388581992123755693495439564091757325968027575911698946383024094649605455130669485614141882945250210553314870279233633153747823780717001515428513380065333603171527612596859726313335130972442958390891452349946069407632087295670558744987043495979832276053479318158718223192776421865407762691696184740832704136460583781312796190390487446963598438353785010717848686356141922782284802871131539976675178786517770357566880832115162142264593120210003246373757780104893328321864752431322814651935815247759398740924919165238255884172974392161519235268869238882662290866541386105322476024646798814523173208804315723710379404446231225315472063284324414798755085852833538051559555970842152277361516594611081950398013999613642994299426;
G[165]<=2560'd113748330061379790699678668912592370520551954942963963620568066779549324889995961998248955937423387200042396312630755284089459113811570441060832596364577960326885132197130017628217530475162913104889277541002532228328121632323488618047213115236083788471931104161785070213054106178472743104801586043680117539382362958103165177729701831242341757435272749522899168807886354055416579528832792688588671739041372970974240535005917589287680949583479710052763905042877880414908386503771898177335281550842042724163706349429453501771166585337744160017168526827641335244563574022064446707146786534709470958585937745393043683769044026006865859213319567332977364912694174684039683703826458660319972687801630550224581232857053654606888681549535208674112432131169622981774049768588325410;
G[166]<=2560'd86667092745900442164330280849212761457465197622871059630889194229704232285412190961604724441971690923994687949458768164078916018886077163712851268702903371622646789253796428714126738898117669970712936242414798511338233374598068315063022859289347180865940676955929806736923737856284810350768529399193076583757061590757728898528927385893216253608698094122890742699748587805528038018264876503884874724493594533045902166618623670926180216743112922270279415908098895041647030424172665846880073535708391873493432104952231372103290105168489920419058997781007910624370086650801251818808705068493969156322522581379642684666641457775382154850822624160647886984073252054347790364932351024137498706080687646853349394110658392932304085211621520340734105787624278855708183175077442338;
G[167]<=2560'd113748355988944199832880788635764573141166607235125770080410534780230645040835505330814449972561918941582820266066878229412090900881147825006819366956368761870053939028807600363596639464353225844757550611788795322843301080722584576619475659769649687771556529064121448355108421994755486094223338250711500855730092419235661857784664603017594200373317135301793200926557097322976337695539058060256965818035123346521510059816006398427927133691356999853974118328642521563655898020487401423128705784857919716115339114709060507994257954189400322690001234143798748145219346167082065750193588021744418132386677254567873276907852159715376979894396481266391657462757938076501248395954519952018992879992790112913102298594678414488014714792104055625319595477778158185190324494305211186;
G[168]<=2560'd88458408906882464469919517012277125873628432622376187574896468955683033195471860297036492009812829570618546726448327320228057763830192741746015142293620198615496523232830917612800937229130642373642157633146562893280618143802598775675673261854348809180887662247708053324898793273919658344913119604954194111640443321312894094452738432236813205010389179614298399796415634554786170174702926617030051048893430059717936936756044748773618151245736931016051124960357571533046960575153645361955213131838286220408762136828279121891980614374328170730915052895351475950806533644377530134342724323124443048994088657738308765824479812372340975550430354462598314173594254773469329910906752684662143043960295407056631002531107296627864480079335427769605953164309855279624467057896272418;
G[169]<=2560'd88465457876017210180558739298088390231195385908864625869265837285188960442730854717686879496023312052215202777526170588552031977144647656065273295976445286819052572413049974723831636134182625945664319370632625531182853790786823272936194890062525271741060393799737025417054513546256233577350276603443814331112038483906093984118947246305543381449311453037901861856098847948560146107693226311911963006680803910701978752556002618560450597435594312431258762843717607939153687776414589444238729810255298865701772650432833000734426813196907396135113390662383220743683212876538376706271545420281791518803002303791682367293247729404250794600150345539408642268815991215057614422847751405106218930605399963152857161881355573237934348899116158230412050752724911676138102494239863603;
G[170]<=2560'd88359671691894227793319936367956630219424522166507737352194292646464006921697194167561539910344179867867370658219073850587389302724263575503997067125210522646966996189472083877146969912374797957975606862822731290482855422109355003339381061219331073972614197163469028950744046897654948515442103629801326695773984946399833149966051980437394026558375310117759861673613846405299976623308887208310031405470245211980611894509377837838309305597076092904172703809595931638102973117681852250469694215851597518623051395065387474005739885366598507464749310670262080692562500694934899139217398859947235910857420556860570813971396370516765971044578715172437022423612553760070499650809654408358098648353925527790428086895104370139051382103962853173125234271756029255529681255703650867;
G[171]<=2560'd113741718431175714024118447237919878448438926654456852798750482116454039604494956403869678844454602291509214156950041730387188853092110253544493856996440869991953613933971262432670862130162610267696590963394408729072610742216307834571769395183441869664673819550161727467831050402302423164140458998282127764366391496699270505898953418072636753765712908324393783260521181389626157539321193720250349757999846000265554856618696068187277881772903924859955351896864639431743555266289535607435701756243016392842100668203995230359642914654161814633204706260106494455308250062206356639958327795132596712315357110360342639167230315771393800581154160719217547312060043895607439012934697668468983407577032718575551023883399563761666053732652665287924972585230516369031608530017395234;
G[172]<=2560'd113741718531667196630705111224937734169333510256369231716623844622243274539376466100086609835864524286225438783119839123498442097596378014295408438960405443477241030538221731699727232371904400235493296131833446482225746528365909444719147279778057911738785247273207923693069449513720856090888296691735617051727854575254416158316575618170017652103780462856155754405360342652320163072122224680135636699041435440028316707046764117748726257181371038320734527661264308591892171286097131570361826574428637815920465920162815081932694704131891988430930842744562672903125011282686589807529211708686767383907563291040888067363895507374886165269582012253539852956722488871003455398061446850914517731261129980908675456970404035541544890195186373393935741279433090363240029938892616482;
G[173]<=2560'd86660481209857870253996095267493893809253665099487406148372942674193345378274131737568658881282684997841936494483420797161729900682270769819997937463165035682258619730506105324464585358802935598649240482443501448948575706008554897488150503439178628617623340372880420141241894076846450180979548449615392639795598738566074140463829573548162394452227940317963649126098685337222890620914285162773977079732629696966815921761225301516524820572443862069708470184450493632193302786010442122908978726497873338136005803573882872535467024464070992001598421619535758986894906735811567233114508301828478395339157828731164607552772492464938197332934580835761955788048989553450978264218545665712953740053983859674798105925189884166598918413950991496345762472038043153541234364924506931;
G[174]<=2560'd88465457983208130975830019325293843907760885196073998519347835790111974868927871214788320175929075743223376392095244945858858245365206860640069725382287311158839855558533735732400434507302440955275153402358439236029495370770695715885004502119826227345085631016711623370338334159733960414857231941680020847100695704388082052053122388600313195783960155846796446748342656960297749531707891780748595254758414790931057074163332984541713307779066090349255793866407385986583911431110002943188331333972761299264731644797779238707502821363864058097965670420947000410207821515250834219868712916235147887339030101962329402390860894062251477167478561089879467908368312089962085661534873544067178847667126969428682036362410368848483651535219389945903492917995578202449640760498402099;
G[175]<=2560'd88458433119418611951351097976452979021159067532142428305848460098302049925250171772866193195159698843035603345553378223080467119797086677617741976507946191378772464929980870905126371891476932428962437977182210104798996674291142985361395315932343746254162095335836012670494931254965561577446252703122208562871977208388427240184805216967151511552394320809102053046393106549318717239883844147101509886604884357652300856366090017480146183437586238258974771878737709738724531674085998339491150777459926438393750878632237369240259280069404212828825828500637579118863196222184552008621594532859425285997097900093675927761874467632758474196378120842397587650404961302965422057259113757278326315838923653659850548471239386492788719375961680534770992213772452165304095885237629747;
G[176]<=2560'd86765855787593793732341937595432799895471165791851582760673985455518053998346506734352370048600054707413123603367969821685458557509741694481517599240136451985684252910788339976059482952343591057860970365095175271569101997052865081465667553432739611906001577146734140000661494832324869128715029942879446374870510265464573148820015466734473675122066915816030215000092070435864966498875652595383585000799220011964641944427681300049828082397510872609544029343690945031241807584218512467886577585841535091869491925457791656659524441332760905014858735394028400491838328010346215991238089805591212969382060559633930097107388193949186039356367712674535206312604978863056287423074935831067957573968413113188767711694898808762711185968575607174456307534351568401778612345739883043;
G[177]<=2560'd115539697876163150195363348572102292445163693093528473837794199984876596896203438895259779062167117546436769739480899986052176435955322691293544009974107743411364920178330248122727086135447495451101514475578049492318875148861138513888509132910837138363285027513196180154953388188880966136050441313564815192432321953364039373473152612046897284454258305520028558686589177954967362847391796411861826729247294083043204159563688533238236395052272563982193794357930010472755166386444141530569682210808925710639952726823892511505773944580928123675045058462954992935312501967232000850041931622330159842236451375990378870148567895989492549092369222929444001064091210686442170706796864653502262086413596031619193692833862368696357900272560102484773811194533667552182423085661762355;
G[178]<=2560'd115539697876189319852292911707030498766353879114962661027504560591298123073018209909085345367518415736585000112592540752818348124075895159690349849612093991036287698783781754126311405513867524986337060711184701149105178509757730878466377220520029288275811926329805882081503186391988118800468193567514089813193850786272798489440895496191777539611847450749635306530436637423349707095472308918474352851937099686453429178002386584395588642226376286454615916709556875134223360073450217767600608681789570686949609064438590744903405276338908855661987914516137219256161494725140432411198426724421650982638937129413159838613731515490515170917182537399787842729685963857918723106071905287437344660467514046565524093620524028010135899870570272205135215542708629407412361329972032307;
G[179]<=2560'd115546722739980474480329526131692994171050579650228068003792669953512859360647854133443976516690688130449049772577394838368026047297002651020550523057800187393930491412602776748657941817857983804892100159188344744045978246469984719141374956385660386606574871078526010561538361395085631710410782256718435215414937164118810778850019367723207026726550543640084678360800567617815314899835064681853501816692553682863595739875583700655643859811255763384261892896560075864915397285192031917554354988619272538973997512064548247797180876237108714588656763452420943987426940567404714882233977524899766509586397827446407919308668663765788622302267533639285925808988886909494424932590802371297834826782551066277879148802796646250023762094250363481992674920867917983074652297532482354;
G[180]<=2560'd88465459597797550774002293444839149696732267880398671379200405461091050511869719583291883958031562922549145292503827862461323345206183830083815318396943102397702722640022010953254491366123021078797060194108539484307143163208235353737582529195267971589855778321776452679168572104579944598917672687453018641021442514176469218302168366747419144274056282333920846391359171726823330709148686751044884875192477418204378514129645495853571715985505352375835074584795361990411665334593406209108133830166081460585111451373616330134789414571715869738377131074551948655914113940648994458669896870322766789700875758965029056980125921482169190665100085235588480059775600904026458900921071861498016822022809738303631632262561819213933556765253293404493506698121099330269350327443731251;
G[181]<=2560'd88465459496911983920334036944746879146611670995229149159429173901286300536847225658974396393109649579354769510057292508520030542768807361216477345977366117370483408115341720226433018165226065769348279496058782867405180250475172939692560074894626897094105440616467095725308060253347937064529105776339549297382714155953829828344874569951955346970489177058582192816132546987770776166346213449032478418768724338583277223116602397226147210514608375662940774543576724146177934525141754335238054068901107386090671980106599955738098401837835709611470241469822940233118922141666167620403208360466267412127637629839387339334542212043203284510449689344183043337698104699828695002028285012303590502738537447336427357132610264373500413241924749152427738269965311945704991366629765939;
G[182]<=2560'd88465459597797550774002293444839149696732267880398671379200405461107122508902340104564912451291749485311799240600923575268931774954478599897199888741823811871830568391140822359710144227806943045336776975414239278638245785139502132017680502523599644118046343488715740157686356337020066763924313144456195238732174541698023353147208210300747500325810666376246135323881583591958851738001063095470800768424171316970699362619825063347115528112846761787337314617938526043666361066694163971797962936807986146875747500440186363429576413224289180212991005658769404761603790397673243359909293983826248833946082303161567955160263768448232087771497794790387355343839064787505494268473402721229024665502361127838918096879267272270382854710664228390124786315686044327212785799777169954;
G[183]<=2560'd86766269014901796062988102815302622931738129319293792376741570527223260854957432704307774942480961776248773698756105412408930811630633088113496035940405718162449796195660525960889161098834479158784892310556495722483684860226598778089843227530742633707031600490753028831544886419477253286309077946109184686551400529785089924165759759908697062750276205614589035508918752575834406010219124366409801785792827876402941633315130426116265071557691683648648109672298338601424648321407637773979665509807803426552532307386159752455732021317350079608101515000090956183532963083654678350760744700368914607698025325886916722271118398173354931462209870784245438532692225037664255641934585229309925181540710176879871425622959543693991655067043006878755321663981165637410566661851001651;
G[184]<=2560'd86772880651411118042356841401889421067330502551072460638105906568899001148166278729042257118068485318320449105993017040506955884327223349481780464346649753599749068531889088174423954538040950838867635524942663342595297650766485566229293909044842178200992648650096723927527445807262767606063344459522704332529052643813990025257640292870347066467071138129434824754534942580181786377870319176557351932436050788346823460299262852928595685581878225133816999684768890258005541285730653390559336380548228134688803074049146933067808492525239666093486561908129424555992734198722191106546764305746728729754849798901198938925026331440132938048007018583883564220540049339091386325834982781676951363001044618315796941102056181792106607031809539565497847468658237178581850240266220339;
G[185]<=2560'd115546722739980474480329526132034807767160513149934207133187637855753614292305601502666089666414132916136866416189279274022929393148464687509833318100827192192365813389044246900089360043787883963580114538231644845762338971875789638396636867339156887053078916593575895935802960009113003627298763576214826817597727872145686181607568771114341289575975780884669640822817581753059350783394193305136261399195294960225490742276204801568286114052826555482710673751236233938231484170472963608098822150825247812273548528761143683170410674011732666452243824768634601124714055404888061800860825234472423533855066723074454354808728333517589450549075577633787636706246444665461316782150403040655576190256419666024063074353475569078830607032658508820572245188258834686435021962326782771;
G[186]<=2560'd115546722840866041333997782632127078317276135992351360474396274200383729588400457315570602681704540971193679761565243027243273784211233103331039031891978519302543700083237420485492057635519154044632836153920236473442224093250425424094100376689456854364513219429052182104720216811886017317699531879666435167452559253650385596939909179194370280312117150810214852604662033316581975115812200441863740579723478149223641882708552666527887518888254538193194887938367708850103328159234411372508001845909707316637207610282782612746211340970472366455915002805249690989283364699645513176546602251336873180249789876231645886858867705636187095476622015233314878503607994470412550856732292934063376227046354079399991062457262877620476163141253364093792432384198804486666902737876366131;
G[187]<=2560'd115546722840866041333997782632127078317276135992351360474396274200383729588400457315570599278326571734755465870332131438942111932682976999580848846725591933742976567668843760121806945725791677139426208527215977492027762114716137966885302961804897975190370280601953833566334971409625187346301402358647392808407328396786754363979403043192162916029990357179804188551025286321611187625779893060708640375374046891873118132823479395135733729873417834243035102770587619050954723383647237963276446799209816723281926007984185524782056963201882477647804184301532924033801274078896432525003617886347558199372162215875322814711917943034624400313848348888960246944659059242490196886988381270510515377193607270098041541741916127985189321039906316704864613261477306416649809406270321459;
G[188]<=2560'd142627985882189567843586321954178700299176010856881572124877031960185325511096849405328942890238859072233089536682144250107340336573228308023644419802292336032324922187910040122774765517593495830634826710567521215126068092581455617748364897011072331464523437034947847191134018859203079869610957298989601277399822976045915816532582923374232888565646532837011063447985590587132457702792969334458889791980303486237149143952599720280029958726792860302806193399314961529883822824153388011255740850046568352503892107915430563572548592822156491454374990856821407353116567844935812609666553959815865856121471110548434652235377998882485515416705498428152921843779602329592592080264407347526460974464535217517782707211767797009054971417630554294248553014802228226687197528292799283;
G[189]<=2560'd115553775044671982963061113299530222941617574771310099128747948182707420331616372522817451912088240514547353524591591980517050536660083790938723388227941513387572525268920202607112963039647318406873898300994415080987240245338926413792941142159159547136954839060701714014090574346722732661481120738463730140570658305523945838064186622966017488059967828363939191366554654509702990494404456782381560699531616682253123738478770918704244921948397725655373997581726675046255390585951636675462691341570231211784907366477995295937373141018851935990011119307347173990805159956797443188634847637248509169779168432779018207146140744466531661264910462614037832573596298762940185240248244107593642166824714046143642600873530271064178417163545321226759553914979946649014168379454599987;
G[190]<=2560'd142635038287740473524525061522409471612043050702934850963051922554183032967348669678980549907746197070834691837840203511111896624466247531147307144841913840709772688190797406417301255240300976425453297816460532960947061456840574338686819636060723996524694500782389769499107053427729478517086752614232106047033686357156041740812871538069217817188619877735515237234374988382065427207396202730808830611450270113456341200914426690636658039556680113580497837584748870147493409240230962909678388729928683811036960529262999491030209252499991295811122805483499522437241817621824020647010596757843175493118065577356710547367617691088924591930208668022890834705449967486584810512416789947276064255528170303113344322531893139752844349778461167330626477643533557788365282941527601971;
G[191]<=2560'd144432962649234474625377460308921317708496549953101969166517134816247468544710315962633728031541483550503299381942149786083053474237331274265274934588404887233631041964169225706900189513968845768018697084879535565971396367979193599865676351936006867102027986460195727867757415257169250592153110631924457310454833032579482842385534984607890840807059425613024522740228463719014349742289908780874560776102023450533570212346305641445900212590856974654291217386843562682559056544611817244887516355125806475547523865889838591774728337228799982249645978375176104775761203319010472918105780304864703047139055522012987415851484378535411147375698506600064700798818275040602866212130384412199357265907396668037193110351998651377131488680506449002967753500604088663403079721165206323;
G[192]<=2560'd144432962649208407568030223599843305219609471852869789701258734507446022350914349852882883535220260407670185941399337446998209564179171703339301043391637316152766258160131263835161589001990966049868608165449363226146012703459801059019547162287486053262443509582598132340273257219277309958929561643392823949212683114823834385356984711402262772454374654276857762214449917550708131153032418802067326218604124721720623806024620565636198393538863398335486961034481290044192503522521912833321748300068203860119982990245238285049520541090716120356031172397459129245506411887030745355854443632558276940091024049328188342955298949938661588593871319123487535886082388643798636316231017141295466653593619819038405861542255333082341250611808808771634079263337319235740292482075931171;
G[193]<=2560'd144432962649628661495444634313124354774782849269215509234031332805946638802264592922408005005779631020208022236421400265342719690216768677606150904421430323238249091635025809658182517728575351811081618215943806290817656487483551049264077442896103077859408577514261709112791162063896578512433189040831708984401622496935128899829720516483168470275902949581448980389472289011092018231066849019525325686820639833333864395335404898638738822354798288969394839227711510570104521542473390800853387145584274428890566848238630984293013917851093854194812507476478281518148638420905632514503424871527638465807291481026503844615503124647965711870688562732045100936836727739061533661717350061394794819004881987712606890325205492980336356831983815523111038084593771440350735157389636131;
G[194]<=2560'd144432964364683298007804972413597119466146602139035604920591219613605372430694373675366810812520829812094869611288494624258787002515987624034747515079490117126223178115717853076380159704041923617339601408995232170979954932718866719363385949968403195072418785993697407422894367841991537900318575327449710384480807815388119192854688836845847881218907065538936161696520679201220520670958176736471152430568764549621216502482624435644060633617882015075396152633561705873341794910418825730094211515478999728034543581016341937730249054303934028089828572776306576077839112841327189065436227473881483973740347552493753982483820545923271967837805283699641745869762074916493178354929868571510077383847871630849800610978882198747714410542830608247336876283411340580686299109193364003;
G[195]<=2560'd144432964263403550696640592258539055204017168665215443926926485816475408688593199978852126381060545426929314564416123044423414454338071945975017491865882830351561214664073581250526366776940096625277291499624955474638974063320982625621184121886531264690376252208208022415059008082816486294676078055252237120874608693826327910410407333846502559074142509481271000162218820238855987850256284761082429836588894960668893169543078561484527435373231524125587822514351473765549561391885283193386908317763865908783501501721478629785782883665302280716241418917739702217731447642568765945378075547030100845260885462319398084935466643954157811919910891964068930803205342770336041033811836983816510998737055807832305189918106453710369955427130318578876924772763213729380372988829053491;
G[196]<=2560'd144432964270103079082491362763389805055644408395864439312047140339444566582139733912534493870877803184672234623227304565834891849749299202750321584271975915183389955904387943000623900828148145868343884224306151577078601127801816762092622921351102245196902846246575572997167561208691995996840792545430146231269208710570992063664233807383141815625354574720169335527040885861677358559573285911225947348032191556690570965020364334417350291351609847137800738382681564137104827163262260305157157727930790426855381120031825942827882670738864615985431534157678418005090106316682646886933525342784940622654677601144742192172105611283973747210083072617675905353458487696205698648702793702940013199712157030618006456950136769296519246193704990718296112421977449537083762258824344099;
G[197]<=2560'd144432964270103079082491362763389805403355179173207637160674238787085223731020878878914324099920060225306700766273212009999202801138194772231276595914226826454697539967571848898171785791729942634454730126819312894889910050223848219927231833633029929796146836673442369972845699247547793938129583284928810985257612131408808532689470530915814694555154149087024823284312901262819424481815587178721950692880380889008114868263946502924672269911761499371752314999878548656695990733673530953935419670469979746208962974155139405043738389965077859338993716821579590870953098950896953532323638623413657185864426958803241366279882650944339552240355271497982665278716361063611648697505804451032515217917431414844015247900897066711753898620338441019894387659283473514299689141997351459;
G[198]<=2560'd144433403424975593101977833868269629983028359553247146887144108186321917675183230277447311366100512616356737011469953456808170085214896096673224337833621271698869899461174035280606759573145294129517215324550726087187904439034554152333697585092906040142063108991926719911850611357873388569374990354546526542079288173840938754439515902995059771792705948543666084190184872656626545011806198061888587254826465741910931505167564508386511506070025829797230167519837443954952937409744422225889406885142626786032137251008950019854329302818034069714717912379651575851821453049247598043514797616165480602847774972998258539490219608207043635160521967974895607192166148236655013701839962512091399957387246260248667464376521153119966185071335160027163657744447539157670371411348370210;
G[199]<=2560'd144433405039144662784159189335671034015088476217713133368761947408388184150454168636927079218965007176632751981845655124040491923101669138001717370436385217690451492757447195739329773993332788690179924038630565915242332152801923252945576586431523506787989565973309530549652725484473126293661336561000997484691414681111935363022319920407469648592806008743631369506828629891757598557181612558269974248456926545204742129409111925371991424618788848238772117767835490583640185165542465542166532452285091145736531181117845436721785754811500477862017232468435687476198849737030789468859528288460448955538031117813267425504374863599782365624393602530777447456900142149867669280374094393255204562390693209382706127194338089294789871723218271907739313170678569210367422453570024226;
G[200]<=2560'd144433430973434776750100551007864271741391955345058377099736429711189101240308987318441284501530128138165317594515671746563749717970900693523008309304400179680015742873477607408711491993190754462412096865985828718870788776272447135911444710423332677089887166803263135887102922468522548475487107355628581454260558779081127613907528281944833492797014074502705464805106542561100021958368689239559037248822583145522171652596229316982241610440574259192224756509782656895193878552524795590013954522637163474836668439743317847882649848509501949751044205525592819646686136175188302781966864383361597334589369760940056447360885990553800111079445869933028043511700971437148098388867873582411782564583275409077698057996954764697239227499816963010443061694265232103979806977594438450;
G[201]<=2560'd144546242021401355282619094036979267890098643054302107817891399230049457496491041898318257821533346632320834780737946864112276557630202387332857999030122865375691399154107839070888189981043962166461608095674462648584318680409168984822544028317184389441640887131280966536095983671627947548127459796452329497600796208939399768161575360953725035521923089322641138169690827669906244849678707952423901474055650201392535789451043221178118388759924997247637646703612103696141635854796139069981749922799320406085940835612643430280170209625156280285761362155528532946623475974314445877371301830150896890718503914588284307165691598074789837541542083218512106561627811233594341894184625783249618202659019361890420708087729668563168525807332144465849894383573273279679993101063234355;
G[202]<=2560'd173320084109996983626232996962593971088694688969614854039871639958353695541733800769877442266251813059108430002327149761423542021619093080507489059446200598382524872487870151356861700093126007770801449586875942784372063532972161756302155723528293388695811468885259456010950119757662088863641581716626351572297747679187985876163139254716705516889880145181144445439455825578864155623047945827329283607676129034676919638103947903937638566998932083894811106361238773281851452146885025165826683889199045297164716165332196839053084696338644606805367809835933496532400384018734326872055871573770761999959264933629465000815987592614383706121911621726511640566810854426692128816860157351766999222721911301225549541488868322447933467741488519695969037005743673452937193257329435187;
G[203]<=2560'd173320084116696416177405506298035575469406405440692603559434358843489523483537070494037421639040216194996198592573410104803849074728940439600282713142339987430416543963278355227907520687927193672460845473719919299652357235476533938008039191999156690397890237443864501698746001477058381962973337665958038684321096725606894848307104265768606829600213519428623602053020619019167965330692745094755981662127218632946139769214403785525629416646117670967498872949057148939091939180032867605909197304325306541339844108660989478792124034345537068998241140130598299240296626455983512415754919511796168591423629082164991603778681467970058263933383208896136088356126025077674422591880751283670511783956835701575649151337807437343126083943378728734884804259588757401554809346168402738;
G[204]<=2560'd173320084116696416177405506298058274028523080712472320860405957010862960683248801888344445420172641491905769557375188681495344590999793104431559299363203503781273112398197467212675279585881804109008690072721416683926997974502348654708352291267104169782409116258865233125331097245367444658601431127002386479471036460049193973381494246676656050022414031913637635023298926978834102083210334930420152146389606278828930083333421293981153150723576319345655845942013122423536574448162304699550631840008045161928680002330297424541638628802846203913293045012190326331419347674289594581486906047025424146767691245406139243332589052656042016853282169490360900423127388911204460721478342119796337269428898992103884262374053244124551829538186708035934654203254533186708700690182779698;
G[205]<=2560'd202093926205265772615378191028203749720578488513256486658669992676615569982820616559272328723622733438024479690556296062743752020717895372786729876262201011305066618120568358563286159433915019459743910103955404506786235653940123726632058413152237627787797370502796598530485931417084593585234581831050215008667772076645558429209095118083122547518298349132190352405620065602619578025808119327153422530088086139287685978610748971267838288290563243170609396987437234316278318035736012598334822555499490835941578306447045973906233799763128485518325269608988177982419879507102197111578460374911398198706073944614335742957964248579630211018280901086032974879900751527498727688787852116200521865066897353836535919622257949022331489606728355077018998767415231170225696122913104691;
G[206]<=2560'd202206764794965836355293124224501824937577540447413110445698446391508729173465436243961296818536339289243276370351515517530341573929903410909136417662503692925687750980209920751943847379026077858930456183073123049972839782672344589377244560682045138011129586004150545100391803666408637414170212593215893090808820431295763261071249344001587130149642170709157462733212520645580365194735888368058250005585039032393685226246747322098111369245858102927292592951648472082899266932571277198101239515706997322342212238055534794558120321049438788748796322118797882552631113807407874620311788498226663324141743242451731244662741175914735917484464494170692496800078355680367975038411206186554799728486118626745617213489627057417142129290927768621303121641264288067408995952243188274;
G[207]<=2560'd202206764794965830741454159581067268657153938321535133832722831691539636963707802406167276498144084768787214470417530950934313155258707618137462266974304619749649788627885365528909955846028075070100603964667821850935003899994356471397865522298993168343988765210219948025926312269701320698674139113549741987010425473976886659548937773002491509541168255974097387548620981422498326472423072010523854482810381591728565024605058961730044707957888364281695482880061766162331437290720371786880570471866393412360149543401782216408345837835777977721587257513457317829889600171090945300937602712508816140317368205376161584307968684988568567202927878487333157157976676405371099900783996562827556834535137609140595175559247719320749395552326091418689176474153690150346343123160085299;
G[208]<=2560'd202206764794965836731121528498295483810995286654075820427085133798925475948209467869620386522345807035507224608471681006365953747927821083333911613660621576924717427939097054779208598241036933712999755188557402245893555708639223050420202521738893873715061784157891022493717611621786860275529709980111994290651577347807872833800117111965554722800135672512325427143069889204269697771766246622429977232107215759564471039422545009512653163316991522658207799910711372284699753747393262249844762354676220962021113696264083944983409454961956727092103054955358684792472106809805034564628246580851553013552847539271484232713207419319827113520833757836138678224819784175842450637198825036854121684940006591681842477378982370514482849960322071237459309095525666047797501655545754419;
G[209]<=2560'd202206764794965836731121170086231146779124855504652175898103063331829876715060597335271966355115306760799084866192070957646668382116406207703518055511500184377973743935385459688912614974297876212492975725879517345946991730813693846826951375461112538082111232771235496541101013646263629322318364485237483992559149023877114513296003726759263126766166452561996628741574146784941044735025370963197805453292889182743195531084573103749103915104129183843920292636828813738460365753050106821842266044603308607590808955103213881121339939165767815051840916734981867220958857857525666170366593104581635925229232655417216273450258064750184302981453643780560139415666231647911827334826253977477093417924174304477555266872222613980286915149211341422686362660723807829561130944694530867;
G[210]<=2560'd202206764794965830340577053043096491800135556380731119920578647859914712939127630186808687551264149538066717641746154369418958919648065685995645921187661765078832764982993247537250419530323527764591967215091863949432262650575634323489171619533482371801898601397559152935508026140164881972894652390007569217929892510078093528070426648106030461851235481700317476593633385295720666961256745777887502738879821028855441367982291034245867039213842450984684949100214048122216834862831010992324232786688196650398878976901771652719506122244821755951594583055878292891507034812705192452378031060102741746422615926044877397347169301882901817837763840627285883985217822277874221306987779827657970213386056573077992073293419169916641586215394818175845411536080826534935620850799555379;
G[211]<=2560'd202206764801271178268937053754885931823587658333574027175746566597140267835002477551883076465502708248231130496332291426540685497803200231371136870510288687143285185754788676093033686700356701779547107756368304848031775484066789039057705012109321540896265545223865492458705988547798568529266726143405251872218112916160213144496650530465112424629067884741259974628003745064704677712422003711210598944028214782247000676543669763262954841100418290661388532785193483288940275133884218386754299884668346370166754838428842822835750091972587744076154704944248341535265157195654987337652211666370035471241009178722460024180101761010300620930518620370885811986847880928811878969060671736112417246912167100410539250692834140803553123044457867480578133300431471385888493075631911731;
G[212]<=2560'd202206764801271178292420570540277333961459855948630839145369911508569545274271495622802072242910382729748612563251200602556313749799408538574132097795185561552321582691310605329101393925622571643703864775541578752744978660392990358638454232244503206845378264006488619837030110503949063806840752584377261048555469602849680478502126192530263032209891055497688748108346450152156527907239776880496182954332408139065238566301007337154544868811239275311392600396864723555124987224355108252644597133059203403764701059273201099224304710142981995169892386011647654744604192380418271190962346695484612126075820560466506681548448035605130010217797580580724896394523156871349004436207740744097876378739446183698779726859013193431926518527785798394647771064001912408695950637758886707;
G[213]<=2560'd202206764794965830365534001907012695023734562517921581926628643658586443086082075549327923867822139449773826546341551801340289622045329269771943087845384217641732088880233981848579937998946204121700664805998864423732468232867161412280121065717600640575249258416198919099443314226927978174504865541044159902009126053284003209010075712231026030297598027413648261974282990074771672588243553354625025097367352240223534315439204268632218565219470561952512092970725574660669192476474644021896259119019030381603735946894886635449917528248844856906147999565936682312708294861247870054005792372809574814420556742725085202959541265502370590097872633738905352673081344782450688354964463300113551896235976849793310534877467430660126598494128878947924370046557982701926088323210883891;
G[214]<=2560'd202206764794965830364157677178864076640621615175008045508491129682400206748389683972171994716730596332151534660341228055355785530583346802979167896910215394636252878589728820638342418985028972484349846431207494033942980324363608714426147954756755481391526403844483684898601692274708246660122347650411904869071077894116691436818516209344706924112442104195709434155568817760925530573810491858540750793708202950032824378206479476812652220214152737867797671006593110521033633174465022348373154921177321224884663072823135866738329056831402592379095990127726810661523460946944814269320198775867548041018831490682800862037962529881769730076750187383619855652383362288501598180329702195482280423299283980723499408599439414191089884463946822861116877465450266135384273476799116083;
G[215]<=2560'd202206764794965830340674520211074524302039061178409244843918267594069178829731915380527842419118826869046329103416603794619792773499705284387344813796402390398616556244004549108255294750088926469768640149545095329035949023961999781250607963582309666220094235944964086089853872866574185537664733096575391869945781895187369451357872039077124053389207372579984905672772795682201503391521509709275992657716278284859241307623886775279046932289370331418822258067865047406945288448771212626599131693482247072929201958155129154717088662993503641150899910279378554083823698666130257078862234040325757599191443473304508726305978116274465496367596890137972199759381476091194250822853302558817140085230557945802670472525999842184969967122445210314594305049168042951139505852938138419;
G[216]<=2560'd202206764794965830317093536257706513907397295767942445827164743783456118655166687420624624783904546229927417655769507644668036147464284913708153980886719809455614489240889489076794021831693234521350418934641294066058186744294057218917004178791370486584363225752976100190876297245217634533172899995617198227416281290369372572993663307631950964992267455794827802725312435509182072450964589586162332309188995373765111023795220513628482339455586333200467251469322281445508644077822630950316827379039650716127188766222428869203214234680155116618093015046187012488860908745967049345900265988978012278518067672013062438150192229586102161044586155546826230708682974273457986952282390242802053286006857932545113629662445923430925182527687549723489587062296202672521035526921401139;
G[217]<=2560'd202312990033101929550557182203175902649691532299164984245836705556977977297548108546923042139824876231092072435117313542242914430154799967823713624336211129961829101556502955491349082394121919083945152085857002082535747292498552677513249240037002672602184895819052458295054774708959617626047694329873950019668850765399466638489145930234462892470158949382415774422431987884691895404245923347686160965774608504074327831580399435673635962779499376867828901949766023689234137889112889398064140012463094567066870990342468447488145704259053743387853746472131674043994504054928855316525359455539523376934560168166567021257070571930283018840678211096189307437502003178521784407389352137846303465200019911192010489039721850624477255383385202363319416769206153211869622316641170227;
G[218]<=2560'd204012182337357668749361991948494569039066604514340880168345875656984278955634877261575288649989561799197200820151296229695321801124553619774396007166494240966246889880242024493276090709790910336632473419224892296927321678528059601823777948997887423831286838686005595143553597124990904491558055728808373071776411485167582949813787949860198389880437185466547064940291060351945567193000535977943828728398236652404325757056278089354772413197242231118708978537989748664817118719771415530728541582196620763855052506982148795241977644889481609461531065960043049571043995800318235658393939243517921106109550825369570886019915675485970026064015826503539581861977541323644027835951476146748891352157662383153206183914269957440783609058367668832583698894474169353316235704259453731;
G[219]<=2560'd231093445479936312306243636679167430106287549127325582929068861819036558278314234707966685888424268242247943669655348455543184264906197556893203746389123718775223424177422172782746245515558558739611676916712892132870327377804847310625763211686182652521327835818694066799969875476514688742072139223565073171804847270207368249229141013811954409667807019357476724763366155651116124474090872837723196255588879855816385781254438786905179539542314338229078511170079796599305248825794987991323836005376649115355726970976205114244494794265797116375538431665431923163036960292194476819079954374194394310420038986364764088333801756491998647989426204470806794222049401629926018728254161257653536800713866241031965189436925116794502818745754158498822620403018671454212778384793215795;
G[220]<=2560'd231093445479960948960756924151011255388141323982689443570989006646355925435891960358549974341868608975610202671620564965768235841089168947316334854598995250295464223297954447972598041652726396783068120855007298353100904935302800895774397398040726178346199636474566274569945654146470572562938802632313552515484993305461088910887764541658304363366013285540528697461788248565184226021561339758096493886134750714400799155374711531719095607616782784424984435877522160451673796825145688204637008537203833971196670947503970279327671213528237743802916923018678055223574975680167212448981222365439568018176467020207677779991974046157192029814424617817270890173310630339895386980065334201402447998224269935096792351076979965001223020466028480329498260175665984495460905842612904755;
G[221]<=2560'd231093445587151870156813175184029428501041557337944740732061488398161467380373290109678832064210544324561612810081239744983762204554049967662548296803499871522136858648922517478683135075426326244536839017008234596739099986305994743078828925120034327924190502290461448723130128810783993663604662118816048346963607139745787285242475946364490261843957777748210749438894400140109993226579906469903491032842762071270293428921200813122647201013650644148252140949792117001673188474220501339100324664406193383453180427080927020875418375855901412016594640849506002716246691250715556798401795388962282806938514549158133092753605244458601462534430880554648117303454104616082960887291987285794670723473725394155037031819741147327423939380219563629609939817686290777812780767991046451;
G[222]<=2560'd231093445587570681280531586918825340306593988528419704784768997263065403931639606862211876270525464747524252044375065721036008482906468345668841325659159801197121618288234368495263958699821413299572623582247219875595204177780212433301631178541098828597665943122247699303666860504708047956276651176616193220223455641702895082922511628921869777698691232967424082283165781013756755076619125099880312235332506230544167302105694846827603058465679160254797637540868934988861470545094548880699701942987044557998830601514775826529747910066171673142869440250289565326770826510246912605298623199515410828010255953231205579435369698382983764813506251639622001104633746264389950265198523712076419906717924877042999280121673210192728091658561819748223432796233900245240661888867709219;
G[223]<=2560'd231100470445082663626908380740093018126628676414713026849080181064951255178562785030694672132727385546201337555271768624804602671351754030328097220938559615510617750612282544536217209807523932635211451102216532226754214623710751125121418612889261203174691495921594145797514465900181619389870515632878919719824515154962893565648723671557117807720659188482625536116214343806680216739846371333927725657435819445583719300390330475755229961811976488902146926537040393203751622232722862059389286944309060280220373686256134595358616587287359422053221647784860879494648945526777561110131804081506983324924706667815391631707685515405783459496813116569211669499878391842847715212444416378997678246162264896335776496030968664694304966481290394553634010851499061586191246498944139556;
G[224]<=2560'd232898863022799410144200635368198198811759139355873013441988371542157580166218363001918169690069248898224786444046028151911616899530489626504543470540346114004085696478995828880844917068186386303887671333794186065504048314204882564572593741303655532119086285213402718998481878351875129472002851552066827816459654578870696236571417778265957112927796626873997574628275414141733730603090651618615420341392212632008187335773539787604102831362756618364052782614281146142347566884240576018536448569450334929737400083926687103595023773874572335879457352589225991792237567117270323014507015174344060541349781332314432379326138281437893197613469269482036769011334564504595639227779642802790268391499174313102015072613299546369904036370067208560533777567833839032256479112071361029;
G[225]<=2560'd259980126165376424109298386359235090914110092126904546495232452310328828763000854042727113322735931726442456185064550299068115002952669314275659912264306301772982272192135378324321120595191480046108868247526283095295593464446828329742485868887292778606833507645837857994990448730806628353277473887827599353857188294893623345995697186780862481737166317853747031738038974988701377587297220589328661899761174693554632779197180579805127374382362888356302465740154658021544686066380855884699922071794609363629232078587606646677694615568822522580914241578668628271072715924421379051023615809392378646614619431967819417787074807984820610174005246576074087841929131375369883279543779007822563266996280009949070154819946467159174618260008198320547710046371661920076328493640725268;
G[226]<=2560'd259980126272567338891418779278284760543027027996828807674973010333374187163879525568396516595226676647704190560142489623998578199528026331028235476828641380597114914264184076973345334906480679058387641057933030896364778134617322600267830786144062024101995864399201869579526442666600154378604162558323507835416385470113091791743842035291528178488803605121355599631220499782316502003358696203920768452720378339247197298623058570589216542171664648455293825995049547421290091891141550133345342449460306116944782944869174781322539019026450771474132605662634716653967660445713249641872909048790466263041243209682342256771749147968548192735246085710701166687917846612813498154726290780940240925320382968827046004063448426436952681424220598930973909459581121150382623446578438929;
G[227]<=2560'd287068414278541417250739956073008756696603323301776897854239173860162483966506780529741496396725935175248086354582421636445691994274515244852102062247480798677282212347607045500009409807372043007595194944495523741005033086531654766302694352896105351086212854166989475532257433148094590528421767828246216075474049262351996872323487423925120006753512089419502076888503107602648316943696147037397379717025729491417796828661772475962261415652771291885473869307392024017469106212002314681580660153159777720333006450763646858723653912336475237231727473532276624359203701196101088477227235068268606147877590409841894453946765815196802112067062788525597489935165492108698054796265203689608112161308697452406601227316990394375523911533976717118155297723169277733577743870926791184;
G[228]<=2560'd288866779301887728839407925443027419602680769892616641828102147264940615674487859030733037116766030422861340679746734664660735246158634162216309172284829376816816711665495520131057736657770522874109240284231168142323981352570123154253953316829862552291142975296716021837478502023001028744129446473426622946071893271594955798033964231784625080524082751667346938841925202572539182841357078692178665119358648319006988386539898167329504988656700387599550626056663611141213508533340971465645478126497785796508128337374252538553741663700518257189042764132763202072596133282015009005195163161256436752442596352169455680670976074628494722932981495146681326795465118527329676726388737459726094909160011958304311154276721934672037448972649433581714641378518507532095132949719294226;
G[229]<=2560'd261785543707769904112868983312277388623199806460468379398195466373791928730507219555183690741861799480237111989897204732361930675297402796136048727046975484478083535069853642170020438798377362695279349352465824374873793691303305736692198473333815374219755391546721593121633104430612027811093845778428064601861159362561512336567933791722057810707400705660437247754877121286860244779424497071373466826722710936831792998320163097568422853330556911215690747633511171926220259455141331681833458955555235304781538166792974398007403345311881474110715584270451296864180121764729558959807550499721294143375777608140927326279604546045490525624939546907518229440989769586097131599474952084433512524354405164307671584129347899809629651586284079465337399519745318607246962020521877778;
G[230]<=2560'd288866806849952828218513490920199325627659169463397388304697593003547991654622017398271568178489230080674809896702041936875788655801176503332919685854289612040004564201204532647457894985939097238696769006242976468575397695540054692935910927830217167648478480412800244334918469043937020004977175817106785335510373064653912570094649598574810038897329547464667705098729068568278620799077708822320827148362347785460275432718762359437740089653111767257537260842189176280198833084598506016643730735270492409268423681386903619473437826077683590753727243333465234954715672536385147343169932671963537885027714111214173766142152015788414960547083881976490137454568095518419627671632022273901553074176502915493005601367919693649016676409750503757221085938208916192762117886094549249;
G[231]<=2560'd290671811064569811978802878580452739573683385617813840918293828149068450377716379058269778311603485653577759387136411074311458800636025620211290958269076359200673873554976518587300901784513022913105016733483239565792419829418697337761713058886193500080637318831752464279926825062681804270823353773967881965575601290597291434562589828287238233142849387386348769304622899358931733406676396498202582002715459632279650835545584183724727425590368946188145571082426071037106723423517365001175792596666244812003558843827689086863785952024299444103334232176082569258811560216827609935479689756380881940804336801979635678837631050686959637858214488111289158639199012553543345994312317262772111371448320729854701944706275070561232886335093154062372179828344640604126427641379238673;
G[232]<=2560'd317753487528640956892551930831839954451587845253445056667297585754098738066703503374875883920130545559481078210584224401090736215989564219510964992073151201782205439089171330265542671686200279581500684783185814037053884484232578840096622186902796321408160624711208359760704651744937294092801459325352192546817444159676156882486357602807147607929163065595786725331329583928363839276574659838644685447299253389027467999933958049087726232038893072781756242283395789982126234659706312961489265536713768073901264816647328017447258342855513427118332100462104997484490017455429932792081763681812681704784539261398331426228645024869424528708362576531672746663443898700909178689698159556308371322387414505319796249378682863855686003737100880665569945753718144611856423952877637888;
G[233]<=2560'd317753487534946304820906196863095721361049656360688043871920598362018641614664162435430931830708568903991399828856693504965212544959383466165884895718453741421385346848173037885631722227599523659654551283810906167362144311508303619376306928948042475204488427239316777775775689843045496394615045795895881578711061400350525640947545302674484824494903291409950875540102316835509947024195755539246535576482675098516069508796038169119767019242440717328063743246318139191101510661876614901740743249320245868951820415520724603923415817212061325618956667696410530667415994850953001290518166060807543351511548426091572333246607163635310654371037108590041650222648832141901768257034933659696122693782035511041816840081431615748348037276869635349793821785413117403006605218923242497;
G[234]<=2560'd317753487534946304820906196863095721361049635716468789376158561418005251405462122663003173329234168634697303392638864890950382230740818640471442232066160458278742919226562859399298578334854099586072417858392104424115943901720240430965803992644703472996350633660937248386680070971644410986843000501442935564996300018319248043650681760421410419478717118433965551488143052474817262472153123881425871371511592416624030338830872422341560160853828155598233093237157815526229563088699940505526578620180320975921089325746682654905149818799857034365052332518219837466833676367603012304589853433019582771589578517912943716508784421894731527331778700406581776860738794881459247415367750368791270347146628488077764014452641173673163170808463287181381992055302421902468760256890550033;
G[235]<=2560'd346633115807664813304606722345925466120590955268164107553135241711410229105460343803143863816138695029930291239723535312302637638495044124732087536449118208536013580401091515188395631836469810850316147553075511721949319069553148550930643220329889967915600569231355664125450328722640315222661840679202924966417446113708606003191529569380907172886678585163212756314613040754864659346367499471473781623487158441167699411603218199376200332153987908614864170589957569611444240833587342549573344201469774545701136323338652570007492007079964881131238295181495944352300053518391526813262381466982932128071434020902977938697782316838151604982382278514466537632486895667201196481714321758120043181921612075545064523786754381365567572390308212203165121902376724600194714790384436304;
G[236]<=2560'd346640140671455967932643336770908411751187455794182028448973678353964023482797298370503485188731832292530465482229455254042050304078386972400869902770679299304822856912225679469522007468432740245698911053047827792055929109042935896014374902501522941471188820091421784304078786110325991206731222806939827524035279413113234632062930178537000800687180173013493993833991600541474094473669868649327846442535330327197126435959490905882159444189258946992308358041782436004994283321926643953323038817571956272184092806582401358485654633411959338726714447911574478389293414254649010451981437918509003840049703488634478698345306008787836598584268297268437438912512796113573605622967854412163673284007095547969272950786742212119059379165224287087202153895426225928443631880814854497;
G[237]<=2560'd319558903362283609294794437299319722185762739584393743815402900440811549555984188195606313626891260603197814920607576003121394303489926926962783142601883099049968794547520523556589463873129352473308065197357183661891312941126061183569771748396866212073929938394845888228381037040799873415290007451441673743220439490939734200913261902450795664551771329182197114989765833765773866155392427527377204593904127926578223090794259755792235158505541679684322663830759015795246513299056878924092980768496219532393913804960821204465577847011700559377721367440163092061523412366807876259234482453695643517886660274164727285562000422856057795822659649293467685165428597921811518129055526503923476355216420226300136264174800701747147429650723353797083882204476386219805577171934781747;
G[238]<=2560'd346640166504466532625293646531712841363468429855998473439919041122008268829779686344654337932926933860967742315936960715237455638003939934529922246944492410806883130005709900079757883578524843668608756517358187192232884265330685006823621520070297236380471601758142433337248160053254856086320680634335139985876311478025031408066592218572982812168465085146864608356385055426811620824642919508471755708588883144512069090454010825852764214234627144742915783705528474575094836439751897622458161123903891661410175657853831582375333952348746504962942179155671428914631210780067538504057209630560124191573661382391225988596659693947511592739096885760250811705310396729305064745074139800326145673627109780677917452549070340025726283455815234707746346686413927571647888032807338770;
G[239]<=2560'd346640168213215815196051365719374220388627347852853552644359060687753556732950158243961029396029608829676582315342786364253307311707995726316143220238164217552882504871426653216210923417635116356216300259341226728323752756515988020089908800583133769882002305705815997246694736807259005644810293993424463453859828896719258813330761138356729876818098255189609228681769148983275076458367926216562045993545284621589448625689425081855703221619913337804236379282069908603432800253190854613661346818945047937842541544458627744053041432573770441499807761924949877342047630626787793567076334380145985654331836233056100879607006855615221718393761621845456628564393499196513478880495009748541504655838946882565489486924149329614945224338474496628306143771502965928328517036149928721;
G[240]<=2560'd317753487635831871674568336370618740935843270893601456383635861227088704390905521266074136399920657789827050027267611980113682219062085884403207437633305100965553486795158684853434026131348595657616714499034679577976465411444027125149006549715592259011800939685759052439683104235929200919697373268882929867739559032382467260336401247544118387475480309035208334159245626582927515076914991292297606031910074626317934512679501990421958683353577979882954088804125217824967394862674942637028472427928509381330807794951043156962858107813777028661905180690624102673977987041176538660614034242406687641303702257310393491746007163905012451919800309284803944197020300786557276218896593175454115824497690487473291623586489389529042371087981901780885628316406642722260224350527509571;
G[241]<=2560'd317753487534946304820808324982329514156719573147504920358151399068033120374315371344616802611882374624057630365710201326569676981855341487030060444446368820952729887121023057154605969925440708487967600213777011719972211779674900974406968458088236443603290395860466677315575003980894797575967120367626874995178456679678582066729142919037304322478962263685159002608596660491313120648424633685077528786002072308887333586007561764314226284503269231458760815522904016547905579754044129311748136322510782965768506460331498522311758402524966210302639771004601137349752734776941326371252117457334057419691324732158522537777106590812122867528578967056912407347805582223372741400785851007975396336618158211327644211894253016781540827960406906645773006907962746808898721823293847330;
G[242]<=2560'd317753487534946304819340246858682500312394912349154612989669455014900130552183720147209677894964172409185024239633126959293371577583395683214086183350512092329604459074647783203211770521242585171574889328885871164292626241925024620533549671996179292665234208426706839133174172998318797910747184693072469850736651869997054445390726508268397316137941623846911495261140094586437988762029128469892875709851984524117477187656262586681848340544379477891131462512017365746844702959026423329827764783689904050434557751054103978105059228956263095114171571322795845814349200824992623802624597572461361474421467547679452189602883858390198737668233317105687185316069831432787729993103655122376390084980610758360663758215835440767199556212152700981328572734424545837325266493014939171;
G[243]<=2560'd317753487534946298406774596573632681860880662713374825203871784740808342479256224383490876789001923965346662407464719498248229013804563883909327895663744073257202605620701626824782375838976887714090437738990040463297860401062140287858180330514917339878719351740893578270489642361690149987658329621651518720270408725944142793491895731738806423796266323596575941846561487522741451999170403814957863916161747592046999180566876414934514415818620314173279381941227213610461660284818447587105481428398949743542031286516793505038738201009897844636228089061712917131839003545317132736583541304168076122494589553670217382858973755309823000948057969820511085062914810482104112060642698665030366955860312121342188395450239794470151583327323010381989147315266794368365131797833581905;
G[244]<=2560'd317753487534946304420022971850474722804381029319755778379669490570899920204618992923194716556560125348442963386345487905419111440006325431566984490355763010355828206362327959850109414899273829977298106591487092451160817622433250656339838101308683190576874259950075995844105683633960763663058256281382573025468675237397429988759605315216308867362649529339566646723874444055012988363183046817326810117471566008255038430437334787244096836214645094845641778920094427274469572287693220829736414222469787905024025674894170464259992830932575228435470799811620966493239133460326513290265114911647551278813457323937485605847573796587975284165357031052007122396806693274698920673498862235505670861500106301807970386792186519831052426552449363148716418007097536901220543001638601267;
G[245]<=2560'd317753487534946304820905814556893761859029617855288594279009145886009901709369308622628529462095656516759098274008764731582372613946352489178844898998773619428015270152144715196667720666256535014413719079539025326207730937683786939847319454547079187607084715250428534565854404511291146873707247942042411650475008548721035830765976685773972114412386612513374727295640300572357446689371975902132517731933426318449656646968425137504644184808968622031419965731894491726124740795375172344433677109435131233504183363752645475637169861777767182747283646549936418238570693907573762437407070721955224774274705412386659578622700917643571198583053485548799656287692538970287894954889837294957684475354606263225829602731872275339409344202535018003744408593008102352424386800378974561;
G[246]<=2560'd317753487534946304820906196863095721359691411162319281936343002134538281017069286086342040967392207211700730031845177039557111461114168356536906915049938231816080135130069086283948192754105438291879143991277899250956528912552926324211430809456420973956867888566584731121004049392995217562298725149446923729841711868498257763605617290080207575916685124727218301456631097865278373387964491271058480159273154941775553785240285333153808535068389146033259631458416781692674883569980638881811122907868913954090800650342120673251790044990011730968404677631146816618757362457649337447345795983223179291498196717796020625773739862873484213920786270523110931303127351069980998168493455851256804520770282666950222772363552742415032693815188888216317983034165528191007038329080533076;
G[247]<=2560'd317753487534946304820906196863095721359691411162319281936343002134538281032333122924762352780547774958672088107546660768234896559746418952852087544378346167516470065611605808685856453589435297294020594679745492849145929085397105062626607936576671475958146060330281563931301352734366453411164959458706219937018553119786433076165469678526112282032115204978782108316890119066578133779039461800887310167527660252551105765215716888166981071965120291626602758516319669537714367142678094004379342477666789700309944572991717133095038019578035001304789599805403827336154542839827580332645252492260864204015747463931770414377410044377558021388400772424071091478366449495472657642097515971501027596469258930766357080708905364985561036198872810527666566119540785050931845798052389668;
G[248]<=2560'd290672196945163595086007583775178341424637251958871203582947346900691342953243384311177692285142473398171733322643100575328497666762766255183903879118342061946299668795787163687125551007788684826563863369366070071324473859490665706484297738655764833093756949352275275726712448624901628979196296744287680295962213197109081716340858398528596187689332504857631913641991633858133551144985034472607992091806248964257010440341555302444171257929477481295093318861142121548583292124690051819819164267600126417771212537545594154930807242507862523878457874005786583216317230650362905764155177399280325065992596229417984613256728800406283809123753750282618620776683035328662971130567362960183620897698137773847726582552576162889344978729510734110280315525568999700564724053157679908;
G[249]<=2560'd288873418594045513645358069830705190882746072404512820394964922756526058960857841996408744325414741996326290199134598982118605957512167641427078468841999628684952506083971873341382095992543175595001539342423603106402141769262175660269942353177575280520062709690290810530931824217454456570778543629861913476682888220206542129956960442068682737189969812661256304895801367697538288330567505627552600781444209352008402455005221469514970718731539764859854115946374958893682688642242964483707932035383832955992138219995612086563510000416595560652844995374382159547876445577406189239800839916525156336861463381393398707168158870610860829120018014063036496425796897962306661355082558465660582726076042679665265371328865564807422323609134193343801851889032115069791287450515419697;
G[250]<=2560'd288866806856650618376266149196992828230901344769810195070124475989712440186637500730734432101534195472004997871028518775251265747544649870451286184992485164031548756069403061657256857496299640980041625143497739594619950255640420570703980138861413258274859280392063837250266605199327664431728121142458520929327180991347831036453464567616353443904419732780585960208790698405181394309554669401493814517817643569138155729757278241806561789925158442646903592749769288453806032871843156016653220492817233137670714543281559820063420688355915254609623114181650272240940872584298250532896624004947980742121114385893588382425008061067839189173753335051882386007296613968225044432022769394462975712482017742420480166353550700218601378922666336249757879453599689110888671493908406865;
G[251]<=2560'd288866806849951186200823815335556125969617539165001141147927011766392144313567624522756775424365606770862116583012218658109586039576554475309237278199426280520312948551758542617425841852576098371371639717010947393981796986962709432648464458750285485572003246874463179163896142377572229455732121918696150572694968446348816028811983574478132962550636771202384336176327129958193920657738177044644395355980534719927466341620650316491833618380566944789403610568657869051166447057200031782846930686262238710413159123155711556989467434347676802402382062822652404843512464914085126276321753666207448093739604772598738459604277194896835661821822877036377965017500910325930511748163834008971185146359624570218123809696433985930070331585686333700509471212581045651595822607927087110;
G[252]<=2560'd288866806849952821804381890624925449758779836803716031103896069753290460417702851177718761572095211962549255074068860133937201460473573320256989675438809688292702885342915954668867281977607883058418040012960079041133293052170482530438462899494756124717939871203481390741657001121140849132867871622374949107250071409493313486510784823596785141884976941862953621535351871185429455347669488367046925854843915803552924772241494692032347894778980454883661405939941733447477883783995918479413246607001792351928681200939283567586659519125068430620332128686904532137188340319712287302327390958505402277522126900937457203434911202866319831993620104420494816639814740592468180094483138325045817485211020435420019490088249368626774081049883400211682698209248081304703811250113503506;
G[253]<=2560'd288866806849951186200823815330450196363768418821084198321681891067064587276912289283259899764264629221684649644156498581266918122102141864141382482941227090930313749583511135612640536330685123973604328988799195212336900714891711925259591690416101148548207032931299026272440678038377953277587297870535432039183763299935062680123965615682938567645723623792161587359006901414654951285298187650529703658232532234989431935786976723043961190352443906126644276737206386116134510245500834816916667413572646429876328625185588705312694440689340494928710796943063364606201433446756870849613749569715907432843655390652847876483968281901340512331561967977786479116901220150482594992951823738975707658421227631903800634850871536158445280195316065202428830333184653913546275002382316544;
G[254]<=2560'd288866806849951186200823815330087019417901282875133422202822514074411421053343516317351130774691181089783900146516070602244424300946432575600732137625821836791731664863897178260620349123734330567590029973489452352272491288814301851113077415822597734217702145266784378168987953467793880761040144759319747870031466024841185001035951667191331749134138413444979116736356645505600517753531012645446029333474891183108083838709254879130743761987120557729807086656579377826159342755069305469901082035384435616035294148824583400392843373480760148462843606794784983627066004917871149246363274224513327645220108275123222281724540005808811645296724462343645112943725356209049647558428533934957557452067192303584777455421964638968017256771912803224170324965256013245337523913887843634;
G[255]<=2560'd288866806749065619347155558829994748867785660032418629910706144487718255251768009000171465173196845750318567723503333292919654841072644995301068276718893067406885654845649878003199110268575507863436117174678153023009414765815635840490322140354538253990323428488285903617767596243051368726311597768793390365922945896944282275862251727997584913477190002505346961584462225289987646667457494613490883819952542033969923250399555890751272300176653360103681546221099252643721974300363631936451004418499847037608580126874133927166599500322915465505560688427460869742379280739176631041368552476265595630861129233885179204090453343332018922204689518468896904774672521687949712839813872669384920551696492560168518723472706566523718910864750895448458956664466314041332529513991832339;
G[256]<=2560'd288866806849951186200823815330087019417901282874835710851290227357013897529629086850209676794964736857525990266216064196636826112978513343536275708516407617657660936699680802974935273879540581048092057187235141931616615117137843287508196531514150333315950483162648904018868449776889828092277057153508940594067486003252567631272596957934245916705697929755248001517419410310979836070602710699189524623860284048390972446625442780858580595146812058310163361517193481411490352770422922190705914915686499971545411583048188484504013404076475301795160158129244902014854771954181712163475970650032339114052664999350696255627012868753475922969824934535743135701667897892052393823233809176031582040282030237779697240296355562733070846656035160082924422940052749121503354171671257137;
G[257]<=2560'd288866806849951186200823815330450196363768087218252565323162462943241697267191316678794105802145149376728691626711116529971847148772814672022203819507979812279555678138754820737372401219529374803832591505864725462202072959845370457628697374952150750026498331747707118772727135613790834417212487435140499848649727295518934856955645007897538201099225485301470186777239756934237363155436448075095359818522992572796607091988975175926768582967226411021040975649390894817484626313553809020147251285566279851232288735333098916401566393676993567558312039010496339500838542127768662201392829839009491893323444203914083226239815063655692592938485251388274507334717947473502045031072038691953855491142172364204782713149344586362310369255356493821863221135177867931577168131515416691;
G[258]<=2560'd288753968354410997286513975322589850922108738490692825520404341418666267093450686822448690502813658763268228520147974815307506058679657786996564457563092310507403865604056895270121124370822756444514703974924053990960680997090943306438943174194018195702529412014504704121608922437253399981436031659688793896641345343895919914999800619165184321320426172154394094478307520903407325060025374749198228025131353672198047223901941852815782533748726945974538298259777699874418435650682031299982534691902027586160256951274858181066692660782432029148901455077913833997285866894537506311478946036425282927213520096422016648227514656316642422658301678200118897561905056726039585869353699458855059530976004672702581260682005475022719544634256511709586237023107243344150966702776131841;
G[259]<=2560'd288859754437674576465325184298362679477532022423175708434219335659064361739247938391509687998740630510655911370768457142252681375941873599687851934475871685870353703480936648600779700003862469179351319960607559512028068820741358480943990702798712629238921324225393462122990947718579246022787890074013317194046560997445357938529515072151951209961066069689193936848372291531815871563382861168544572461665049449732252279462458049804180794763473545986552174815854515423837023586907748169539636576110493961840981161925627331388600768242992815911901905872005553670373614040487150730911176555500511704298409921488016362284981666128539591290082481563996117592418909656206916845288167004601322302655038233506386055285563718474381121224185364824569183341226992872126516133028507665;
G[260]<=2560'd288866366074185540084989624917427652937348192253971142444963996651003723191795467772825051880157570085497946996492612617910712103914352859075289931776090975469258625873647002236173851630573344808598352377360094002072462676490070713686829574755566707413675342381883337800456998634815258233605929464435444990912580375849944482720047455563001001209422001214231217954683315622763910400308306614102695112971057762170517607602842439323256627711807760688009065392235848329492786876857048423077042268528185054258225473855986356304154489757092021670584752301500686759815171058312317444270307700995173925599977809816020085594414466663174243294722743821158898250169502047637883954712963969747520061803127952465890353137809263046045669230406555877871828397588943330114499510460743680;
G[261]<=2560'd288866779301467372710168249295366491349205432114369159506536445585034517644044505990597003182326458313939767222387229808677520419843077369903492395545653035547824780692874747835242837048433751628447454702945494360827998830308449564652236277322395561633723276555898813924050351383773596588235046585780449510605614011418390960770771253762821370629772686953737074772593820683007090070476606432602710561487490349671548074754043622202197116576996738853098891178580346514207259494905481939606887508561915010458508662357840369301111587984979647190504067934702301596783739663781545361641707803778584373780393532396866088576300502934674811694353498004122334508193149894015152068089403502085978179353519120177103869764756134316724697491034083380453874087118458352729928863081328897;
G[262]<=2560'd288866805128197117514587047170309173288089411492498722280452012207287841401659968952497575416770108089621119765774618796224837792023120820273290504443750426080893154094256549263357105037492329908487239769582475169404221254549188878952884448313991837377141947215722314666541589937132659827150521868631066749269107226860411034930585098936472246855475348537265237051321542521851195008239884214093512974260724167154896991174739842682904207755448885106001735630987723285585023173838145611078717632234335410516673032620744058761830112299043558947836354826488687299548757204274708733835191768730933460460449884244235781359834685015840799716343749417792326137484571916888069517542850519942971490642584463769670061897324925509206212155732523981557227402477271447986213861111994131;
G[263]<=2560'd288866806849951186200823815330087108410211570320996007621861642151374733975357001624747737359291639488807931782693343896967867928201506212027261417257009735569120094117393727474010032830033799144843078741403104088867405076962815996351445607197797762034070271580601588566498057301992181646997053680153103818410705551572516546616726820978099742121766519765972090801420748468341975759302383861540393010189570247636250246850145358025858368587461536542788076425206023728843685879842052303360575778752888270238207184698534283473986177916185914373923924622589285090289798531157581166102231772495065888046406700661050965689884547649244912042413545636850301734917186091924239881050003556612808256092177913119866526869659344615593419031615624414408878449460479277871098880355222786;
G[264]<=2560'd288972593034100338246551656083135978626422822274251894609128408069459470186683692279474419481195664822074807256602501602981106734659094959729417682119658610637440683738754564798097428747217992296632163317503805317405646010880587302980726873968512134772973930897304068150478422172583659041109837625498296980689192312435189829569162527619503645163484471112412403909398923628735832340194060027328686272765298823595857820526933850015833131447580853398230456627347456322057358937516685738664356525708916222581590094785423467901370177645156837906312566127853713577160294163359985262218608088931319397424690404876034670228983106738650793202750680463551968944449319547173185180857268151436873169967578570498429611866887194356886900834734683329427987350057042134554157048649823540;
G[265]<=2560'd288979206392363728935646414289956602697065626820539360300630215794367649882158704765439077552394616161984979863403359397419825661077741590252579492986945902360865170995459268876597790498091022080130800477697042143341453843391109848590905268587165358646458907180668407061742920161170260216064825319918225897464353061603182698521966821767102694863695279307793500330115247336214203302981656187266533812128583596588249504153144075796508065175618707534767019293101322960415184463453137414146930237731536892079409566035985797739013994292488351779107879274051958129684589421615337981105358299286351137433635245943513074298921744238856322858352327937571729802626797963665922639428629237583813298544267340668760318619286141618171256065448556913010942374479719031572420592174039607;
G[266]<=2560'd288866808571731527170089275939457119987383974558214811889990736112869658831157526617836584578962982542197840324368761559771738025686959391318667213886656993161035933091974972827903842298193004971862927999962608133391728070058482639388293771067728898391206224799602060667527060766200380769841010611187079770979995821309539775798128045154362257581565701330220567086728552341089926233741539036955410559729814625540435352313605278829623435502551194015846998047385139866344742913572763234580365416051886260591578843154024714249465510368648202461015805276408403932853631579183003190400558329541162725521174368970429697790422581413677528455675843923405449078834088628221405011238823373815430344808528228839856379754338452760219612299606734213181769683060444085480775699979055154;
G[267]<=2560'd288866806850371542729380766398837403878526764636698880405354821774460572051629806908208243964932161628903862107136205383966594466234518991217713763829810039049097782813832926779663454846560872622889655498280808743905164390183472121721809222568792733438012370137776047080319561557515207705847647740220327935731579339487687014813030115009946935348991525041279417524007796579793866130564634208841057488378099777998053780059135173317332357236525139080096423775968696020357330241692480697558558317638131954172660013889114464488397576224913878906142475667116336720019361951303563666021593140115140158474425595237983991668381262225155227674230761461546503942273983579541468926055480174805358988038407628127814036912031758339066718844935857753428974353912954388809442842254917668;
G[268]<=2560'd259980127886738050567702686988765374387463685668492741581269237612928300188544289184385084648506636025451550350289017322002953307527880435977313086888477334301904566662313435133386344850893739429575031195126393280935885252793107524791469693001074910667954726859593859337827640431173805275172856388968468163873997000516384164022348452410826961299324157935298407899820876060578647688201404839739811074916872136715986299843765866665382072809559866946450122194001504739942651115042526950391782127627733776201205449299688729933098037427814204440390501512556393877987248107001685317014031297806161318530204445991211635076598920562063746427166857882476181174970510003304744060698983887496647983036201211342664481043920630484489821728572164479001228095067700692986059954400207109;
G[269]<=2560'd231206284076807068072208925154137932499244762979111942031084592826962664482239202021839689082367403421846017800157422778836767745513475128586423627181519529100407948495094947936399429167723501024157897939754719846169382088915521243969155881126885214566387779670744895074149332318370099855829547497494537702356422968896106596595211605879502454881328711686562411243232974389030727439056990886967885760448443549645436742042755582037687890359611350354400477652440683847418900778243702965204253166863218223498614571488829153570209364388381870463212893737595274602171150241606072587081400303585834532550369858755260044204538083152557376212466653856791970864693418594202670523493451191068372906763228485665152397009456529149076990546131722747561284940659583078366900247890313474;
G[270]<=2560'd231206284076388353160458806969080815173270010969867922426591326308640952126204315566114774180626188682001003269345552202769191233411294597675085320149888359175378115136827975609519612126397528066749981550562019199488313522879065744771609349595020739473572099354691980745074368640336570958254560438580544826624359008894451467627990498333220698169075529616087067680820692456618470032535813361115815276247757411328045290197060101387540762584220658740356729212164680563080840734810974874601506426767866903444414699678214439889651667522772158815487568205660381741767397284113544974692481362880997065421010628365015162414097206795869559462558087648608323083364811682312091368286684564321375610843936956973065417706108877289401289831937419339484171633021250335518073081741743168;
G[271]<=2560'd231206284076386717556900373256709030610308385603339582079664494033135822954795041799202521645853956483294035418899958677300529169315666078520309474361505387453133825796889770515316921102273355268614370136431467070731413640964972657709268900787920458378656626867458919093949422658060739786735338348420880937362633227330405518084629399062766114447973274440390926297578043635288920053593940116625549932043684914930982063644827470818409306044374801582693425637551838044345904364059026429808642112399572703395439811234689259079474818695694078043115273941330278243969726421128337341030925304253930743194328097860184781329081025743971749962495718471346745023699849906678613274806921697263836330935616664118145415981202484817220426406297083852719897737706953518665711571351635216;
G[272]<=2560'd259980126164956170206944910402568357759739897830253428175450975477193537511214202205758539072541944510705842936295851007667956349498338884441766373585211773658374276291961896088670179244196207543280331742764411749213944983505639941838562159550318713209567893316103897570889214801604840679383399364426043055682684102759738582844543572177349048574551992802885261760996890371309338105880240132843955507327373078240168954020568152144459528443774839881613856581715494045710659091779248950790437998583934349458295649539794643485606172400731671393377765082252668401627420085294658472382138279710688357143215476838771712572587001684582403573031681807145999688873281490313825064781274753536117915299900290036356731109052330032787011040081454820081255164868660078505676641227313664;
G[273]<=2560'd259979712937674337581668796455555741546955857889300637953138093237687103141966446179436402153787085687687900759214031696076110782838035426117092126857459535059698871752351293647165499840997315596489933186102051577948155651180955562808071513458125679188909936151846897334798803375168817651365990073671971561177604394501991615783373792713511664197172769297514672278541696344882131997530748153966133720270964841078631506959499469774492895508082819900421574127223481423397205554442353955871233109078200217665086308520376671476481572244677009292611009618311972887637082362410927358915433548643792462754571171377837933669145274275101969235652226088620378995013973068134868703895719750881841279262396763658787669602267576026995896544600585236880107954586328705071952934292854049;
G[274]<=2560'd259980126164956073994873416404387771879767764713084839868115769697150106840967097548740624325058552166103961773884170574196666759042441147929355476836889036914885307465010161558289013008780655111844753552035785853738621853938442540851516865884935594753725048687498767619511090898233527840647089531510188623502524400671990664446147259803056570932913373851312468625094533473348926560275922758108745528109435709429667047534470289669479610093287967286971841244444110661777429790903676842075140551310479556393673002415115328261822164071689981754060754332370049349074751036844544623796514329011916871716601847963906082785218117536502705260948888024398213493285340904726015622097572284269846746741488860637493538949941211904735187033122704822894118521101243452115873519079025296;
G[275]<=2560'd259980126164956073994970905973460214819040537670920596115418876115233572016013264975497022760341401074898160582289269214402742995435381832023836434498918134270752813241479018343110618847102578326032908861798383711226997470467402070189841421695902126119601733553253427467539784650364553378619963200046358355364875833553991477187330633663197941580940246974020682600475245729868755589492200411392413799262023645399450312079331346621994753891190495309177756314301294844968722077346784586122763601032561409730997851367820522186653561049751777644329010960439338464333149758130002755632998914446340847614803496201282764026484350654261918434423867464843242461812404478642757107072218419734386667315146304506980348402389524508473834306966146423312826537282199166769833039757513824;
G[276]<=2560'd260092964660496262934238075663502775748204722563419237099712572647322759733495569420634504956713828313269241200588294461971058037293557877960347321812615908442662872864577076845573936388970808324745513004037872467000682419691993218281891067796749101998703985523906639632996421770375629531771064229539569616846315156104988913536250599360697644407078382454878593209952609356500333731542854933953894722723531379295884347934057925288042393354999776460612463025325802406853819973734435649675132961456141571725513549513963338319343586260679586334752024459435937797673172176934170848442098481667348776585404569324117761840824938503000160569737364584128673329367493890070735672650203912727238201833606486467690115823287762054237823465613133196128257666459911649360638045219463952;
G[277]<=2560'd288866806849977458483858624777375723557523307046579907333923193189318291702694349702418715838387540870116326564592233572951875095367895680569159270676212547522438328233677228936714241600006928960369527023511195327399097328390450314955582545191444686278130716162292880892038038887970019951049201530748756447957443742823233397557311391392338412730620520428074921245221695580678292072519529865150139156214423734906708598944285956002378170050282301444088488103219300650270272776247460470634327930047954360149340743967064497800702283916746999418000342347274250361558757705776818443462852701494062279982720190198610585924867756817068941728804104294677439074183400431185028313282784443833107945738681641476875289694369122417309562276796632136037812456326151775486703731416138576;
G[278]<=2560'd317753487534946304820906220757597944997666702310340914600483378251475314198117132096086744285405134186002470671315687952942109293653375299047967771292747631952511622235956735494338414074057479974124482479421944578103737956870170053665845089798971491212525254959532212499701505860621278977856016621834916902578354973162603568293732661559237865066545558278037241149219402416139049820677912163369051688268885090097064009528260345451479238509113959961625689136013404425416940046882273636659211640381953773487413716720830022636615616997487535212760470550775123154261761624887513545079637764836141726309058007700847133251215244580836182188935902750402764174201878356931787317610031170522585806227280085222136320957517731139542476139142262008240720048985358204430457456691497989;
G[279]<=2560'd317753487534946304820912313855664972681365945055857243956279001569936844099366033337668241316817217175665139972853718176074279014575419431578537422048196320706055417926821023614574034706568674974614136631648404596221608175974820207467028267555528140961658698132427384663405766448321310034753654001299093535861317617134597920700269777586402765804742580374480625698008757031604878045469072656718238256598834666804568019829063199566103401546202714953006330527039606291238932241184905536914134507181264219320426675335728562553113468873188708259631676288272932195269755091136241174043684121525167899700591697436303115530918449321085962392848514237981221317823152159711494164909457159118889760685712013620910724509387692659857120327994901953238397596333795647466134595055085312;
G[280]<=2560'd317760539947222914957288052913274678562313918517858218355133984480458333121390479808294016872729976557907709006443464120715387705431074455934692367292110082219542560035226217331809024015956384077966945217453304500626804187229432273137530723620886309524665908614024640995583707374822529769872825486628675651162789281450665901937847722151386647305100592579633632052938662111480545865300285439156431213946982940105240071339966544199331454353257816570767554742353925268269865411157865026609722798411503806446699703701728069690957341476049973513636153288921870590183392463005416064044780826202857962024219700911216179681651247065294687131931078391051075737374745921831795925062836938915056991209736072814104065826496040408726739045825806873734943845190185919687960867428049011;
G[281]<=2560'd346640168219941423440988578396104423301481539449802853021534121948074949350697667340640358627512172922524706403888604697671410056553996887674398893406435558470759534212475969434800666494988356339875640795165506646675661852933549876043897486022064776921757223760732549642273044228712720332803539585904501758242942227382639206070249380717303530263505842716964842420012081617538984756755181043891394945233883686873286216730350359184036226038064648804285405457713336720612472909227432506660328673921646298071948835036632433794836224833587756170165071126054270526236066095269338256471831463950947716172142017924992900213862853148038629780665776331929401485330129688343156941455923676635446719152277845161014505951728248590963957286883190229424892514648686396088597128139911723;
G[282]<=2560'd346640168219941423440988578396104423301481539449802853021465111213903647704711959299071332830110145284250048598603537797485109289721953132522718287983672211473042671024248976863898350479720367322640242297407109029197988359681530744583600477328386255891991410114549736415609453925336769095809245479171259470162560156618193987380835689880864010880806095006626072514386772650257375035620476340993892425927682048645632602627204344846695989160410369418013444044171908315860278023771140003510715840110797369115120156926567547661710960400918175769715620380559834642144919213624399497743570416378709920093632993844635664188715098968096004237927874844544364546822777390816731290747892815904189772368154952831488325254370450544466803207691421748324666729311428351386061423017100291;
G[283]<=2560'd346640168219941423440988578396104423301481539449802853021465111213903647704711959299071332830110145284250048598603537797485109289721953132522718287983672211473042671024248976863898350479720367322640242320901313943997992422655923442495717101394746904960090762313768277226082751875568884825620916857419778142904351332144255965788973845704792009944449650600585740075454214490789079052852927751649388053851954882129113600537121492449426948123271526107517119031977250112002911040867988387955967284660042771022310264683558193037534237404426185709226116124780655608367726673271417583573887121405627068956550485834352145776917008927007952655436481757053458158182196978490926329984014758780295522293335941389434837397800463249738568758545534885691463169378760767543361707338650976;
G[284]<=2560'd346640168219941423440988578396104423301481539449802857828072237613142319219053929601647797749302551322723410724669605205868826654722004404641882941704886196802133294319660091387576000785252372675769620273959810566613838198345547973166811634210712314730790524621801969710371264119007869411731703426914684768365699478703876970965795874236102534359866645088235844016725795574074411442640960378703326067820707126659776717645001182822625446247803692925801450752642460711377900437404074449107369804056113823786597903153519328263884874518298521278094249492243232035576679983679021611690308978628490053874712688405030396945165036516332731163641649252661516248569509804585764562474528427285539974772027938801934551346736290822384458631307610349157187128871852807642983219686753287;
G[285]<=2560'd373721431362124347147315811083300081371909784719318700913771655560605601436611957779092833304158640157070309326555537447322635609081726979788141628482095565756166985381068023356502526014204050728990460763670842476444244708245024563735308116297472694814990758187941658269015728793364311555505837576614936148720628953016414633904466658782800323609844154999708400226254157174630735365859050714455038235300406222203131958752643349355368737472355717870871871066055875264434821180691243469871169120532575566769055312517309442180468421265067649102681094460294424936177422859312552802169134157706994168119858130440506778592755907747962973104387740012445813082052417973885824700432577991174320021994146391604090939432443188875801191616779885087815089899926701437160024248936389376;
G[286]<=2560'd375519796492659931924689103878934168040649160381747487687938861325036711822610886641135682831421566998159978053986320533553070658359588374738642535909894970017282729321243620385424078034155908460136200883953777664097027243730999661533388438046085173075770957989269014502769471846201737520969337562952115274720104346092211147499718757276765782942107702759481148261191316162059667068695560921864418037892739364528646834578630602521720081624752550728141379959203882712079161276933199971175249857660327923627176140483657985128649760473959113261888932547399212337220407902921550084348991386257208302533625757457463848021455792865405340228011510773538101657182766096789159338178926569426713009799386503507069991070272071540676281316140268353754344850988814693553599765387806548;
G[287]<=2560'd375526408129169253927547093925976940418107761027565240581595152154469300065050805907896611124987064866206272089334022383401282992195518244198611474369284763476946661978244182143014002746638880670967854573410808900732338544526253774296211561890780289605955600115986566551835874849506019340813345168992269510851534242545416969818468898411912994829147532935459167398965413905361840671038850386373076316725310708860341686496094764823389017232380276039130607389608627815212470244256430826470634941368238496964068376733362986010722351160825861205670523467377835946453894587937060491560814926489048485790256874471772574893166168862361754023038045383880981594811767043670727293266822702971859669829885379163175211269913123418991224844523980442641124214546100720164417571813667636;
G[288]<=2560'd346752566141485464343242665695923824268393373271121733154215036415188150942111237476568056988555651502877292516566154085675030597451940531929561151019962591856081400197499188434813090127755752407478985185912082704958526045490450496172615854134765043070040174802726516823701409696622994577140524091967100593695286213935404563909588255378585344955334379961521941291795599318146601097635443666797774380479803082702967271485227572673864863232018062104129841340473692508332073490680335845438834735389686970476617146565063606128344516776451195915115886161177030934888203335921009403560502864511979364826672174303685045255934832397405640887609227234827631422017538399886280818982058410149786524282230174829390387930537479256320361267015838191222832130450155406652940355350652004;
G[289]<=2560'd373721431362124347148875644188459168398915927571499015997451226209997055906817256918814009716627326935660996909025068783668568661264818528109737545023349838709312108497881808517610875315077102866806455656282182622867159621773205120013674159340918952266639154211703449866172367108935249129534701496433695974648463547385070058330865948831677421080417329874530866676392928063595284947805857141795631461542431000010866906869410227833577609732237756191170101452118778470493287576501382431627149370541121698987206082968556190435500160550373580335372449243103484906907493925033038841957875158047034206102096114565088907822010008369583964384955220055093304508193038326147156480505318041463901712559953215342688304171190954457169084196441202122427142802539277079827965770405733203;
G[290]<=2560'd375526408129169253929113042530298889789414982076551930409923439760068482558632605409088302693514892441681899446549774963415278933728174823722718733133277122899925408933200306429203324529774208553795836072766482884935256296646592601451516340407307287510328660532192014204686294693703237492755042186196829262131189339773958437155201666885207322569984255419163719408110157165959662529328158968329878530969674314401961525035110057702215433177642764431926021922562973172388655670355180171115593900576704401518128611247899951110583236493759097901609846858125425702599307922090693384160405274564640469965214352853474146288868734337715495623407051449659263710777081761477175221885568237414413200374534204160464103162698906228401944356186627611169387231773751923585379576584521267;
G[291]<=2560'd375526408135474601880956561520521519737196886325436384754235895324169030419761988665777073679377503397863365000500314179856839278818258852236456209745357574109791347694505947546612741494001113573477244016048691090551571148402015366277436221967841990349451231363594949092508342610167637097913823182453591819743663742123432834145006006849178067448745847287893365070539403770353033615227788248206245752402313832896914583669903408925381475896483315599167589295581679187852508776186095050920406230225082688654425070151407319823516393368413080015441510878151796925939132181684560424542234523237126457301491224043222146040043131664903305496838223187765234208896767804176770262446477998975984108732851532748587819597816292557092793309817685941516003964956321427565808392238967650;
G[292]<=2560'd375526821363150519127485350980216382125986857065812555824160204053813673185976684729430719540720812727115883033741012718423631070949418756474964988463660424895977049371519920357857431938322457214483751608971709800251844880473113018456598191090524687287327051083366419554009147294276221383185891512449670818739002823833796718976821554780375863089413857190730650145249048145067859929811614613724333310628566757950105028440238235586201014430770878956950307724126193185467645603751869651609597261867181980354464632313439806058325102203249987510111589251259764747541967802903133155882431037038854735477715992162923697149266592144561477819593051302154611328876753704941176678242300583980200443222250179696377005058944232976077237706983266668015207679053771634598770250115148624;
G[293]<=2560'd375526847189855633666559015004202244124685344680385286986908383510140360225359778383926600932986682321432518024195657998733254571311601138885626025487105466667033324887713287341064338082346473038203208001683532548277007853417794530552127865957312009935926957029842819875057207958793591223400182410379062630744912375996286346595764920386935924647818052480677703445172306084979079839975779047316927764803536327712249962879786437287870577836751503167937633065039484773980870076408247758254265520475007446235604381450519477738896696205924679890065361908690446806694768636208643154491413576648720265490914546825679952177358048049510425877932366515891837035614163693466313678732028027854173951844096633233819220279493721941519726738860870072719499360753542541716231090047058528;
G[294]<=2560'd375526848904936542061070959929113125243186798137565353548021048829967726407253442370302010655678350364808738927299958539513485699262617651380144820295669769748673247307688971112162148309042557400011196690001809683950963517309353977788955233674633212980233535279697739321895407972240450244800389160939083301065222471205698227064185071808386007682375602480808963127827827319258723570115682130744722535488360548583472724555560929212270949092463344501576238891435410943109365417600326084782615623763794952943378901189864082705977082980265908197387506996028731988384186730335957227184960210196982169409659559792641263085569430221147836016370493133950710215736849604800896202176347209894759097897391214147733628067224751341549972324253546434835495634796314995681457964835025300;
G[295]<=2560'd375526848904936542061070959929113125243186798137565353548021048829967726407253442370302010655678350364808738927299958539513485699262617651380144820295669769748673247307688971112162148309042557400011196690001809683950963517309353977788955233678694581385293626690807966578880572000045423770518189129141529182506889641914886363884940699627779121896113098559384576008483339385082980139506105944585763219514486311406304987705835490695270135178775470887535871887463285494505537758708682353562861653222269689184345862328957696784531518207190004650934816268860071320037860839742985875405788509499391853860731399407327644136907457452417018506246839689364471676828783293391568566536779728445558006788436703616248320736729443063562580835710037118991798002969599137251493959992279347;
G[296]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374651378681544973288907532252361076013666096184460625399781827169719148772977610020867833935195026032158838317745569339018325945531255002668281394175289134992069567765219803847188262940875447481211034710193756054284083414598378595076781963247700374298336694176296505078631449050348818831928461717636340065956134262017483659170151933945715108224488681419244071933931150853042323265650978273513731356627087126287898286059351509987632559140499298677305962929838818147595068890991662436475534209150685066187941648807146812574275743099734355392924225754987579665208658400645453072;
G[297]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657039402917386276938768773586998417597159149295475539205602899633491245905579478605941723007278097492554777844616307919064847940564548905239597325536668520282737166849996844511351964826138914747640122895995307320016870068502197036245286120807295476568815801598894994276041037261027836511059993763468117425239876393218907732926459438863983131164352222629781775799407383010481503767578556193448632884110341213930884539055417183982716567472085382810774105605869408473109007752797907430731421725926151122437824997318661331409208903707680152685148165780140389235223615978646784;
G[298]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657415310196023076925218073824657327233206299304039806276713006698115550748452450408862943291697040146065178922830559647560969230955197467482495859451973224166459711018420976279694516823698429323433530039251591952575900210307235613641752465367851727253191851699472077409305280991582571120795226137069389773322736672190261405666787114976557665197863418949667621337990339366751316000811626871960934573522331479894904366433421361869381485268922025878625569448553630149009730305105886991972523666412207998587243199138503237987206745809923012982271764569890465258721387882486369;
G[299]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657416778583830251925165141403710682348972108483760760444959530553836739439244922954968104308422193732422518963752120017816958167695556549816364270565742410309470784660412881889681199867100629442631847299548386998922026390361655070466133948825978186902654570632102772689301682343569086865765406792236428652306369554265815151318186400990111638917134098570893080747479523738592761982592396804419497563137004095859950674641000457406655072687577916757231629033555527067911899491646265038676265057328732403817690636942162861123360396714729010990816811272903091609242289207268147;
G[300]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657416784340807954113454800604208751712865204558928267058124904247147456990264372992380310034971286143486938080533102542529503327138947648814757532578551161019686048354786133786222001384160223697637909504794077060264532835110628172001678766657792595884410835988962785442484033862763246259953755021406557369516173528710655921289938212232047277381545929758557019142581913197999673696274658008760248408734324683115655104846805822209271418042555022580056421488016602067951372133531777161637441893156009484039483856886812587697160892150254082630030760821250750643413001349584434;
G[301]<=2560'd375526848904936439835848580223185723368693707248157100082245105822457809118348087590095698571469869739337393181350835846302500224783686911464102222087831713236718483888648648631327416695137378484303943437167632533436369404056353111333448490539670071129943162283606802345088665745048015127786924780970649583853589505013895673343080842715588017591407115222790310215133293792928570136926696205489051728739569848045865499798068798311719780622578545671205391694619176930945053443916216794194576575640935047724543922026320256350274631671775115470674585182779188461636508280767310479083835752947860029500106679091560263950992563802132672406775920761465473616174596067817435358563544241283821325856111217832102198206781047347664301395876781295355680520868178809398917750913118720;
G[302]<=2560'd348445585661867949275853091035897794748149839136224171230578940215639490914454518039843152578157003246839944395160268608908099119098937901568080856375832185224327245835263105475645818408940631064137985811401507183319003828630070320940670992538815182664927142209200341533879712428861603737489947019917294894079407954102091039928873948157492963581443548492567893982982356051941992225144188123257489009060485290944767822471287531863836413681645623054904008734210991128273930638018544563640090339685999565385101480400222529430565001016634400841513509356451632150296292280938034492404634630877764736980979315890165616368472431826203441893118936315982439421717211475425951619831364761713253575643663325826845652598447060779373524336865438615150143731280742889588358762053643376;
G[303]<=2560'd346647193090432010267956802042950034872640746146855908410108296943834601004200864980790016116858921587975876006529338458176225161212403691009675054665081370652454221438876407352801677217745456613387348009691088950666360349550538333011341841793823262495258206632458665130329923913735046728859917565057734139732884660642238178221274713474142907426250618121605812760024984851743789945026985221518093709696053546609121753118067284308696098338398792181791885601325967876699408151047158636774805062909631684107866471220203442898486100405168062724175444223589038196604749655612514716518143723221536677221165708515203073184998066923632335357761155760454625071730899649540755308674863195176591697600326357032125843163380892911965153724282013672871182996847539952878883302471343205;
G[304]<=2560'd375526848904516185556003642638323394220460995529563298783069367865548540540349160638377207829113661986176614353811621435524714399916059905156634154703299210657778061980939040198585328187201013062808124396403385579164021550406235405817873845010591771897856437457259832298901923178256853356240608899885677067216524323191963235612466331177598795013976185570779912942148109393077897140686259594937430375554704815254823063487428757260446688405317079478717470452528636146863610583009837659453994256362719140015621478590097671317771784533191650175625754629408363481274786482103853738480692456232234736253023019342794975734790470726605526275942391680070703455930780853629796144267402489074736213949005991911391054649860122339760956788252155173927901276154887559840521174484821300;
G[305]<=2560'd346640168219941423440988579889146211111029311278590752312994453994577135627304058425346045531358489929099089460949648771657908088388276447827388096230993387996665576942285140162904845669076679144082551440924803261203120529727031550144180410252400697003679722462655927700229138830688619307145970714505889190260167892611803334569077628999798999118527912559814921104423293503369532790182301809001769278861922074724590017437709155499938523209608720739349071930998661622215119982818015656217160796918451149041125184430656280282622721884277249966595877347590721555959079009776111936730352006166178532393694915652301833499124234522894920215025044807607649801645544756647582956339970950220054684215168839090970174249005627237546778084555195646492754499612590443539124935773798612;
G[306]<=2560'd375526848904516185557569210424016154361537013906935453260438936936445110651989038083759123860745836583806238287687290754724860441261589290052941820937719859614427395109211699569844811125209627892307266329061090947079342164810385520301054401171004877333155035255009624974596020407257677440066085636816585407049769528102693667499570248736894968066906632355349270242131989853521229533754503044952323888505828428890230910040296815443317085738834319074833320262895604571372431012870338959089498350239229101660937079010932181776226036483720065908327487847597036024183673239260232959550667155003741179667665692491338446566745497368985127385125091823620687185653570175214675605957491090420487546726263757228966476187644150886711650583877524631031116201890775994398784957363296147;
G[307]<=2560'd375526848904516185557569210424016154361537013906935453260438936936445110651989038083759123860745836583806238287687290754724860441261589290052941820937719859614427395109211699569844811125209627892307266329061090947079425960239853770036559982984385467456116524404556412408359775083834176693272294669442183632555229719434578127044150689959261320463959677189936808156472337284582669921755904406810156970278640654458130389428211363370876306953149845264023164833557099384472406240629086975014115971819144211885174261202435711982559776852635481429865692633411224340531386240649435166748532315138750767364784608730233118568993117047128546099487489756895001552861479218136295005469065483952796288394776448079727294381945963441917392255229226398973495563490376116708336716125395831;
G[308]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723047641974943817133278623886585272814067639075285614971820383723164074045292231231462044710139670073055070647604676300152927754721684453797438305567538907471867202414181885530215426543722039371047253171835550239111731494467613664552029369450720266184134684662980353364403277553696804778779132330345287988684121520232463922987098291955588043244508765607847995549332978622459149880434332531614132460930553048264279533994686950189444704395265945059760282060303707359988458486018557038977384667825297946669078017425465788623408493459748555301717432;
G[309]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723052107496729862771239177481630005718846648118712958013050939669416911078729221903567595356438561391772021921686877284936732953553713683533859010177111371927686458635486087837259074930031822078156784921774099477765045424112310777406988106209590620258513102241520343523564805679367935701786885123442897082851292310343359021655023975668526290037319771221771776044698344646350459169777207587404316732783000392782990835614720959041136458510834527174229636966160218705708816337736647521009994814436017885909635723445392363238809493953652261277221176;
G[310]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723052107496729862771235061177759838348197284202993201177687066269862770303404057392443898514647609247072966191596754797761860573278479714104322581552656585198353456918961734055669536790294831364476699297219477604839034674406160610354342101736789382235711467157564832497110347588636018353568914030902892610508978303922609837201255740407519890454120617359338299114073807393176900651909508396956952930053240836125578907110692621964716837593867075274367679850155064465214370648859287136372591510594936232757263878883987479464820439160426939238982190;
G[311]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723052386591841490623611453870657438563174370053109572667002577531568320968048763020180154273845619082618629380564226211690435244469367351423590419871220667266970834424973878696771591127051561432873154439612586525037517096389998399443211256412901619855546465234714211136371514609737617441472398747874418480378650530842482186453700831188746202791929713950839881885451842957248714493351461205783597237054270720578342738441831138165111979791632901827892493633338643745707861532370754612041306198518742905773792238515446056540038405858310385901900037;
G[312]<=2560'd373721433077178983659774043465613524924801110993599615069992963155275820076615329483546461043819793951744042388502183442891350633694048281361477292991525872657926344144579898310437022143955696896366026922127644232094721293202169792692513985247642791411580721287692795094512308871201313573323488973309438302500259468340161921149830438881342548810943427194346022056203402593617091337026873782899874401535266454498896872089472856253004781580114241165678283343465855848321180349819789605583738165087363964568954099029458726360047846220685466188104585336608086870836608229043001209542299938130751477964980172125800743196191202587941107024679940939944254987438836815260380180782490596554903723616496558229528050557135090554528007992172401917454911788853494198591718952745313809;
G[313]<=2560'd346753005094588486669950423090141556831270931236587125728652429030591608673345959649455955031653811663935251721904750449228090575450056127101675945172960055888461685363580268264044506119840750807281081761388897619368419335049043406834130895894610698270269769161090870688973330402985541855085352475722969025000818535565406556830557157813947815233223762735511540954769754839529322040220319524428675555637680120731468334300409183596759161638829938988547381162408712648125240563404603767590468296055412964293827651868763644635916362592247314272124284623804988464507188000981603189993098272695251365251176740311324143203413323031141594687474479246903753817068954182580993522079537960998438902233041918952060217216840687164484318756869319992242902485944219172964622790030748050;
G[314]<=2560'd346640168219941423441086450276847843280448397878446792590461653617842175617255904587188902547472858215744061801939558330603441485461287807182527293142884159101823060870283554753895673607655605912436020269543783367467791647097133529064074407151573117042646606905085883606823380045187555678723680679579562803448935391735558383591429425455394538786520034605072689644732490411160447499794462515893546241794947868384896336299654565257245550149262099655998730497102169042028996278067220784992976891196907369152346282674243526188841944597236624354454773101839516737818781608821115180028728613429214872851613116755024118242612120136731854521316425134439881502123118136101141965505959363960093866815483037022364575421059606167214102626651403350046428313727525681139908817967999956;
G[315]<=2560'd375414010409396346732629519626342080899058358993871893160616322875534162469465899776576919288616632551578269200109209183135056948141567630058938527281332722272110616959072614031629531376579418439800342801610532554186712003497891829880739530037215812692070587435193310602965401489655207720069408626151812429832963720252982811187524887725951204819700581383676497087019500144762939372633856757179644229107349380387455863669597079327446704620035852971639730696996872383804767960251616674345601117013274532810388601517987104021227455416644442113391441927377043010696711132331306483612485648346697046214095045776441930478060724851917772448464521825957788774391874281697877140970461708234507039035198648164999129368798857732216838330100723128739614158334944280592645054188763250;
G[316]<=2560'd346640168219941423441080691702199335269302910639842536700458005944222164396309756752642879434794206514572032290904665845180323790363793555481396649501267759562705865218498394460832823257968686155584401297841388683003465787073992613012089622363407788145735809484120244301817049590691043170228152020713586020510137609497318889746450021609580376500170437274694148590083415418434832647042954451302782390847035313840995138326527338296101133280059138939314224657543842980133709906860953706035846389888629301867728621189912707555307292591012612543318914871487663181346028017748510713070389310075986373683274168877555357749131345149766306035826806573488913671530078288467162631027582014304413236441582544335214610320005908759414676087857644320322607736437930616089235014966969424;
G[317]<=2560'd377332266441024674534038617167303985585244482812850037864277405454706906936976060827567322522515847482713631764029872220365961238084088224477748256803143548580879818416097378953529607283064010941887788800807396761176730376592468896783202412144193467099377816342359056172163281633880165342604877886285656525015890761329995639098286429011090379494943191261367212608517833808467068225120630835995787715088206658001687663449383568434877421950823754890067076949152201831550740773624532261085565698702696307515517523173673209217699121617813531319638863974336542690962268556735197313854218745381328097710055792149791764519373760634586753657851838388820063686927451090223217865362050788865995003530772930773664610003450671668403031470197093454830276622929149971537197466346590212;
G[318]<=2560'd259980126158256635406865026139233666304076468074305095169198049654743741651397094953947118451600235760294816559249018872235399055713113294672479368369742651644303149117602459630681565040709667717971939391900074360034738822999161431055795162220350713652074458878819684623833748285238489363611154500289767983361768241034472035920487485002951817081881273500699599762242663168971685170457385566076741510989426617725016899368838419737386848694780438810272967072510186519730748321056051679406893906168173172514425350925482073336514346282717304278813564940831046970226549979491771743022925071420018668751731900690972091253436052256487803078521681689591422088605159563550733749468618114292415449857487805653059304908669591610504419790829727543105157635554635299165466843037315175;
G[319]<=2560'd315941019301637840741606719666406898370318314340297958116507573339952775406228458391153395459250582762584154730155643843551876890452632677705620977118662112025236493733768952927130702545747925431295125757531736825927544269569722923832946344126950097332490215582399251696040538520156072621762269372954683408479281866713268152949056611772588120870756657675114494324868484989443638092545212584134592762384191607545833056625965677764043913727659442988916030831092427863868166448530053355539351903380250578657581567654106251023967764798756807623009632303725622229073049735134146559764919349722069251469844105835348409142807007062033081026483547050461020415162235295767316665553949098958968815971386788052285097269474618754722636014034361133543245480516268054674380482746205040;
G[320]<=2560'd375526848904936542061070959929113119679899335218837535980752748966041383386215790409472540008891051625765417479546745746262134113710067793539858982358532168704980829821235471074405012705906548985063812969361550487283981037675630105635799696843133416296996319322761206215587210344018573302701787178724609438997401854599639298057041743497564706473801999298083892330924111559500017281958527232364289045660260654608601705172991965011394673953779642340681262933582337612005157132188598045352152523375309955972977164892251612680441859963566581388043185519495145561341647616756609350235336319945335656034597464813086946654171203608950988315914804170082949224322127765708583237474528729053499981908111331253927734227055769684720504653723099881635396722702515815931061596905623683;
G[321]<=2560'd346640168219941423440988578396104423301481539449802853021465094361192219946495457141142565033507453897452850181595683976286092803514052172074760706681739510818511965200061610304617990129984846043256177511350570258251860640880652062806320583015061806607306720560327927678146059150454415416736147314622973561432764072563359422434596608665527785035804915366289212138832653620871501753822318006497490525815686902382491329036509812759014086562595115424139709060711614487732371136761543375240319835370715958140482142817962602704550055219524932831715459181515087731047335403964264810513916701825419226348017738901395820901281440184819306088236508616823137698774709479043196801944794124573324736612683534838654435454115462362681973731199915966058616792880897460701747695179306266;
G[322]<=2560'd346640168219941423440988578396104423301481539449802853021465111213903647704711709828827940022100936906611478783216268957939562764555288225274973611746392107185252721190639162962180130164964029177284216985784244453299952104949753710335492118381791155131842906935767485498729277712287017043249684757671387459276787418233663991592353172852986355538450570825600053759930291585796790995671951207760298035061458210539146948426540072875072240666284227243023702372066282974865932387859311390683192190995295682746561970317698185509103136405238054149203395383794356159946455506593779298837038536864235005996237489822844698148403525154519962307860908577801323565385210282856571033500841691256443744426974331689234215901573845314542391869954925090227334047745962270121620355321807402;
G[323]<=2560'd346640168219941423440988578396104423301481539449802853021465094361191148479959009337098245242486631442874245980576612397687610053193040420820426021028752497047976680783540743429987919403100002450269510362213986522570622108902775284739914934905919306001776762900270396754856194035154215714681515312643378537579207795652746400795811399851342512817109215014537269089309763844835099222047246867890362472484554955183396156267984388925848147149892052950654319418597765604801263742690053140946263709130023340782575987191881207227708671193751401131362201353931822561450797784321050984334944254352718186260151830655212088882281641886466619045571081215145932957328400865815176393177890736305714660492463608645598860148010755101835071559679226997905060604997190238873542298473603841;
G[324]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500282773366044883679600277988783080328995310218200089877372429646475606802734884255207548651553430591519233595158598425864076146643599585119309746315205823590098202634844335782132701435117645960070280869337191146978736679013038041664194722638845128531933714093155286445130949464312190849549750370006781649315134518380793965947533579202329638863454760271761991347379013596704377721705739169415432429181549480307470269024551257567795895257127176809791664667105680773746252001678868849689136261350204269744661048518238451588732412715234575187525484489075654345075088641109380825634974002069363988789370869215449753253962345886625085726859536091978316005378868928749445514547;
G[325]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979699112508105382867755088050408990184665037417058460440429474492645488999355748919373060381364373316207943159628206614875076560219440309328276727581979869315180385012819741960925185380895340998914104908715704066102999420046604102879142903973591471352937643612950837751330118585455803687330260388047502089502333821476021364995091780388390353205108444819474592136580346234316958360226332279537218233389572212849977683880431582668036393847077671527441663071028162850164524743034383787426415422533576529409945787139819878214874927741002318767662539548429936768742511936881189660909367968127042367948732845290833427699208751572;
G[326]<=2560'd346640168219941423464477829862029498531691690635577009575698627722631792078647363085263079588409114283765262656054865106275795697842053424395408592189042852404481499917277659289075291717724433915799482678770567422184585568855856127823342343638569452218319752471314986026872751617862088843989562149607280589473722184439295330673221902545745124288394044657617511390346868302409914202413576426586838521510737033794353587470586750853072309984164636651029780956423522043063441765605738771074190646412091908546914536079492059956911902863128050285549465669791208761106846875308403704081093745889880616758716404124086604056411172557302419612230713837096345701461943183340478997726570489337289654095030992426572284870869923008089185175908786875225097037763551422769848701459437750;
G[327]<=2560'd375527287958923489225323248330674559346377387611524711638634604634970123077971587919760833476594695461281705758322779919142833332497402043435836023313169488676931035304276958499035353136160949225262753783569358694867345594133357169585681147863189005366124658613748796736257334697624939339596796649348938341023444674343861611212738746939938521524281693838987960777965479358136732021709250893317888276891150828999133989812944621455910053175507442808374763945233285864286781541769572062290049813973322048383737088556945086693053414396550589844032774025018940179950313956040778532601560017290843277244567726323892030301161205440208570064766907258361091524555390409480736955459067620957278982098700374786965757084666300050083213769343149201406035544775802957907459189518675302;
G[328]<=2560'd259980127994347679860592485004220513219339050643260884804360016519412004006960913784636810804791333507154208628635783266028628230259512502548326673147421380346776586409466930890958266309055334770110689138141094551116272496008570328131224747198448100145273616212045843588824344111250022290669430793377486856382256077828058980814187376303906820812508929410868783068750313204141300628675900014067973590604335650104205944852447403275059449687049271533580576308902639136609313503016296206977045044377208168602945391892247727041543536006343464687564481371576464296663203331754841609028535947021772865322338501495269859062737198975743404004975069961362994070416931450407046849650149910794442488483980900135756421899848170481779541525606293929581439329064194327532021724875896691;
G[329]<=2560'd317746435129395399141435557912922915528349966869745531896178056794216570062245169126153431282803090798434426217887605962511144850857554686827662706009533631911208691926827595304492300910046310621501763052736004665215142337868771377624286612753621676901750661214658646746348787633501367745053540288240285474834442447244215202891349938541259508420806375538855910476970051852703559444908954335596460874223204840103450077239624768693707703279766491187991001794740515411593395042468017446407427594961356688171139363430336202476313489791148366924625336391017611217089251856034387546278705264224233110016029687781792841108327076396239232007202271307071319166538794928538364779084087819789011835476037302033296320809187152291003986808305386162929496211804808485326719305517504370;
G[330]<=2560'd319565957490035109871043584065289681934422485167754676826192542481141305833073855039119864435517249614909361964957356725230637500220812425243906643748540363248596504549960062295154822148483878375515465197934897164523129299435085806695285824135897744869823614970527102557583381715977474112309982627812871863902671434822140780666881572988361676477604660099866912088149750953260486228403953113472636263104319770344395240118525199447374295416434649970553400602873166156972034892273898455002956337732608121199602242429411192313774929809305041882702707014700975340884369490720620420811820626699246897694871907768577198259692984960681568193678179293363637852770364915126287239578552204181811689055074568575486229754126097125859199648683434543495531928491545054205979102411457644;
G[331]<=2560'd231213364138034241015058140100484796374131443742472390217035448534456112496072872961159101447784732140566130633039000340623129719026467055094909058685300602162580624333429619348088780409114397522121000354162311441543048340410660709353776568341463975184591528256201143628690909740014700215389292906028908381586428988753962142259298575654802147287825902078797325541455018305971637941268796321896883631502902332321099229777748606965616960690107610916752723230309229655365202539957053062562144755282860104858285033150853909753312977112444912824622768554708899815906229838832918693201300622951775096312280389037862964190304828712673578469007868709246648042232997980183832071217928629470577350464011996602124940243639537434205679700022606600704690999654489302287007365738575000;
G[332]<=2560'd231093473142809652519523677038597848083139368407209418500205612149754757593385154884838765098567465601367013585000046926510336050548163009564920088799203859748031568393108301337531858587748579102693570737369118835432776166505922427928305051347262924033457960198119599039518308609990930412394612691091576231986260927679999855846865383453187396553880193995450892432294219832448305393237558783263671327427086377645366377043617945443613054767241130569603458701598129417223773753704867671036878165324638910136549230712668261863550364536477569531371620412183365081675871777889484211956816010164681873300630640832138709036218642257068236813553448360136253577671019240342725545158786001626328187925609875371780660085572374100823202433298799665044453215967328997557736583626582905;
G[333]<=2560'd202206764902605022391067431222359007799262993461919324246545821611059319041744603128948280439808329973809388558080870997266049294346752451668654419565604041973836748139969024045288101576186658685711930412627214143013602014883711051258196630987556747887041772363014320602269990752844265711942885097616989459559037907216752911218529127769768030762764973470811481417557002933306134943535577300215441487167107163375951461564429106117986126982827900669129128738474908651166346858160589748121681885528295329666589650836837959839079841688652123091766647579108608939408818970409683038218867100721355927561076168176395755954856741609727424984269247810964453829154269231699357460284420769909132702075946685603426628212894998844262990535486647478359866939861876665349350082537105340;
G[334]<=2560'd202213817106356880064049139230372479690335771558318542245979225956319614209301758826160575330499100989788001235206929953773713185979867328160907803062047096912555999828486132878241292260985017789540409063100926103036660140401929245755641400370242440156125091551092802482519812065794806622881987385726258769526767018004320428917197279353854546287156599475063367880889231595918700997352512958287019139814420858686155498856152081383174147070766788115435372317309141903173546121567334626142957994969532487551884659067482816924930654004745263859782243555190332796561929349080778783238893397146143314116920703311053636612218354230889153529613976715696284005308125815301328216916124976192484539388891409682900885773291587514537345382233429252782786896508350603510545315804239271;
G[335]<=2560'd229288029658953732121682396643270210793679112876287959704719155356122284956587881513729214842816093146060917911438725994345069828034162031524460514438613762093228769251188881007610297185265257026896510996058254430297747611862890818494921260346239901106517374359741597707580276940232581409497188374812564053979104936738307736478233730970897493002322161549597770602096764598844740598625169086293686868232437090739647076900315416592421550399588267513878105497514951115515643216205099396223574154246994860798002262083824437407881455439055700149413245778574405226799440899456448989445048999485773242607955597837203044090222902113197872457644521436584340057185107379282292052373502523249860967423218123654846296622914977522456592416072596594318858743698162966153778706137303144;
G[336]<=2560'd203899369568477836766056595285055287061327936298050469777005617163204429617265137685121957730154756481668046413655476154227019157956216510248901014202679442121094540461818008755469158372462371094647283228048329083850024088880832238517561473316735167430411415727063286314128875737258383907551739696970301292879479324146904560595117745576474463908532994172526150437337251949866497972035906395605524898297812633730740453029526071019667662972978742793962025494066532782640187258299866833652885659308927076377945145480086841204990552454186260537028579376925642756581613062112965934542410670585875781150217353899711626913573717640963317877331203208877125700649318839828226557496137779156504247172174141759891444585719261922918600461309615052982494283103178983105965029086231201;
G[337]<=2560'd203899369568057377612861736895361760200859565282768434459588093221777683577267322315156621727125531170812870950486435560203050371179492722570982094832734265230081786938662713465652299557145522651898841177148077920696824713021489813912917425931082723285192833869280756578218704131868702755522857523142473294832868550546609572016395388354486051730494008750943930411950109959841573747886553609017318439774010906545937247293468072096539391611037107748013891857205839174558770539019612426228644062088427900191140131803013438970268525196059383947144158095268961260413353084274914322412254922885605143194749489978894743910853124712149882411112057044843877859905015821406339590494221164409449117040268065651729783511014866140305870615464949472367983187418510731026189425587180723;
G[338]<=2560'd175125501659508611091062783262764904567696519346202955976703954639031329085300366075741684755028344324125037084524439586776232704703765563793292582900517949139998618455789554993667354767436315485701378219896216230217526702842088462493805512682141646962436606619661190350046719622612598862943390910583860466985736717409047146281431233132844954978107097806695217957070198210087871057877377339284162854756000449107672893588686333725480911881927918744075394426313590315549977825794625488839900842250096049245189330113229763776881821822281182101575798716068155717652170341101887371928987027418358999886298642843789964955975562146524614365262326380578305104358893422912181607594418526357499187021836527279051709903080668699143576681263844838302926845510544057666374793623946331;
G[339]<=2560'd203899782795365482519411348736625561287471747760822015351949233954961550190387666658020230881197431834214667160287708251087276913909470734582862567757097604784719543222349049627346167112966524711378405315092616226042851684229190888818322531072280441926811881185853561400595592162855024136922278015646856165868074603087228527152938915247660410170112077434288841454093930923132579037332989317458425282698267119550933018732063224740366038932361771771361968432578836257523839830832128733853138767959936296589930552722552972291772591727728028612237504290134855351187270833623082612086341638144956569910350148883189391068982386263652624292195646816988748809272316637491130542047396803428677590281684453658948922854638921585644540217740292912715417139994886984226146349171033738;
G[340]<=2560'd175125062699681526300176513193175894891206165179899961613962716975545489034451908493261700491911628073648422748552856978655300583055143460590561633470758090458660263230849982534328759731442706885747021266315313311058862109341055430542593198679403116740151059520580630265948656736744968803231598565496574947447562669887884585280786894911623205497951507598621758249801484070485100457876508104363290869884216541797734088810922015720382058129322267463624371607130782553573604373725902688919647187721228847932648274981204418734509288567289926468978234817707863260748761476875847948132017618757752927166878677919506869574900558758822803190907650773224220112040471449427116501956434478701714633148487111941195127818865094332549785421061668717187410377960553615236212326975196439;
G[341]<=2560'd258062309079705057649129236559732929448858679835146770035648688992295325477182511194167091373109335367841203169153887884814740480771036109857506036165267378572634910339449846160554183414870101210686517197184239566157106901876084758014144859286205069037808504029675161960175975751512619869087658555052853481449886490933777550530202705311964238901317886939371800564314678406829611409488492697787924095655845328139475129957880297079970392651069758054962498820937479007648174776453122727750368734827519178908029955805306174504944062827669752213758127887363397481084757615506471946076546714427570891052746996251629829705958822821582190217360877679681453910544670816775076886065876762684259734111865720774352489777683301663703320189551404710869967230824658368870453298584197973;
G[342]<=2560'd177149074138633769353906881315947183979968395198623594946467349968799734255548500348790490968646930242862562811738295079761892641107257541767918544808954686351654154825194381375097541703955024697281519714091398650343551576210096634256780359215271243638544957257694487454956545109407072922795844466166781802073561908572952654578917871121375532900856402445098693616999251242434865950730890589578108568232428494093550384536019430771665222619166394374144790282657210528796672175274854368597724581648343673467709435192763021101015419607574492190764033034298234912336929670593815336706325899426463467519663526306659785377957687562325503891848571552275978274296366648668057335709841838529069075545666960354865770132624894232118614374957207054516087073703576400268283687054138979;
G[343]<=2560'd143274299016237833007690268197125428216797836150202233068653579675122025926587856618466493173159944219948666549879275945824836397778556224792857195600963423208684606341540350403281135100811945852765427374944440053632168955128370836609715702941158087155700676469731785188797950648638846046203662951370708752419496023667614578953341698768340345352062098471234766592933110990797401674671617774317423703364810800314375588129162958418073054937321771198795522769925049507555261959807760357622589451327766571198497109324372779069808075523966126216507344955840558983281005614013388467384427661703635612943247172742820653404513420135285302860447411713430712116780396598821674356507078974985212432260653704920654845485446951062085410735959100933898422144670865041840447336524438;
G[344]<=2560'd120201790053917272393622337381051760023410450845603600730654865553527868615055119926463724584758926560842775541495884199624683322889726253740389581569158835912961651449538450834428413262766944568670934987164711833745391815234276218528163205326849351348504820660059599436896496677007545677999018122660029559528561171115816791909644170420727052525577112404594939841140326918798099045108315942862559448080773755211092644160829695886629653093544214663676456686333146258540506041222924947429181212892621946609413358414236746521254266892696742986312232851649765325945433206115014058704422226648162369513442928502617211873266133570539744328912093734558940047138086909728556910941924324155391550264482201621538280242361051881023793540993756516150293297318699104065812001653;
G[345]<=2560'd7613497445223497781101466999057813747485980472406612769620292038473717438857983851964823216654939849034781152639057338441474446696420814417884977344693411405337799640288820660018951849486613474584561079206897797589700573349167294967223233732251184462196649943630427411953941268109214444514364332369719321683432636900582391245905793175708035048834850462940487468867184534007041553277755499693779889221113770698295367024348532364592800798041995460341355812742155116749213137441839772668747911836461109702839181286037178863147912664791668099403152270308862265603865520196697179843787575216647375251109921743378795810526715909893377905654054289697377798802892920384467401535174800160340147915050991040072316922649097893045957672178385847458660471003347858543728623897;
G[346]<=2560'd27081269040625732417464653287115421125953690598544427549292347881595370241624010954936334198933735583434565431742723273016187364091205029932879456818244044057068327877029397113527886685753853923398174873253328414750521917045592896310354932899830624278916874450616248198211112669718903952390670303407874076176353138200395727592392615879735722520424369069000977754096996472741616403615259298848904196124107782778789332273382688723490223673804333708081301675682221833346626751439826000759090660141512916616066326170143461687222227481119852853317918261366185216075484988260041860259468959478537795190400004398001115373299279836084683536513870384836964812330381468739915955843104365757568248761425916603233737798198128106584529913866380594108865489795037518543984493515311012;
G[347]<=2560'd112405434157560890358499200341965259584002578630221989362209600832654810079998887274370094391143277033420270463083097943596250754370119088699975183667417934280098664639086962350506633127422903861513531301419591085212698060581961201547278189605107794887339406970056654882713071899112427238201591719183115718905710264590431254528880318688470586668296183073605268047646820895609921282090550188666916266319130708410650502844697981446523911454444044175861954651309589356115892230753477405381776012568826570218509206522924658099801070432480047600003484376135277455356923383071636780506590374196910372164551747523426761876394704015122037892763446670743309846984129174031775959128023041153321813823892827539734675157741830300343289911552231723062086499038606017186957906545780;
G[348]<=2560'd1692584945741080180168639769507371137931388075081459600562560036027464137542465951709212441783832476976452891024543055661413835933783783520463065306862150747185748140199007552492613965440394164749546128799331221188278566034403950045414144680033652854553882558651633061245924852675154344096132661539665919076139441102480202832458516969235939283036497559300397325516470657223013017014798581676744675706180269720860930631773726859372507798941943594089371877539394026171782253312885876297823208381437555581666094716259621231527880095893690106297441952863114583962394476210499818373652503520732267807294166831872843999529729142312214839826405553647953641005614695730039608527824482525979054792282093348618306124306013640671082864294178193287527273506838625832435598544143226;
G[349]<=2560'd1692589788222017297576501823972598245871106886254788143216516394323782424094606953498749069192448427543505223121410157754810543037530461598141885770874968303657695295881081277349962684836879462662009347873950465589675647837912331472395730196558317154460852193154102104104705493770843532323665913086329441318744463016110015341011951673431897801546027970251518957452075938744455742416319954619399034231254999463935748656911299580421803207736572905050705221486384352315608830502791341276706036785666791995794246859329740606687225228313506712293574731353782984952475230677615562395659049658122883899080521401632998489386796763508371869563681954029811296234739606762361498558474650620814700189097135664467050434124913824070193963360732604902242901124501937928658067709395019;
G[350]<=2560'd2701258132438165946309670587038957502927495619238018910458773837813198137029635075074521890120764520891980739699612466378086581767556224116323269489490485874847910992605688940676767514727803946701742632568324932340261423809962499620051569180010550545138894801707399655602754238097078339960043321882283786584051075275435239551990369726687205275350371714601511424006387656896768855307734255700454040145592668147656694261376584992924544412286404827233336933419878024568253782783239910456193093177462752584902887163727918189377529656583661802145695460749105294070459439874815366182060547781708860029122926636650147058570911048654602388552314951652526765605884491486600637530406591960930913519653571607582672699318042337358864584435733580206143106599181558389758987776792;
G[351]<=2560'd12305564096907383965118454744745174241888746486041722538907866859772013926850738682398951830824294517329787788621264525507362418291483017471118379052291371009177380959824187825489366226326320796019203589230800926371681666800204962015793358513487814681253109336421843384134275440079506963730342598417586798390009030759639916119522867586975901460254017039876482220392793420760953921774508306204673811753075558722974700535562824751894285192315251625420372111851746007679123380672090248466422370221784098848981008679444776542323701059083043960282312550686785461539826381120748934765165721470546295139267718808515690116202268845105842601481473139901083312414378393064946347912600009724137736213718567006708225613017517556438602785109921428017359686577773019039567825969547;
G[352]<=2560'd3137184666812866482646569288086007109229579844593183884807664840349731007910793662576251725821761916990163466239305788150407564691365809219975892797043087405118356353718410857335600548286808838955686482778588246225835990622444497676163427953656089959559440724366959563390566241536384848493233304500703557166713426375583539470524998265560073510606419969279316824025602089547421120438832993031079001995891764488953366821292995068406228897764269895590411965722626127697269200729546787023497541995177775992003008942663087260014488839886005287413268713185072422240446893673070641353501063298077634010002660161905738337764260007897734017594604577587483539206164885942036428826275801698303915573031530295651371887655324460060967762438697583150264392781780143594822009308517;
G[353]<=2560'd3550311063078637993014447135988708937736428788978431972435408056776556281780562112183194344223706610489558629884629433507165033298303721955531596908043080383444879721292908878985503227961104353533320550312760803449991714041732177611084251507253388716081516294291549411510276700561902193741142898032145416962885768826076969233059215122439316943046726706661242302375625418968453070926760610674514233845591724360398064749671294887679712059596771117927663427251087292198336494596505907851344699907337114538586931516236633030391534867951016659181393180488061798433661893608350408782519790960348786082776952368083776647153641899915610910024631329811064076498651311305738290687366161847220883526022590317271830558573719279229990094596072939075232513621247886043249190974241;
G[354]<=2560'd3550311063078637993014447136072159522392602710432389950934599981186744173099271598362305211224496777713328191523732246509896775714719536969459759160306927677032986222123380129993012003130831161457203330312127740118501175133554992772007084866389991700231372243472776883500168001368838377291105890630406608033380658896997324222911796454142815115783821962522721882484606122098416193226053909976662454951128279427809712867188211357278189983114912115062159737941007424939723871970744878557405832080260412472365051430932292159419225701517618786712245004368492447093937651878956721789146357071224019500614896080126479019521152299230382181123618203960883559435485997771356755434289103254716873143427055307629929232712748788546361032222350445788259951053670141312945291030582;
G[355]<=2560'd3550311063078637993014447135988708937404825957345433452989312123858201021739227759742648469604645754147182459071368197275614832284563857763029099390395387018749419982418934320441202880814060550782080480533115876496845155411111383827295429415537275005271354011097421106307297675037651714593437422949252515465063766303258201740353384162009224402123692698357351873398265361809979364909473933103926205485909755509695387987718328088019704029579022769633949074485353409027999708231160152841682178970216217625198305587532911756359262760728397457543762586359973935670104743057946250428748952885078529958905452312128919753520301309794698514945693266135973558056181417440920272947375992085372756971139283596653792930428772592719498749742509962371154780998352030042267440928070;
G[356]<=2560'd3522870188894440227246422038399077487991688511324486384609522584568205025544895202205796609207873468725147419923017261708828699326661912471573649605096160597008166563460602052010205453719981096283456631879193509896212287336060052734009944774782499482433090609053158176449716280915070627621079482644645283537105324175973589073464090333780182144197410923377621388665333855939015877230785250113006278918700250824595651579533964045225222283078496829158189775666847648235471494120371381750618526402511723988379365262860087902485632721280447852646481758599842936436459787790633033133751661266445225629221483528563025668874070040855457275172939561924347038296322545767362973749332926199604802717509934651843587628207517041402146956246872347274863767226907683009912052389920;
G[357]<=2560'd3548696894008979300910445659659907087439347284050083621140114254381180679557545443296293226957260287489502840055844856415794935349408624214725856591213527066560112241826081028663065228752617347994779355386557503460726597010443954065101028830312997798151757188856218721503127251280291051798983245568783292602378626959404746486530432835085992412234742894258332363654237366290575919139607100266916379334041063542471533129780301756829123768954211409722137451508737034454009526819835408626983051980131503500086867809124433371120173419722043848462349281128611089526574433546457614040792225951083906789991335300021772411393931983331140365673154802843745177260327277283864093964213064216665719717320220960492277906667727189031555238998584400424494511966508007336537371984912;
G[358]<=2560'd10573560685163607337524870642605558137202533465412531957461118371702609577667444234275259288954141196803580509521417584578863637617557989557243157182562308611225705478326942943194848099314922826459307534059264484104959815336108400852699461539814732165932599077414089859626843526321126567180247484126788550904822924133721987613776011961672948334653963256156094394231227946858335165783149413304257354116235643020508268571919644030497472605574702293953841450362275470339498814846936562045020038232432550735427606966497705737855191543002967094422278289297423864310791113589685271384650435189622851540749018934589107250866649479439565396951437030841097964667222727441979255130520481110030053292855047898483416003021531329564360570841935419840314418493444106035518178983939;
G[359]<=2560'd3548696894002588756433497418880088038182367602582547460146395524231554770187800651632611413670330814170079905587996436024052677029998169995346728936573613656058267117786719679767236619354255698955474554756145729858085179547871122260605945516341082283960282759597932799747128435235071258027789034853359351043619875949293421549546313018948110625338876881956882395938014298105718673167893975224869385314146112522378179095763831789789715989077402605203893261545761367970900603017627593496485926275232421386312425918097361362817272713665860929829100437631697479123676114679945721137299220247531689784664401570893961978072991478058970012084603625586577969771852615173588883738176998971583250957725897268717408728237341688658028630117789706284622691541145348331268804247825;
G[360]<=2560'd3524484357977680397644003635615023943254120525215776711246447596300232328984564660091373151175933622165939569685771267841123534466550308144051771369911864601441674273130822666380833139170268628583142876623256703123303602094795703442450357166000344844227942037318474769233632329497557190341447969900886857633612026631717215026046423606921692297988251133937922054075930255529477698260516652105821035092363720871174881011049518940747598330127818461546070008707087335265234271832197771167655618918175190027067328492382992736970820339097205462766290653318570110910128751077312833505029031509396814460970692148188730371022571703576672880367642535585508729742418380280618749441356256428640409729825025509384575890411113640099320045794622173685943647863592891939400305348880;
G[361]<=2560'd4376859868590985324370685126902846184393011801907854622851068234864274879369362524481722797099566176540787253315426473000774618212299299952580281920747444662866161398605750620060866508016605704165647709202290712939766647018376706140353579478645702998164096369772992410035401904301961015838651617401380108438855215797951901605069342207370009995097217219836506283803279400806235392955569491403451530786826242528762187223044179245215709543936640795571250539318124451497593515474195766640490261916130516048767891029171602211435994244469398907135636361641795538832536933501217957141070057207039398988840058806676791839078822219492522789415399134525556630378338553695721491134011036099726123392646700355907401324000124435296153591053428104872930398347680130887695948849410;
G[362]<=2560'd27098809920412622913081527958890090270555593111636312499943103938055012136140259060448948384484900222148308879169244290092453286096193162113754022573233976040476130907337770356012398952243521160984312598178736392269348262734417794044288130205655063015808174790814538072742248724852498359840056806599966035481665838117912646067178650730063709920772406393648331329494667312192550187884492443858755736236952414555321086300399111689680688961122599483290901856327906610012824312077803457122853977461069114122273465368074207044579315738440901350321836416316071055979182080810905902963916926833287611559817006922033640116430619846311085449697676747208294157763900465028206024430804151281829617829242487974111686135245220683789922036912190142045474380373088394325565038182535169;
G[363]<=2560'd10576714357474915621324981377013977593336247741313076091434256614000551182353773535984846664931985636513986251677962104004875621548143434962562512807447099941237167671161660660188324210105096062495159763677944166319122232394258504692089556421582639182829753395783048385017478850953127261554153979582928176210109318355370472055201619578335030111984407593240021155667506965284846016899493371581677060805533565997961360610445010865612728008400111539605698118406878044829690594434851320171205627393965647491876085647880532644970233497277122519536680888658941775377301890447169548770105208431399177112311449730496402868900983990409437439374960532975193695690069941342839414886332074040837279419923343912486380618978524612504189773996106478144568532652960710190666331726080;
G[364]<=2560'd27092200411310148886147691466406486094798151457873300244785359417196373449680162702791701962835432321825688238902761297356736237540715895370502880446112789231690085879699945692540629523356485412261287728868468542478323432831642064088983787657498866867647033813520848851197102047961519415086635296186608753241612085830578931320224419614710287161892260822935391127206151745925996505649074163514478842105887054307053587033992491924724124413818847180454864249159357702898956668282322860775008481494365554309777331809767810275705732455318379185986852920974432054906252015743874192142465829783018501578026356651337045654571391220924764938900140037730332602816515761717578998615353569956894498309389257640687963455535967772927562030596052829684063563636760661275095923439972864;
G[365]<=2560'd16779892794043018800058536356847281845635341092123483811357697625583236672588164988191702785858521593240950989620340530087401582779048464397597063941165922330702537479712557871475953626950496216088468698772395550311623382764603947464416697111529718140712482342704821369724959270108171352077903065345846665867955334816266549163209984072547323521951217563698183358774423672472515107983833247126254279609049437433805819029731945132925695923860646552482352058287673773732068587305844890441193185907469360457527425215732405824872785105270411475834235564209340103039655734644507197942315627482438615737659518526611418404906159088766065281117101953842407559116685350808139349389690657642848484060823618775053898011682593287537638537164932104533029440297618664210049639916049;
G[366]<=2560'd1711852125079697282962856169020494542296527249420747694139009962828797297051382313486418101207001788196081425421589986094090261898597598298590352818155031244124813377836212182414857846276267671392576782871888213304977070184873190293046280664236218294752766989114681959418295158759007827977175576935030287270897308645487847230601710474187355485648881209820904533399971809475604394364554802358561053168675452044547607096257753611155007834299748699007652119289034216734283051553179591026878525036877980056290689138916340266430037701249858908669130256897338341862613064227716827102628855265736499872111653272575153174061054716983578994290262001777451277144648277564029320376124082940716399293662427787626604080109682648960357084223763454906423410647524368153701393934385441;
G[367]<=2560'd27110602279193046132221003166316809846262049193035654484283437390771407327040492952428298289840846404031684971656287893222966546366782906652716452058675608604616365884830494836378482529284858973159503827199361679427520269693867955027705287286015904979379880439471640235951745342978410348068110094588517294979858777525520824882903502562416151641145718550084247704289257838305705514553047819812006229178349312730174153200234667193461457597297990900430424643711105870421575787898555077129892910639888937036450427272205809980355676180037834084094680200827616289001675560949621972999015043602807159917472081843303974482358353162207591117475403955609059524423481667565596796133034480859748453484069575632402127524039966483648231360054710672879899657567172783914040499010273281;
G[368]<=2560'd94207886959121087535283553749586685319992172369941124020543116429115270087301361538459151191350620341596683314066329195680081074996787816816010562539196764494074026824389877695815908738722955718603228533886114211152854004439475242823397884604942769326043014986863122080110915653142657188904719863861611797898015426244210709516698727739806060168160594896413094473781793050105669163012921740262232924194156265652000457084878126445932843820134214408307513969669462320315100216519348814517031820020691290655731171366728034999347312400662900904986995957057980859991221543736471524167777691094504141531948724647577584644922710413951300001216587697136336209444912306170845521757988138968064185679604481892403286789583947204399049678403821121793;
G[369]<=2560'd5563451585595209175416538786692741015271238086729517588251877848071005255856161728748250345327796585628852389833662419682196769920416057867950624600803806184124481572319898520017260410073324961332437833144624621519081653793046553245631111811965019068609262133188440363948555808437457254971008607247624609212763456976230826641348067364798656001180115574629431403547708544658413750841052265634879237396970313047782845398201229590390515402662836321648401168444431576135760127261128509267375608250413083800195468495647036278015287413197617717836514179322643633568721065110958424754066815603675334841188337343188087175474088812626341614349725610985772655494689606070488934000884830341064919025937925387457649883728104952814434479493328417280;
G[370]<=2560'd1363549467393606278976008390815821103062068714058435599896488595889099501929753530770173431829562062706088175333682611897974244517513745338691196088264229149630987751957195085415665628832146467942700244644309988442750121121727727606553585463057024931961400749043110158212240610851094686455448343901851349091623361304045726555221936735636488986881044717512735388047391366483613781389322557929178801287297518948244875463493442203002624838023986332881543213841412300563103026311453438148492470588205223455862779553177670122405229445743128442565190391152266085084964384403177767000414575330856496167173162797781450457449852959933437209095024269218791075790522600219495486276955054119474633422526956979291351854017835295916494501894422784;
G[371]<=2560'd354903159918391446548098474093260125879838002824918672182813326543381924411288554847244226331211156275022321376137195624801437177392399008634648996899359966851329533429307105270284305916876873461113808654637253438933836765091684830408029862085958887809653124066466888540327120713798616575427554345775004075732044215196500342464912148174213945564865274466057715447646619259820124325849683067707589830816042421301942212784432227141416709549150464614438017751159812137011260561346220194047570877942670358239323504345202448541749797905772871598434655152948108834167560119466401392705886670907694274580838972779250493667512003855405024885018762649638219097278684664207225458763696783021794678538676529405271401653371913048438861734400;
G[372]<=2560'd2671564079244667609839417593197605206056135824187364182171406412902281836209443902496280711049957116598049022436932769006278204526236450097461426406178043411541084988581199708546454282297003685103268613357200669861128708124283608735776590569136179552904310701247921259321711241003094959725828291284100533823841702844368930682434827712455058946684978674745725499987877241605788435318339542575125573852270045603772100903263580969470593377504914495458497692072537056011459490740646818530293947933431108370073828090645521003549350116490091550208176365126445565979069755477180763774686718106454527759879171189163362095922652397531030175664553676538633799616882334485095989303038712621643506550417004319964872151627319118281962430737;
G[373]<=2560'd15811968010149373620696857058364560157395978975143193923379071207405439786211493537620895136724089603888334335972571369856062770780123405296581693326015012909969056777373971108676456188435345659721872592128122283953444388416365047349738532603214107532907249823857903184812714926382382816505564641232252532309324161530832303575989262011685085203314959415810682116841938876170532487358236853380772471441843308129841633205079126658043242523300454524575140776280035027847282926866753135379998995551441644276508067620432844101604642059903167350618977440906249562370078191404898604717285155986469981243288338616151906263136930483378163312301845787953658421809727223782587817807874847506981336193198317437753154053959980284937044001;
G[374]<=2560'd40842962419026583398267838919353303601451783888452366785209754860268773926641134330802021273555987269511660904093199555301352784077107657886671062296994262406056540947923359090974155609806388296902005643770944556245761223659808829133256044915606718049952438733533382146047604544415283650112386114431853234478778709458869093056605532798675213912953386962250840789667722889683493178548482474988463861670939819741900956054137109758774415371659781697787729692645255129333699538676060415496308045652887151957351883030547097283136374320006269023441797180782189709973277896558525610498292957452159641408958804254842429469901699961042251330473166867879635055675608254925454675552535689176657146828036647573934250796236615358362112;
G[375]<=2560'd82353202080926885845223337108165536555809296830591425626229192259091583325297743564420679470064883821240187598063106207441214316582271454872924369390769593810591020509355680085098843741966203332929498795068276874029309240669404631014072204682458135481538246574334677814261490172853427570261503113808940237395262759834123668948101652750510337972706826590501512681653556132496696844672072331981331908618073315149197780672114176052661371508277758017934891329652121668245213802055657176622975695985426784487546214348686524979681019954654757666238634009068133468339850405762800211430185934420469832039146958894781476265337691161335877405168203455612272347580377179552594952221539822992828995560096221303436172334014119564548;
G[376]<=2560'd4826781358949936194836026256926746496512253851588476544305925792164486316928721729005994448691950478722191114030035682369702576438773121323206389537163573893395015201642128053741957307091443137985463201650364503218282274030063127664305439837420368240068346985867789009626842859905915168660620652187564294688064973698685414092014276019172288094939062862256521428407034073231784142912034444697528726997198372972954726391258167363786788901906981185909954570433047057345516468440205998489835063746308689712070890567023830537520574597375354659395734882518872660950448013812119667577682579173799529753147525426210953834248381334315868798487661898893252195078710727504601981455238468452618013483854240103767355221576737899027;
G[377]<=2560'd87148741318084025124055811997096458145160558997076420112497220783855209730030143015244131987176440242786232940037080621032926921358047821726582214153591752748568200540307976019625341009074546911905089046957771266895631115442600863725426841910862069608262918873581028392221743505031956218533255304758802446281733994742422072048685367061586631060822378535669552596881305370080625697761017076007997127827342249983889066097378324159344540387757665323768970338174238224809500527636028862379605765510527971100432706340311888766250532160967053898861434650464017050503161689273990516346151833987286280275316859413997189801922581174567872891419222071681471119809987821921426549883719762666289087644571183635660840937533697;
G[378]<=2560'd18118912087321698212399061878847457579665563100085248362949864473457717304716929089247228164545746223665140136209880050906215991351561505525898948189465859460274126483485924118270924785686208126899157877983839420685414668115597800381114615765381926869088988924959267219759554809794512064442567292247172875563088390403240605801396696912405316124638081769598675038328459068772858208315472177039928990044890431585141424495877063378083364627291915983016897781643443977208463668087990779081401367915309582782497627797726132016922619204764252132133067240581964155748892791351766694410096694994151057874007912453993870311015930050966711979066052280268968473364427014108489762751382706439836792245939030141421466065833984;
G[379]<=2560'd18776132729502845738900953295118508527321617869445447832685640369894452072264650389360019236661667124568518698628886498511430505279394553645416782912704654223933633933528488718361210088644740752282610530395057328118452602242332084326692320096750881885780679935478768550661490824694675157256264038526184090439629342743322933007160654872453504645632678378920048433643530300330480194513953602493336335460459852899231727836413637281807888645671655316083174109125627867760636070921835502931756198261565850037902028648226219420864575449698772780484173829970872421931255245843829099900448389388471712332721316918450436040903407827956610385535639633756843368111632619788997703756913014909562761034561569484686225663092326416;
G[380]<=2560'd19170232477226286970019011297562083084679009847007189129621457815850685097218619922960723222902942963283897963069250433231430100189796467271778930293767049125312173747561259722059792265674871159864029039048540738011356171594293507294465633638024024618009131252248553119174351788449526192767523779300524973112563816689436177134692959825905502815122805081793295589431329772536032966033538676006355375021017736811759399745925912295306141237500868463300712925559089461360162093883676382134882362957891728347823685459437442023839895012654948707328927644020050823337399776510433037051057790247160840503177442405358569497091703551191946261258149936182400253361911162706472834308648663582773360403592795282296632508432;
G[381]<=2560'd4314294691240418387816531526335713783616456948575505491860244906147635242884235747671870111960302767666933568401845239970966371898260638334310012871953637808313820487400088377205017788145800442189562188475895338666092619843532862013699752367362049861267087542039314118118272832601451902266677613787159015889714839395355089167378971264935317763728115191493742249609925793355180281497020254865172965233529740612175703205048327035639283853646500550810549639880729602308670723987672552569589848212847045944895006382407572869831024195938445120525907070129953954868975205794254799160457869104256303084542802703883389101903455547181673847927182971955272651554153259331252519952335301527092375430471380420423377803542544;
G[382]<=2560'd3214660180265199669999223687560067855603769167660064781131483644717957419763782827263551814254821731197135807725540399068195382383235653391166771609396822856093602345340817810212246296991923113715864363243846633833274566601574219835653711331422368062862513222726252407066072509231118002222919570933860272013554151262511434757249061996313495134210203268079775692976180762157419796454252139955693677859190545764499010793499203270322902477052105313109228011436220423055202884722389739190916475374129161480462925525186553013259810597068242366403505295548164677906784315693055013496806465315757349029352916328947080204655013278437716428761030807463142414109851106191307075927285704838571967053363151351320576;
G[383]<=2560'd4724878830212479338176406827669293450660401657838242488917722710388292020502288625385418137778623826528780637279263124575461386409337301873586176739636873426986653017247055896226576509594343576793177271118457212209978092115729009341085479490644226234657915175257783641309214447386976518615623852545145329700774049154392696121869499345490622531939279129511160381140022893650798354679278180885867857073316570684580391301138892920833332614485629571869016795839754586158390306588513231850482963960785990023567433721703469594853017926801663696102715014329724478672641230707560750568171558809641087722117793032359621802877699376601826643945849903625493292877551920468657721607670128000689925648719017934848;
G[384]<=2560'd67244596584852928864970805954253963277735896813354258169653861598808835605608722804558397020020597024322678630195093516171675580767150088853580992794213405156111218708831810873518411429510154441370643509461588253558920738319510191868626129332416161574319127264405628263355461347257305217188669431221117547056385183006152194346122935635015380386486637182855657644020560564995201864972381850718596184788820378530277527037841891806717616604612404738043193735274637073371400841335171600140529709218236003445231131425650886505216608688227358624241629532271204492371173969837859339549480715301374809593865845546763823398239044208568428631877893057756945799599573322528199394718587285204258949374673030217728;
G[385]<=2560'd279023236836088257776789828493352527866902977639050336686766049498481626183876556489392998284608830524409589784893769205386973676968020401760233989727361742580886776727372078693860214068569071519418200038519542171498220816093421164300830328048660988283425851472862165520616129158257527538911885310514900562682458232956275186752814520305581135419272546596366314091941851782239735887658631751686575860813522594340148773318719035763192029514595594500876818415719444248681030811564285740040289953530137267490089452796595492874302606257220456180643617205632608164188866431493804553428059114627097811316966598823071236001936100926755907137231219934641762080429824672264620488566799246455844441393287135232;
G[386]<=2560'd1089935489575696979225819286325103146118529314825793551003120808861031248781224032683469569913387206222553737481258158397547602000078241511599330852817476012151620280409192027178172612959472145652193241626274434786432073314361281378314464583810377815113966482529985051039687033174732359837840749419439946115933799654479595182036998604993912746826161261662172199594673706439591798250464469426145723836967138549009542441975316989731327944441003256423655781710119098604130498218950956654609150661277642198935796144160579714941511796220685475450487044777367728865708134603557357768802146085078177547454948702421856933396338860010269112249715273157314501582264927459379576484224686994905730485810364416;
G[387]<=2560'd96211974004429108142940779256930945246140557250370221326470107241811593578039555559184917287011937276993403556768837374743637664711225207464981371260317807550165796266567678196554301818020814866190657786627264953896383738388255020070064084664860151998700379602540555373223269604777416606794672657411695910106024818824649717936193715842724205515777677515228505482199470281384821151871681119325608185975858102603356352851578610744008360836139614382255146047972738005364223064196032852807944294990147467812467302056101757199065107353871921224350095720641707059708954914518212869636748166757344874251423051544674689929555871280065560629596499813532986475578906771102266339374140581294116343351910795598848999122750385655522769502878353582235498921178081263616;
G[388]<=2560'd16631095785038944292541898347672254812496280370455955245201706520103338407192103421865674209592451071127605507359053233092082852154635204165849878981380962559594732812643360782989895268702282954796275008535437556174029586046717159685795931205461587323244120757350392830753704914356377498401448502063868662616736675820835526814330981972432903528624792386599094464399899926758824540365085829949551222145880279655193605964722733840068556469305649771075032504330132229122844428426801135556349116339832476516629975905826934362951636375702405758173999323345930904944094092885347005988827470576648631032414871602784397702188614626075079976722161215260784248482750940361657068107326221419833563545600;
G[389]<=2560'd400785353137346596115460704607271546206609682149521948579808627057213119412188085727958431154388211259822261408786770645745726083133916144104295437061404390348168006316328731761546822202778088146008197833362894141141784363899562638439293508081225614323668614463832965046819778262455556293535185823039098975714160642334983405125044471188781605460675859541457051720459034856226661417940901726169854045480748390135347593331544336672303492064318033990701231579784826001555660633555494216194266268874232859654644749735092567566318540991499844493877072758738873993478450497179855831584937286150863654336170361901448542773829895945780561408841213817156678330581816225776995511102819696283864711310495331989602201355200264696645782189776205112349666046541561856;
G[390]<=2560'd6814910836440051220989838121175796600596044167191264580326951941449685698583935097348428491791338055468593440185173067299972164458451551391865153115833797569934111138255577523565785830846080066824830096018271492260201511223237845633115519025473564878889066129922843456174039417601902853721944918667444000689391353387669454784906836317868336758531002504627968860482541297275747554941045442607487238261953097045116393843783147319230716454202921810154387854665182220798620595104863267693941635798791194651993764993947243155821884773161330290104881904111295476071479777067955523358708158327326689354253362571745295948571314528265990751184676202278890311342058013544958939980506484988719213487026929161711658885362162319311868019370562164898588754523661008896;
G[391]<=2560'd12804767449820017847632614557476467791618325434020036711819688469167638325123599566963347271174185297355873968127254398172218615867118710791307371511744660441974318768831627692975146544901295738944411315205926547962429608480506932994783628188603622563763397054500094932881496725443491641465338276351649700623148103852684074627456394606475010820352637068508299873410409650036755934253409606312670882281607182648791832821337552684360996897046518303341635350834554042945408324579329882691628749997748395681218060748902691735052079690598178828700471071205369170041922432135094544307461405409913772835395158145001796252409570504109173760838879486405049971903184358217702943902754528945550731953381528802806557919672596744791246891246594723609281939571027738624;
G[392]<=2560'd109016649699360587220748275806004343607459842709646176188026838200528108551258290603349913465301215685443334753417691083138980797350642024284081232100223858111329124426260085796009637493434956809916478724377389055290096660069014867006814716025307405458441733696938257990945249257318153913093669115616226997464330614295094654728336765438091094276047952985611582096748424040540851142468405363980001739134123477671759832550894209703936136511459154896834578319497699427711964188871344695912008152335559032320999120002765610784544471933967602222830588345284127612282486286924590172963688756617287913367501549309581336489604996503499148666130714716393149488214308487970697550480834982855332067475448919240921949824446450626906367869851184707787149951234260074496;
G[393]<=2560'd6815008326009123663929026005104057870288774140356851546231339772638052323473700564093741694483064345570081619497127089564232539616992787799453659673971018211697959514940243625284190032114510904985443270559061299493046905808594763289590000211432703045550604658049374427622781224584066353874486085672565064622437117527045056454236552364044721742586055344974122508251809146765631204467711064112154143298830726717747425616679949478818853833453621554827670421412156581188734785808783052560356558930025200660126873421363327013942106494159585029976458483277037444381245488874078579883909626616123569647834133482405803314161769973039704296525615189170275561380315417253882123229322501727387275135397301608791722444702226564304245778279629404912595871540952694784;
G[394]<=2560'd400877108025885365940578713010340976505649656893603798842761878908342338019575149885012886291445349865050995366855335628581295944219534200990504067696650973987363725621564837948302857402506152904432162759772358530524469458203534511931919725777223177397333545278819900209940665353679471747872146779288323323683074523445447687900029694783438919550520777099126665943181430931755803850494391928470231794595621769947668899900468052378165514874522542377197635551996668104389874093066769038677353820647645706483807144463210763478178981749616621108356253625002062910523990106994283044185052221368868738393096312483543761766533234970036520870666824460174614124481129628652321477849174828256239683257763178233428957866345552724957341204926044266780170103317069824;
G[395]<=2560'd58856462181295883324680253694024899352254989735633295466412893232666729575246432109908426866953915920006242715329874419159619316501882758222238966112789344691612649366724289343290628790475895636744992642242701850323700801548124726968725288713392535543378423498590724205833865094280262526410513637910273973215418716279572765493206685811504732375759112454835633528574520214686661293799633298186263515146326692899419027647964828246570178878778024274628712833575187006738701476986781812537881185863354994210893744190074649778680931204396556763453757164350927962581260420562083419359353701345691889123517180153027175683625697740676685457679099115028373804616157595333846833538531328;
G[396]<=2560'd3691999855047665944681715133632937924044506934294680815005636931981691470830799321858431751119487450525758397123407679253587090572888832626994011655019311029170691296201900986664314912049440192123151032718294501551039070020946098271723838599283909252340795679836384029272916648843502144512354383441393683105591504579597921968366237739537679874986201798109096626421859551311240680634669679339093757289248053609790663960924050372231619330640369532306563311807094664308633130157572444409471551548860681556723566006713073067474837583063056301195945678795083875405795440831934127774037382958585234012882733688722263722708490298590314475597446266960028174854742612458747195461468160;
G[397]<=2560'd1493041787808189526630419137355951764459199019333429443015935368902126370371429788383988891427451548324366382609437907753494348981960929530884290821062713729951648007588764577745777642453336035304868597309243034515779773580781037568904313532153816616868253314399116628674584251535223969897505558311056474776620954413639749303175458656997975893806453781042843561294427646296584337384264914498698880782464541447176651521326205036151561144211362293502062755355255740017094585431055946479500133049622114663338174287501079153685427639985307221518125203999306368109118319670973906554296496843139547729537208472057063402015036398306294685100852847429825992750989417351399625359232811253574608940020459958855511545839410828845230470099402976629876588544;
G[398]<=2560'd1493041787808189526630419137355951764459199019333429443015935368902126342531814733941902575051930703646383066300677952518675081117793504780131392184545663830876813420128951727318137704324816840792592301199136641088995574495877269034716991629847722746904478434400765344597978110390315371595188529200975601064636072304680733160466512449062311405592395463902280376107766080034526629301246617283280668531211879081814740565517357215372565854320413335957061095623575794724360464243691348578124944289104154589587378426728125998633421902439144837364280869909553594001605476408749392777519234059519282010161107817695381295299186855116594704542912596951284454852067035320097296489890029984834693234808846446907781425770010309781226230676507239317608857600;
G[399]<=2560'd54454047507783025985249257063142195026691018582892565365786824158889650302959761759180363897621591251521948313274797990982449833407559604944349502940533962502369381299584724940286923419699354573883902990082949092930373116668398679784286224603364494572808273102925559774446201664460932798471053177296722959937326546835006846142180113078723117580550484776456772984374565852226534275969927481597958507261035366400867483221513716300738071682019437557000852965392601759132564400032056601877665150605198023891388146313493871049601755693239494292032265553492358919227968916707778411979902724969874877439872794146036234366515687784151811999045463530238407890855010649642891380547718020595712;
G[400]<=2560'd862759462764354276519207056356300960877884527116956796681339931056244773812638906081158618238895711728754083025286869784223435238051872433757054367596226583910150172085478720961770777476546273004505274965110792530709132559177565798084652881885408727913952033726062130865007654523909190221862688163458165641653436175460413905884290996583855711484660942173246588170448639010104180380327473852227021022371360199982029955222482213284335725933315261720374695790537414486304554455181683321022240992780602861268465419576655232688360711332939646276208178139051039679091422478449240058712760342083005167974523575465042020534370465181069656249995538013338768968148611659464704;
G[401]<=2560'd3554603770600170577398359313318491409345385255235375741860417243772272293790017744001645857931504379755006249473795577932539824954125306864330577890584368758013338038103101307081301716644586797485538766697546972443503536536137442561165855962935021005825369586167900610089013654343449143578997308316193786291331520752214936145767257143914879492738237767147654725580662801459241004136967250142564283481954904199385253621941068873955167965846032095639596646604299903238602838230579435554750558952442598537993623555121373961368424157027098152222868771504350440084005714647430168032939239148434149968588935997903345156447902008861953902054899200050933047814854967033856;
G[402]<=2560'd418146076142072806661647774440807452123948664284203288376519325514438189521582194352561449872868147790510761850621086506514110953763144797909904410645465302637412253107126641004103563274583878757802906650286099634225199672177919735025738165016054704430320896976079302505577157913026787186447163376211696355710903684997410817051110715308774091792722237752038368168336385506908947492695925276008464668328347564586184391925591471218445367297540584168425782296596016235510123578500991687048806855465198068833010460803823120160912525497228753316709328923556215289308324847794652060033684992981342732087460220741464254883594111350926207417992436079324007970699059658752;
G[403]<=2560'd13167479080817040158317739695105513500491895454542910997115979167292820195696920533616404251527491186426867177057225608403896608408248335354189062585813760941864709954626455990421363898301080045936019279706926196438282720170442923430142066628426366117391058293643525272745907854552798688703559870996250962326282863367467349547019141435933923810466928847030635403477983800514532592126032773014143377446660938007701305957908067344789094647492596470531022819466292975252994266221191694917670713116701840927325428329188921832988139788585887919787327559887151837252732079061254242576924783545849552357118314266722738814521829216638251950139142628505327216154625703936;
G[404]<=2560'd54251363602570181252200402101072270441645334662295711558434758147152296310700554327701543364834569766098235576887765112169166040621638264975974061154755187852906479232691329069871259118329358968588012093477697607352580753687482965276787784609067773615828259155567849206328362240231894051474670416773187840127052588991850975537476790699876625135278241200058622220597154919984777668143596954653712817856030630412862663280675642358101247497615164003951595970614249860271029973054643758196022300814254294649955695821501923274052003173483719967864746525346632723313039739211068688363711080647401716396689578219212743721400504600968414935174040097922110823329693696;
G[405]<=2560'd189882796098496690197432474845988369511029879101457572603431027004697948127467961557584046909360805703173437855544355826340532356797590507037232018858089539284745944792754241009232201923771014060530542223297418704772419623788887836408891002658558443507939492804153390874411832542176092414541432788798916070257166706398876065050075288541756928526075484790737872986221161995336548765344731461844559487657345652075581910203262672938715641001682246404219195692160199889298266115712397784815571618415877579655267679454352382155204635513879458827250566235503350433231408173864520639313404368842643930713475734156574902521912486776468869593530462909366495808061440;
G[406]<=2560'd781990368303030078359196724291483127667839304523906606318060677197288051842131535858223309185891565727243167235301103585242432915470394644862287069768393393754050428841534322238709688627611574996004619901301424771970092809178034732651013120562666787837981830455805048923731314762511584336029503409648873695810950445741019810722259275458675472954591511817336384017776939941472295682373320793478566849075722067721347834564846175947240416979298658382096520531076192693280573289552646063322103863193605597519619572254355128591350970489370227587104596845271761004112849762525837451930429835203834816258600977425930138832616937270622897536998763392645449383936;
G[407]<=2560'd48695455434986421465480414896175926863966434814920069790906724106928764660453846758748047903419062512135842423890629862722953816598388441996964272841832181624027960525907523456732487124402244843662386951715642673602166087426309100793895899555301531191279476625746212598052620685588571755395315278063990627051923579093045254147935218868477805306295802705190052630269375857315280550138378296850387721940646653657329796615603564621544206500802876089207513742320494498435738351901734321478984785181980121111971057252686250314762608290851945380342821995266465558312797841309071406472382783435258521212958350367311906272627316774382383030278985393919701811200;
G[408]<=2560'd190216292072548167607381701222653857877838928407102084057400236602703050388264941318822268263946740728901040722991104747049284811289893915447741657911912008086623208344470697903757101960561604210081877074834478740048191368341736356459665209752166197425784936806567620291282949772199094594630865540197405570235464249364803686001173607994797500567228726588154909404357200860054197519109674090197004210286864417906231594691430872478844328934140422158781547375937788315612212622116046236995703996286724641891926355125371085838718392478599563602831243032822672849955733331170436674489525979730378063961719122712876206206743612326930400508385446560014532608;
G[409]<=2560'd11230671110092207112322984547890939793483457866417335729882341523960568370673023966672873401997583746144008755164710562176236691139031401217916345998066361985050273038758411432005134175803783219653104449129375635893636981383007882969823911616836858429596598133265508112683078490569929939395436413793687974569253173003544919253353204206831757835167597267509267879565251332862125347948162722000508221423877634746311509171755932178267589341181847887960892297185827363604475616487012344207716075234104317613668493681193784358357875368903963650525904459434942616093867550820344432265514910465385356033198638971613709827226755696171135023447022204142747648;
G[410]<=2560'd353388121884157953162486170473692293843033106755676087273748106100233176799896360171866443962667266649679229861116259373601823547751684027736982723402304124324463863361671570226908713187134891644810607105990961294095218004832258797896030277578022766244141141685474971777941317326689544093424256758239223702970758890695795463110715546109224744993439659338233886456932841831833947590863304608903664035507498009443064962643878294902320518075867887969790005263177146959025950057168079088373000975069584286990868449028923274966111899194279928871799238025105364677463671931798508877035303384730962799179687079971267923061467671772170270192870820413440;
G[411]<=2560'd12085291463313101001923473518510508160510972280974237465931984750726764640495820801284879731979505373106210966209950008546549388061482761699909171283672152325614946937928951453307492573075289882467878103586186197382086946656183351648086785728419204462667798192712174746231126216073728477396308873709988215769653376332383777899271268250628039171022558894023655996249296141776896310621564442559746961192877545135360295359292809820868952656840674279630347926724736001710896045408190778359866726286969516131036226219415995542447102876460560352492519743527064381022344442783422346549929752441743529590584363042520215412138120158350234422631645315072;
G[412]<=2560'd47208169778604693865393437337901749143273079816927695950337891238931559863250938195181259520033206864714389471265285147242173263354709938910992276741853661147855324523948741114372819376372615876333304947125181563220151496855116573475046526268372687891745512710046026527847014299448747998598980917746634162378794762676636951900553810831603973890689117073947694861316484714413893885617621058257717931618976470226251229940604731105991877826391935898824271117964516286724222741115546524086971352809455356101104851359824997962339144314801207963760224373563824007846329080463362242364771171450072239746600721806188296094167973724704268431600386048;
G[413]<=2560'd183771172335377129023147843921592167878081122243790383649157178779758889576525030163045210922833035117036545910704782586375500740748153426846314657728032983590027498156398500995553018189025833812918389334086229955804617671713580447461107232352159204069729046159436277889237833755713137507432582276284028315175737425927781574397791603279187046398264065409609046083565613760781100579052842988901216897391691310413992982695692571287698271953232968925395593081517426444066843220040703108810514365065334748681006881825336261008760093341186029848052371947739775169219664693826935945948437908547964926540735293440320573401449995642922194924732416;
G[414]<=2560'd1311661331353718854917495765775617134761517580504000237568875479528161307181331061450898385029366481654917465199763421378467039217025845351698951592677747494038609576224764487869636664738053762323358587545728568196800942939945741357456377270048532963172400053917309953352123835568396556416500946388703403053158877778295441658265225050757742588707603068867848602825282519774463461354922055006917176020113559478500457281753135271403055221971828704026423743495599935211263805821146487249084178270959264540297678030135182316354427994764685826791562494575212054123547022609896600639513071872240928059036697154433021323469176007035090481709056;
G[415]<=2560'd44866008861688316278356006068964728526741371832743000349787040378394248413834583187340626873136985032338087073322660614162118095190565000515771061614600607616321129769784285921326420438255548465837401734250701135840311271226586223015864143481801959281683945359794265584261220780881002365791727634060224624047985868291256705646837672948350827888091138528823802147617226143387625980052405061446460506100072299846378643137502101797451314184008228472774286240093956148764741179316273150562650616003959354519691529993950856722732288914217053619081726368111728800567043450967359701500412632153087662146006997171995540404382885503667292602368;
G[416]<=2560'd175864136882119903527224338504328807497403652721420205343223799490133997304233735919937300633600833428450955353744314569238319116277561670618268334410407015833083941438580630603295365328137207150476726551764483421095101364930967437945297732446531697029381589984910527966753537652146128460354521189071554493384282344381615183873611722550090664059239150563484330184241310734765908066733073920906600632932012176790541750003444668721011933240594536272855885412294473954365124395260740612835552555598908171691070572259210219524970775129511503222032107807962282355045806739440626102438121115859013585325465820375276145314060011182151958528;
G[417]<=2560'd649207456311934671352940814733672112750689567363545427473052128078848310326531611439229755716718070969601770261567649164372808129866326744684818560374514336635060378283783216639930738791994757776352547416055095177632690187532515156509592828612206923391341454387369540309248217582218149434033538571105112231272007193235902768778186347745635043028411983678496469406945613538902169476052897674967606351786028708441638658211145258864353209377090830111363863572486678579510847471637792343171658766287166049053401335463870707181473229363323050639233065009901808263607854542898179794061966201431597080384154360893259947266715412600979456;
G[418]<=2560'd2665581518493582600192521270334081101956713046680200175430111130889646243387518478478246034714540987527472272924042021416848175724195531196038795053395469885241797271509301566295030820224070756221328215937900525240994170653471551244069288720996151004766783098371532577722260462878360038742403456871550955564435288417934449186531065171261004783051917347886871930115368256638997141674308769357807895302620342746609470243880686074374137765714450855650660287182268616045160897484899014527865654010062716134340385057005640371513656699157328376683883652901261581523810586246529042702940693645861941789935511041230101142506625394802688;
G[419]<=2560'd9867838649083348961383117947360202536396008939205073965512728078310014870626085008376041989371641204876961233619957611347703981695399055791974777979382030470954822040974702296514374605789757326223717667637663449800688740919930345726594974795556558094366923045837557848940501070310892767900789840137685410160156631878229284748968434773367657670104493024526172123652579168094815531027933872719908578544621827036576398362503207623551122586254076690791998775555062029399354816692299324018369660841638553221265771459859030077633227863369086944119742110681444756206893873719442172183133846885492408634622395648626722818804739473408;
G[420]<=2560'd614621988257817817252073664607650570613140151124293041016620088143030603238392144095700279357285809717791890027775161125653816895791098494220034456077935061116181084330367066340934392087843257999570059396866554916227568671755835573183713964621768002199281068882057705408792230349463664375440469383040541386898650777206516977096670993833752927490137273026186355028869841005132956393485393173299982775514073590820654563766208381116399549245655446059162954976452019357402075829575658544561454535790073770944335004232012114259083657353810030906189099940089792768604647694082171598613700113769008329924171476296811982604078153728;
G[421]<=2560'd2417999329097099916215676087533862648944462021751167645542637104046497836941438133340362126406733728339249133691338694733596367999266259274741288846763407062258435697598738440603767340581688687271498862974690878032767535932725257636021892161030538093939384004169464620957105193311895440532742772722208826852458989475618587303477115647210651108350232799334596954201902683272622118822342195514431527398615759034440761304419137546445379973664580914251313866701076613922592584560837862625376437039869767674242416677764351615172135844235400490082731256295860781604173986057243434159268335671269798398428815615968391953159028736;
G[422]<=2560'd18235417675525524868871209281670982779006540399354570754025529795868144852742933602160642756631306787029371175704850299852179067074623843443353606822927029039164764131457576991336930867184636567017876748676173329121352757341629629934568923965448059989496293245006699027986500949605335212953260589801775454256283447254640172027437690063017541458095822780852758151073096918403866664517179410429693689123870443251504056936719552399604698170452828491037437082437235265215575185823326838704087222103940067271849223280235443036995650775279407822983365507612514853305084136546393258018679612617881128510275380847411110896205824;
G[423]<=2560'd38923444618390563941556505296694389560578653808393771560941068577334132681075200208915958090407251226775013832213138599031286959407265190077714142760843682863622244215497469491914972094139573731607050396133733741563294588495465211729424245641532628639571863455121117045091959947135404290025395604813230579020803139795631902069910361966250000858615530781872895832774185852599265282478080073471338958642490597667890037958682452680867223013751049072216531105573777822627724928677135045164560659548246522645135930753035170102605263715361638494861604766954630765398608865513147818065523542828866023877034597466796653019136;
G[424]<=2560'd144122057343212079671132011789414135931280991204454263090950091070164564657255483536170107808426531268903469411165860395565681072621808298413301611466047698927223267350492790692421706942764594034849273683906725717869183897938773685836521640861627511203205192410989499359428559786344372057409920293592718680938653350638789875675494665908132518125661471277725011864698162006529182662246037167371705058974689269415222812784200041320252205710586436227671255632422764974334829927919195098404561606392146402223922113612593547820241041825882096090939213896954647585646935627156909811137303774999376313655315087683724771328;
G[425]<=2560'd8450823270356355490187389786611762758450588210052241976825111696492936573245091711890433497840335510560843939682415120607245132038268750384218851663976491491924138607028759401176135239482660065257885658868360242526045147657782990270396370273850112934841483869930152565507272987511399111482020911183450486738407547103472385544362266825617082343952303321492774305959028442787370638893516230660740018549766884099406683330995968448905637553816010011322403131310986666324240327031715832654822196524193920483291385958572071949458808568442498692134094979258930920863337803590297889360129142902395304612316845514625646592;
G[426]<=2560'd2191100219964868343251200982822876921781413438177563934861127948492337007413222619309883803106172037745626381798764340440249651599885233260889092911340793342237652056894497621236095827740042403390128307183398678156723379034155054191505406613694711739257547639712070058926684114029254654385704369412834662343522109788614992816744301394178616164640458641258312932160372411843987147995705380737414079502805493255251954291598154862859113256510583240906471088126228291983573985081682841726325280790936563681379098616281778153543494873226680854545994538785035002274386332849095011025569731836500480726871678864326656;
G[427]<=2560'd136975237328983873300432165710633630479984703493298739902506942820231052713503490548364135586207913138359005798652344248314307643931749912000002178478296954895781898183432667612235486515067118942277646223213258662605111082258110741041916488481761326700495739058363109826448939679830316378195450612959474610453631816079852722631299811915899510839855401088692683200988867635003237792185611519804374604369116114680228916097409952748275656857424618434929589150111896197521994779766060728765942983304863801592795429302996128834507464857216870720770185028378842339469930401690786578807605047619470338688084839759872;
G[428]<=2560'd566411114964159908047287359688443423391573498858615818056383364505829263757837967020307449623213418203262481513430531647780764250369687203663271195455594628978621616085587381477388458467450607020828859546339109503666956431796573964893651483782520130218515272497266204389537773023521637791279066495949429330219806664433968279060581713214107898874434909234155398451371396751301549606867514934957195083652307479100037227397392443540404787034058772033749737080552465888995144048507475980409448175136262924100343380046469879100200510784675977354524693444913966032590991674458842238938711795743384149206914564096;
G[429]<=2560'd2097253821942714468063510913820096631963095166941195717018050536356780203664817510245363507143976140654040353499192640887328079816875354406330418753363298376920539825242623014667538658933024083280403649918650597566809866274684143948499866950775597384029462407389340929865875539437500713144941452173866663253931670699720403857715077757097524789774225530404189305893794940811427796776354537025298899713961765724076677540575187510541862737458805721641608972963173696428292687283585973181656106273425505686927108449262273025311582219768557862085469805953877323221822745610188899013041528761219505517498466304;
G[430]<=2560'd7687724482730840618268383820127267030730070676450039415483200355659700170200549796341013970552618344549864215537379960261350760421840978023404216512062325789976672079802829121464851241684266300417633880926809433201750266176610370928792521750021667817475932561202390123194454365540710304910453948777943312576187654778203924472932153877354937792232408307629314952586061713353311875516936398906207171960103546016411214668421348164975268347151472117777455054721711256189783807954322735441644266343328216811984531356596831116948378574724429300572656762089610196606640441872833965446993306707743875612540928;
G[431]<=2560'd31884733053575794003346729589434869157750505597436664408364970179656241472878201303875259579970962397245180824548260505993285962657067273346464002261751096995626308156241718086019311569555928426921649168156274054537882232211323778370698956561648028648976766466219302015686981752264254384096780647754625585228765459969801369389052626201638737401399818926383362129163871891207825957337686907763784986151700685333296241038721235192664843997540106682916024800875373296235393067765006597086113997168357799579158180469807771352277201520909353927374322700410706260676176638202250099080328935620458791829504;
G[432]<=2560'd131877759614534645267330563836845296388429128579824446920848084090195112161362379010441205437109621906573958512030439860143039708037802408692360803534070185383486440970057646046656608643135867034047085245996525648402304532936316353096396280166812548028797853192307236928461783330233620262788743924775923676220736133281863631489428184837576793176521352118664863915243714875684068405300471750931161544309169325180953705194177197321385844205986461804659005536819070308923777232228883006655450452857183260991787603082045761995140305689247807385025021487141819483052062564099334924215563548191287672832;
G[433]<=2560'd7786147748809003077865386273987468093383596827728083700393910443325307034952244738668825234942860792801484186206154572175083519848122068072796837602444291474667965113428266101789678790476922132619923401027073335640137358346069912724420633462352078215022614221944580486567222758325522964108430077117326039365765652174531209281940380448398498818885311042701762787032612067015811407685101850725298318525941650902080548629707173764918436412670955528260017821010630978973860521119728416009112897055413226131611401903823759604166502826454716473565228634331140419050687447627766971773835137718071328768;
G[434]<=2560'd30414639544226536895309685029687086649362395516116202492744441808548221364087790451212783193374492241457135205176743358780434757224913606965069503945896283878619106932566888263162350632351302713331304163403122883631924516438050528129281911174997946297946282774742923941529399096076554306780714971010173468469806599546328897687815438314599278351351689440943938785009518753646254416508043554861252209555000282631883912248874083638180694906114006680537268812121905933415845777979749736109542328389455105939271035711661662362812579139857105869954840785202447476279582038157594146706066726096732160;
G[435]<=2560'd6990457168743211582723418222802367476729289544626533691963745739293933809366777811000862428187889141585579068582525624263913883411090436937357725963446149688554104890035764801219359771251935478881853017435189419968868153827366682523613712384847502615656903913314499978456863194490315896664122329143944598153226775754754117822476412219817531581963609028009723942315901305706330547429407514143618096843390559138939504432497518320650063876379046261832273253883610292082750263323667025283519260592572539930769089131116030740892707428252663571315830018184526141164590009432546950823300084793344;
G[436]<=2560'd28998995779671344259817188915661462555296675395702768223921343744674997946318425798789088452145050893849797612965432584695557673507444627203556173679621248989237652480720907714424751530311499456214880982776939460429529136664137590515322892256972874701877951502993328040631281211245379192955978526529498664287676178928159675051973264957631204952022680187419879134190944026698832525941469050774030682635689972190371062635634065298818203464210839456948652304449896346860375724780391557415155330651433093126301244031408205772044091937881463021276917127442583575255772857289003050566665895936;
G[437]<=2560'd107053298293772992817906806111933465632776443445406876148284359593019665757219865135353440137897821024905970720670873665986056686039305324692686538617563329428302521918565318604587999491034083920414689888884106800948729422980985241864957862950473332495578249989047612390432814590522053724913229864928881481453055265163165586851415312815782089219777919840124385596301878025755674858590400839644313716523379093336802988253913436418035856347763464508028500644535431373925287046617657475601557957426940456008536993440046790585932642158207329774100500150311071000246704682145503224359026688;
G[438]<=2560'd442590837449500599981519648314114960093641655172812231205515249378587410071819495021649560172961773669383124277168487870973619621108437753158165560601778665873638052087551115812889825330306338494267331309469866346216495490921579382482391120546010424497635130073228457893540655284468019290664830166198775091750275839184607047034702270940193111652594167009582276967365041159765683925748097904594114536495411385565064470586849584792706513724061490390555105485921813187137044944453031958451238239531438245606450699070233505692854657749446756798766023051268257793584640543739922050187264;
G[439]<=2560'd1836084074759532569995027877138551484048119585985326447504654387268221438123886574512173297056122404125318094939812144622209495883810442427168664038679916931805049959924655700821838609628816993218713451346688342305042997150621059694749573782924999690704317794823099474381561060770727664477945101904027270860972731151805067591763812854992811765037938987842574768232630171276220528274170885949271154430777108563405169724628635070335374890255137581680229139506755479148182945454109705622121622851875318133295927925644584379106939026320830438248450893464291373537225503703854215069696;
G[440]<=2560'd7172203393448820939714182774628451379751224834360858683373250956031558924054958818272259236568806488263302590605085281825522145015913216418399755097815138150142589086005505407414382582472009339184154197277452973894425157494388798774208484502057360359724446838138548033026191095906795503059560510707575754873337166153925889684798095042877475943627793736976068439276366019562255256792018504716825565214621666588817927643422277807522305966911063021537454280231213442554164360251864334137657122507612734570179388574520503482977307241639640578032946741658729458330913045652246102016;
G[441]<=2560'd51112161323069988331627226215827222810092816928409239874812411820556793134322393338217069962708418068657126014948622209920291392850366686974182010772284083326429067165277774785246345211735949470694488659743275161792119008741628719344904446973369798882619079809478050189881988373809286836202171472887518966079830718065197878244957992205926754554045229963155072755242164666539938934259894730628535421139887480026272546023914655791437124339336305451694527289413181989727887507159184559112033946521268625581521018456962314377397122657042421521451303424802110104195268574797889536;
G[442]<=2560'd199633299587486091274277558195628147385305259888871243916227504553796778955266918398844160221078340375231776234956421507132802424964600864660159912504969312107286085051618968420687910863735015452642798986872884446822380282160066933100700878308086864392159845065230765925083289740913649309374780144357627866023971570388018052346072741615107574723463931156893761739500533868703738759793468404305305414078951972598720113410428188182576094314795078805195094645953670283756623740343738269935183724149455077801024222498050107043194023630946165815493720092239660676042575518367744;
G[443]<=2560'd6415478822172442691385804424849829335275437240168293701322752372327057503900417050541343527396990503974898670459630212729872494857954362082170004982706656956925551863303332218140471525641811572039046133428461077716281897052893588788910488599100686326334033089646441060576004990791483220376234374952984583936456020945299910036920197815516684587181656437746787386748154614657246160569700781094623916946066197409184175421777597671565318194670604008893000879547727061061018767085370404826212436957275054165162414118517315735899995903152310092126615478089476431857256081915904;
G[444]<=2560'd2570999922049101427810624589757922076799569653180204733358992781382799042034878782027424319379434527126711106117171551149820849231125946237017585233768738121193778266252791000378300860257087733325107410648821340658465957308440578972576395571558985679268447875274704790428178310495268345107590139168180888173049096317510385420846296267438099001960767371512879860882064859191481110556132511437870695747251107643372459792575875225539347946592620706415395067012317184;
G[445]<=2560'd2527395763998834195447003244848063853665333801896035250464504235008559628584988606457057043391706961051340913841968946793436386768992044479871328251927540430740023020954896510537439070230054936694674253566460684334529257272752629298340383757652410215916376914369291364528372575686706853451733273427170629313580664947569149949057500735577193153869988367960643908268970077847978355625059246754232781167879206258337534506890650408101732429948292547848462450458540097142784;
G[446]<=2560'd5935696575181333391653631137056414439340741311899988945558394590919319454037270122115077384345331547087937985971750382275458050433999320639461061995483760085053624170250762512835773288766513860058263689479693350236960683056570341106030359493653640516922874551547384147996969433004038158275433630198222485042248453056150621693368885138432122296719127741495475828027115937389169777630326600152391562438904949042308021339316657660068371138285340444453768298345004159439708249590090494462880662379424904804118743910236800168956110624698868447268260081285967184146634570366344757248;
G[447]<=2560'd200240922278232540849726515757695833016074064105555419586077630674078073359514318033384219625193150122168030950282630606867592104255085393491958604773718474647094352648363794903855664756699434714116340871226436957160526197013399364211831905507210508045409892893312341364304533647716195218987750301165238567759659285078087764542160703426747556715326353842951206742901561002656841753161672699767536430899852188456551060356317269313846188062966881735718128607110160587767231994332562427104851927236608;
G[448]<=2560'd57869626538409204305571641484234199088989820139015679862063956769528497758669359196777502821589668255915338558485664205284960825507918104779834777395979336882189483220789055366193760084537380160827283436113619141580434508905523918099390610989767888997726736869313699447215558021063504025006291708015275842406498319699183010893433815568650257945683315860947993284073273729181650485169854497506233756559308889899891682511465448535207213464531667866873490879423646759183196690874184808946024613549178880;
G[449]<=2560'd223914405314576582991685433713546748905705260902739850180423393596558108399678035280180151434251953352637256804907088753327965315701802562957564530937863613210785647445426615686825083683696089505693545348768098112684166478810457971752033251679791570724168813627946858772294075761779951183656524424816787600519774971155957426090222917539845107470944389707144340089491738199125403852274498777952192244344631076395361307091049422656443739754085934657071182213725428355146331617016768522127235067426707079168;
G[450]<=2560'd237091872442920152429458039367608939986687657315386814375555048119499810060053352816308669224658846729804611918523629128171985401248856992335427189479149862153785207013764160488007349662411632428862366921316759666813598808021257355094193753263419490456857542851165644895394878959699292309174130902434752159011097160599792861370321499026572315743822508282463255341714283397009530922355067588215665133886324359594554947456650506667705969021228502002203847444631195571579513040549243807053870744542115790848;
G[451]<=2560'd4061368405060091411110227704044861789545090709218669599457586256254496920543129079902935394722253174313662485817655351574376771494226819161780984003331040582606465770872482159202435105657528364394183256761475144899660695053983219273489416327456784412833395038033819403372676704943418162402731166079824586680801709760109775061090898437123544459177644442376735766817438084880986221902989525428921662530986994536930294787193979550284711062865650648379864727176270146942242454703368331634959967105830679852292272204773127161145982976;
G[452]<=2560'd259156520131924496662368514636484344437290429814358704783398243833470161404677611549870512400749935984893921870008731899233925107730229626619864164916558618240972555685894416191854863021240697142237734243612834100452977030662461561160365460934370587370356304889602995806363924253383408227217278086387469422872614931262942040095770856357080739739822755978587261666018170079733931707699720227649913660438614262257692560446445491239210658059281312737582945311255789712301657946798159612682841442833810141314259171032214536192;
G[453]<=2560'd16926499725022794571975914886494747371974439387784807282019307431864964265911406749959556206799291061544230678625365062275571946026228528077091783261259112728384329990120349447526568103320181103556427601764802547082188117005492716176536678741618413383994214305115317610161338308140666537967583163299692468339032057094173314934075270379801913669294789360184303112223178585359050403033298565286165638276395224353939115878696832777301431690617494148786588580196301593645181759300667686730419259288842327582632898273895915724996608;
G[454]<=2560'd541515772144588423057452285801975925394797829064712875734575371062907906953358582554950369547356621068875153666306127853440855746986163865803281295829285347244030475702826137995850150326848233779112182992229647865043260417259239433585243588158167772302086877932494040437064270363320796579997138102633256692453788297917605428525126072174390292369955951125134810807734305401662221563039980945570482655633571932241499172140654308630043134364436206382570035368206557380056516478054961172138212637506546614935380919414034502319603712;
G[455]<=2560'd540458140260865429959244538885814854235108406854623886198861409190371681419884888546841942724325271033769763807297470112266964463367966280433310021803130388472860584415983305952439892110044788453940946906620985779191448836095172447328841900139599851030898357926408808999548188922796351290978112355019360798677579149329902902092821617895755315230124356047771913203080084360373777181176112441917882031537708788344314192837488697177614290615770192077985858443284813521473718556765881654774585923686240871229499064154188994544926720;
G[456]<=2560'd5148396096422391593693210985223229948801183492992608227369323946046571732449655968919144750263120290927731619490550057069169514345803180878355113508912121465536504128346048803546586007534195996790240386907138137368026304828291887990441335709457591138003493714347746164547597820851404101231841895168911536784805676027879155219118696168869726296715744483106540587250810835727427548367510321337165796419762013236770748476360308301649175923332805375842025558938124132006931860904076809850148118702653006059094398521235458194321649061180156519882184062741023555584;
G[457]<=2560'd540457881104345298034751683004320939014265623911169199561708504745570910673736170903213925449792339825345750192013605983694165758530947280051327086405010051492853838417370444458607632787479473060218366957146366110660774592202057061763041465001401252364915258442078583278461471470494134514084600505158316962565080295730328706587946630768500645882606181468046687315183785766074886203139043314224987808084068969458297234494087729837585691627385264981240582397539881024729763879412402177771913174171108858789282464123835819663294464;
G[458]<=2560'd2250297766757528060363378293585466094909643757097628584125300212809396786629648978675107528687434264065805909716933873409112118247433758775930778076439384675731689337155471411861268032995121690307207800787092740597213301550786429856410416017749721412417848999335223950243971096448926576861247855530555578028716380307447389791331162274252808261912941749327504601494086120642560843053794888031697834777840660844978720039517007171928392204101521100026042446374465452998548131278070570996302668278579761812953604852192976971862815836650860506189662786861020749100394644879867266621229343257607630926246192445393300775292108800;
G[459]<=2560'd38255062034877977026177430990952923613463943870659685930130103617759745372704032637476827987681779675160737753933531249188867250244690365388104509712140232899480083835658999352571950696720260952409822501085365349827937117804683546192254384938800250771891269892497179022220514668245613993539373870265921013852573923170907750019121586404323920591055504721712651864328251702819993793149885566851796554588648918015643367246477721539934481530975179833165695953219959152462084162995328177145745075330507698483385044226024248983221274726457028958479685408077236747864240638236189182396483506750354101208191308116604791535542730752;
G[460]<=2560'd578194155599816621627484493316547994268548466529555391497606548797487059581520526075940878236620957890209353950297575690556175103117663551561542462052201473254458502115128946391261744042331387817731135145890941409345007598547426028425781867928544415091719386100021629981932435004259071435931439494790781193305616426386684126472251490062128554383486111425018437859611377744598792386415548124326044221717593243747513750025064469894055034739725294218157593084968185397291502318249261883934395706874407678524046988114311979098929017852420577077718466482090584482629755137352603189377113791443629043662904000508604536526664105984;
G[461]<=2560'd17892249913945973697835124540432957712749807491727780027002857620436413905766558647575242727400475129058422710362796159695297865768634597641993173189005032022900344170620083372229932931555900900233805991461453681046629609408665910581346646227001245778169129650961853874742667970141775720422309770669189073661110631662033577056060011900630219334749983728273865692961263206599990422799831371834841450793640376514150784295731819907930256460373216385771822210950292743875662492176289181869548816135839621224294683813744831331352454831735625921276864671776085794556530825349708312683769634499174257890949975652434684912110386806784;
G[462]<=2560'd156692734094860193899222757338943175120748314094222073569812904440837945955972595370509221404245306525125748473206089943471967458935088533955787882061084148611031427744110168865128689161021328336649808362295261341481725767962178651629486466824739306633219152542046466207329410193653492170953509097402419084584210525608428976247926379427615214535186680970620426607785328433281200597400076808352703200735908561407380080130278771413845946567565301317081733474864794164371359952173548939444108917494159155918612016938820113051228941719765085071377178731999907040607467775870958846684455204464841587129296566820763831045568179732480;
G[463]<=2560'd9096567331764575249338341290715964118267998127207668515915142038468677705151668321797258846832086143402953483332016347708320295818309582269502170152122135215730839937575887007167754573580630387418156459133592515261019079499891659115918560837064983413153343548161955237997413851141898324311108587744271240287263109761824146892724952305591134553648408178621174706014987682113866069432547209848300997373442168830231134757952619282305731709241808433702302441005320463342821568831843217460932913872605013663433926023167613815694263600809543229800137869492395570829921238272843666995596398650945328534252860937430188303834905246222516224;
G[464]<=2560'd26169656929204717414879891957885217106950231572101753495264102900232206525635509345928124578774994910368010802724137634578476214282485102568948680360294486441102000474363655577959478890710134971395886786586525915476696523018611854066384990726898682894982011350490140953015173564970752801234095414972916446094718266466234087062132240349471780180642896179669271078426413734504248898450995291224479643576963079822567015236304476860478919588896914823346991060471579309742240161411359100982557654503039978701150557468459158364362405522770909527545844991985620072140319633216091542420813835983855331969024473535922498222559449501878089216469838201551521313449716768348322362480080281849676422040138703872775489880679263936434961376802404556064227852669513372794880;
G[465]<=2560'd1715054636911677635422294878265538158479251037731161574604105718356279101409783205953049692816438299118657994374097321898870286526331013614230960603335725656586616254418120654962298556859794952511078649399636590747283974665215613257068199226126740574921838220290266990167442461057299777591807046188289133133211290556218280942878895589031718050923296314624554398254486439055641937607543557296087406713838944170721268238585767193131173545456784895374440365902236068622358258367343874512162649756470436427878385218819397817602603560152802100305338291256356546476287304171264853495818787168097062778826709549727304950432532771167175317503718562274992634450949341197121260064011034734677468704687164124612581740832367441401765947970012519977497988489419359130780434432;
G[466]<=2560'd6414033728414507668645369341665142075358108520508558082234834044867338155889710105995792856128985261600988745265221856275393748517214419189588307890752554074947187066546883380326881423311668835448145264103047266748949461103272549698630168677559981574403578143000974764554918602723865687680340648467313015841782783612473444945167943677027981711854909069622788569746056708161765984251266938162027920354743680129509268877792849737399280771872056357521492634561001284470606313346236524202203231516574652477184166760873890030918554661468381717008222290060127293292186034814326999124281549636911676365465641302946372395526721687216330900239041770001010629658495661854938130475696917686602689008820980489015641901726211289677216402883498284241714065648402825216;
G[467]<=2560'd6389076400131688952283448737246274975290435855004668385233278674386290748764204230094497276889901313533946703813967616512256509906141360196470898191656577380832601357339312133202601711473785109964054389581026088328713863340002936265435676944495976982271777489413445998019768626966316651603491862154849395272150546522331912853391063666658350323832001889167793429705882870329774606940912017263640027597996584628948686643433761660068834592831429934753875971714149113199151936262500844389968878238166429751829603503176420839539266974076770285930504219411128090813460205980522965913560232224247819628386479829829793087875370586529369191183673431108047555451646469069972444080199137047940758506212253031761486392001344724974849854320286547531830937743867772928;
G[468]<=2560'd23801164324326889450166993203196462049195877899178066839328406206275736716792504664642063710205066084643322872620848213614561601660001783772477809422605512390736123165302634589293089195442460444308410851421125945951614862158762300053357048604453253880916180955048568963820053477240580850934817888146521886579905366237100389259701569389902820802133133427279047268203272587974854588844295034553673506497922399532725525333834216782648932166207752239193302564944008473612930443121924826329565003949005700743238481004270316635006550033208792426611688737909460733116486523906276041058317098804328733833351519965802486548788175237588323104999781756964340554307177585472071312976426155670174131959592611707445871312406490429381380640736521506545565958144;
G[469]<=2560'd27081263148906986145549132614622857820845587151436015033669738248329783679323429629872510413382199494492709186654536608767532210106738659793195730012112395735875064192337375474826263468810581690072685153017114718227072447076279337753460979798624130612745892234837033321824899755954883426479591069775961465157473175112809341949148262702901814114130602573293509282855130693657938369835981434617094344719329969453385033992537978259657599621605978723002198148078542842974230807193307797440240968857561044227388569244428964116502940960923455811308274048173173570694058871031736512792215256899230153606581613961237473629820060525195591507219258635848871405145016572505709220268130159801775096176868125568143990558979713102273766163306916850878664297910152278879836963747135488;
G[470]<=2560'd6725704456905100107436900048412759051446299402703714083074994243017234843211107378434145240430525672609937421601789231315900479047501268911321559462641114195026617233795307896913564805300462710388341959363099802227515220758684483681310646768843661400853022354993244658153261904180523366887949995853073212291435016647439759200387183738751981927622746791856499742595267172667444824245488643228432681043450662292387821621260833006625257618524211554687692483898785293199283031438948853715817889874169750395269592259370764662079808616643322588441263111486645820663872892665550719515230323653885174085306026358436798135165450985959914121447509581243964168147584666914205071264400049879816013129857323534572467380493525338767337911394834063854750815642495974100697088;
G[471]<=2560'd440775767288133517749010930110449356177159600153185550032804136582307805670599195049081805596033928074933671021719689768955141780051054137084572029904856521059186542815108973894817421991055897505631055680565700999994633116682851293618142065572897356338973862059602226159204836977437376683380894172724569948986324863977870090875979399922672476029345816640235462461081256477041409118414018083525460365110255250530420301761340596320729697006630785658312821731955024445406998197917856370167015754964133506517734395657592395104564815111739166081503358362543111203460626020623946469423799277496124070214536286660603188220171599657082598483565120385783711173526425027228133893427828268134739808433877543517901324853048080865902894665317565714731471079651193816895409094656;
G[472]<=2560'd3611274132885632135436222191347075631203118698096356600648985584328936621180693956754555293180823117171200928931701583157963201801731682546419537612132404030768448834542013502006923758251949339597895433493491895572169507480979610486985863655617834465050224266790704744049937662730905926714669294747418932929313686987688225859757041087127400701404117380522359737207119131232584467932551479850642956050114134392360148804254513796552079760718214645274404159039969671959506689988104377757742933399398305785377907523582528078851733420831435337189527324851923499543710989415288240646048866491272997447334534402835443449000581200240141953695612846550736255799237619302191000677862988998946188262230191157112225784309845513641195804404500113857345825931690912823450681577832448;
G[473]<=2560'd86660014506053368153161254918276319667183510037263371593354515210027611401429623672625597215675157899760712413517760997958564418619600281571547909728778637084935034672857251246792839693749112915548145542685818444857227088007325627714861116120458713585499209342042936794773344711861045748706322617558313667420892598163050002472872269106278851215981414249468888004607957032695424991168796820876406026156325229276845529372747709540454003415212121226887004200574823528865633380773427304154210251210589343527590591761256034761211453735900983389447241636888557273854170796060545411090024735814376945619075864618963883369611255492026438758432358144423691383019478638445085191155196951802192480187198032396200776404514624159056813851423807681314771815577878047372027531318263808;
G[474]<=2560'd86547203451807617339068553175111847483203248429525817925444716230171122584077505336460183835223075195579935896647589667133775787201358275844452731613147779140537129034247911693420752550806061261973057725215330401409033465691871697803938914915113655263068197542397853451087989555341815403220522928653818157559322257963330167563703711463263885229989392884626068605532949259865373988334412826892472021864256403583468650143782602648661390489452248002291690504996016593855628566407889617696074888433589499446425289001575419692008989639887918721426629920868010780816114891291026836999302419840598272887033660707446724120907226112954666857493306230856824389071180727798032686032180872448723532096375730563949159544707934969684197316312878433630220650703518345256768219543240704;
G[475]<=2560'd86547203458561133094776720231015508752527147505387292460086214498375829629551932836911835896275577965464817477833785305598060528996253468261713745997404624106324712400663521481105869744200456599545208802379383745249173190579021683556204429920843148106805635587726913121622068283165672293431221898745970736783967907619829920329414359650313262736283960845644333173988129907441357031578420729082477973058688921896173598136859333728585020920953187522436364897995680844932021656549708048061875559008927817491694370254625643475023601763131742959041611675894143951646797194990810082448650167324845751021659095157708558113519576871361157719376055521086115566083615468799861375315452082371507203293680567223302095129145936686004225646219965136980709808996436443775759674295451648;
G[476]<=2560'd86660040339956985216789991750574140328768130912269355472458207818984045659242915299202783393444888886316129209690444801534067555373274285471098050284345768275708984379388765837105087551760272404179220484070260130423848984123420891784999930833374510064246408335304760194229149234370843041347818532553145446760503689076816956538474931730074912955624086515352456264005203796736461987329127371138970312808073275586643080160221521900215874088308087151430391115296474578781618123520388513670775318258078420175776515599932057241243859950600833313192587521907036116654584548033271934316221360383456159751925767842149674219732180632699417586668306525048550749366162544818630319514623358779834914055883641368035282951172861022683715669023793912938725123934282708194077433273516032;
G[477]<=2560'd1805858318579483045713064751585408066448987035408982917159919296859136304684080491199319840028884211477879684904936965410629053824698457672046460002455490771828150619974613129930207826667483937841491443815951129866127363063663545412608666566569821928635736537937780622311883129271692196759134108362436883463159456512173844725107659450858608079005740265757836914332449670325469891436971517070905648850610917734224650851319192168665248898630412698243516839105536130787388163133433573476694244574042723196576410667036292715412942124393647446949737017208463247622953976289183220383874029773177014767316834831289053281762083789570306801714864489694622840786445210029846334231132873311309543160930524801951663805065014852470136048015129823198847267693330523168705110639387152;
G[478]<=2560'd112866144911121476921100899625632082105588157381888021623574623197200442956829560524984210130458348608351248712090132552712238043179535558533917875399335871662421718065507316209705643625770185742532915013819940976433564500234704765882291728500020550758347958623217325741616103375150028570841505310007477673497964698261959530414947711685285596189574114939471200916108559784974455578569820721371883303329896325457033586972913269076510382460973800773498364929066777325073082646511761435584929387753210943856199219958447228804208457138161337743385079455450588125736176358226757901739853186090513075773173209048583176523712061455822838726734883102780071544996594068497660603192058808262103769048285575963471392551347918787674089642989113900106226041334102416047266078995507;
G[479]<=2560'd115539642779218408837167996247844404590773723290894636235768497392070131583542202839647541006867163721552951857953958893643008095599012651641011047574416935525645942940295295744116384358134284863418075126994816858464399063340182012047213379958540768928600247887661459645745791833523268686004309794539286451946497927392028946903612126949942034099983131999773666921537807691959767855179479041048218034668377844571240230257521067916534576385927718641842697195122054586044890930611030860817781199509136680249627942525625295591137684281082009408154434385329447583426483470264273005397812444036162345925851753017128247558075107790400808707708747607676396549657825012208205636679800160006009986624926029824784248751525041306101469124752377495244697508595496469801708650741370880;
B[0]<=2560'd173320084109970711720494289198052211650740438203027516077689659649862143493725683782486328302616943953466672165309524793619658785190347252447722591712549664159625675664650224604670752595972979134294131742828139792591649887812380222886897358289271213583401051430472000582462636123383600877940612198146546979821905779710513285561350675180051651882002889447609141013041912101708871061651780089771477575643289430630959965066442758212233198347520473616549188506370950799970806489509943039138652694681329579332798938950494503403453276383207339292204766616315269101009651104608690998598991291761310838010038342516524812817511154628610154992468807905459589352649764334914435793507328479851263766351633550541905524756866694157583001944015264900332254359673123139716386759774655573;
B[1]<=2560'd173320084109970711720494289198052211650740438203007828217177875666530843338786299118461633778026724839448259586163977539656354413907908213964490148101181445934151862392354204253629554080553630890129571280110120751109176624498780428731894153609352810938994883454262292413716286976227422579580223267292983168531976982262009542056952689291446846524601802087596315512668487646449718980882774078040283055851565184778880974058429175830081161258965791768064122521095177023208580855637293098233583236563675682095881999746880973331205250941743199289043565234841660968457654171980855351311515762492738399006709550869252110324185462090094765311427709923507836386986373625484119968675000180611314502743993937524583724482881573659973269545366706702497678056132091484619034724968781141;
B[2]<=2560'd173320084109970711720494289198052211650735795682407171289411421624922929077728256950965120755952274031775601325178452213485954039079880168231486770553465955453278718862492008995589414630454360645774817356161131583449474932157741287996027390474386105784278333121316187891408794705903950732980314517118121036057291448874232541403781139388079835184605789087491619504080161733859863532357154524871971910117849930088777697202017530638983907804121834482584329134662526543099210364997618357118855582254736038495194188933042289643589121927591183795542083562638676464093514437885312430341970199844406038112952840460704159887886649544704081989663656881525449554250888067250614732856801622284760058120225434035241400728495756031079825331007319967999795357905798206063195050273494357;
B[3]<=2560'd173320084109970711720494289198052211650656211002835011869433538234118271593113107203110399624717875276984167660117641981658420861943254809063404979882881242693314283248292132429047712111767050893106652674634980650474117971848043216521094905168188180986133147595269923345254520624375508412103470553586815142130958496040808489254870241819882632507776312309444070891030039269527238486301692773546468677102791248827615519713574356422605802866557634366316444247561671834854844890296827272799466283411776477581851734190946756324096269658424558715207691313622334440246628206856589988376742645525155792089973721877495182721364186911971271784386756103510241641031230858796735698778418217731635356110335296122644750827457913147003065721874409187974406066280219394099972230838834517;
B[4]<=2560'd173320084109970711720494289198052211650656211002835011869429223939992765489752419159223103002252843797652126980400914265990883224682294223179967314719456578196961536109441097761953329378960113936256086193727845082326131786225646044397342485572347097685261275307454163737304473711751891980430650747994681170034954417847249008275933726992489272405385393142227390853208460940386850133827199181951510316977884984601626006458513595637208028015573849342434615979866432820259245506730890772312872394732729117484136302715786981642202891521116921240321390101825901992325492692673821141374664240869798532536090861951577160167496322716539362061959337064076467535178518333086135893168599965311410348042184499095680169116387694867825414451068907694208265423747180637853237141730317381;
B[5]<=2560'd173320084109970711720494289198052211650740769724881738649047274633370102096933092344972614463431600781221786003800645802921504545159422768568658485746528330112212104840729118515608006659841608743032416260986514956518068030590018862647223707791966316094548498410768842675775119994034266537517599926764508266619312928627962384235186995929135615905803225444980895727814870670871964128251421568453632258509893393701286156577704030973396331625777782815842965930450755066620901783383476631227714187158642999226250972406609199340011374400334907226807448616558892554578132852063441376280846214977769698598889307954143151064443510130571841227007834220856427011207561279346698127615934242432294383087219680914113790084618931841710261583903512187969039016553031856488372616434111557;
B[6]<=2560'd173320084109970711720494289198052211650740769724901426510732546618839062381307311549436799747381490226331993948465845761319110480813439421894096896605589110748448856432001377352793002142209792041236928805570809311535958656398515000995343715810008576502257137890186512469790614845864897665141857229784330822344387321588813332643537535097542742235948686158125111669330044865983280650746124284191076491452311331083289897619896966700832443382714368896898364174133862735246990975705488500555983151501958246980296081795943929277975369382162635834547167854602139311585554579313197874656529716112098833405335907816070799598030439617905892525580589735383991658298412384496936849848859452346983495921844983167237157071773391785523996208078032841659479293388859974023196822683866453;
B[7]<=2560'd200401347252153635426821521885247869721168684686909202470915545420030226179911476063947707838601313171577192558036855014346861151705121824362324650299578309066475891496557140242854383205042922495500079908101005000229137475111622946096447128475205288646500323532461757842619763751295952853708316044682922920928578971607385535087434087391152370857723337680033841590464642214619933896652058646609428832201184886696116692034158221496681774354924911934694325479423584797603556665847627862606446373583148010277047248256514966229045279613073967703537985522208811329240538901555994107333470484515846792873546839985522376500318293824956429438725318876292665888986199298552505988028001528806509092085781252704353192760778512177900104894917030201800980763140312312817644337687254357;
B[8]<=2560'd173320523163957658884746577599613645753931379924037761644977758647394904611435758102979031047081113643955744970526108230722874397877171552395173175469590598179066490577743646517741445188837686920658097068018434467403745747426178892336773137925072715595714171724168554228829506716311758171314527635874337350260435484498514465978279559075426233528373074956611799594732535844501781504720875090614979419826618903074310216395468845237588463071468560998144272747349986269992328821555304130032444700837984300031680752069535950655067517887277110599031748292008695899986916839533465989180033792174200908564019896941325178941328662780789903192060113707329890573334783408419601982206749574491946948858938781889244349731682838390268069616336433510998228819107543858631419126305019221;
B[9]<=2560'd173320084109970711720494289198052211650740769724901426510732546618839062381307311549436799747381287369197856921960190968869342589853960468996549745257647175182812605221847920225120086933282129971310881270040290862643220720731232045558231021267842012749931876105117626966188938099456607146953504480516630532801697068692121286452835586527257368851217656097421761135853140502591054365709484603358108176978264287909661067843557948479185669453215881801198956977853021773563115248649440902682238765939674084465164389395132162708848565214101049643337864764995823434016041933102467353940372296990598213797876069688304822144932799382012192269585192701653401239752596166838710453527945662914086124605203597456821631768931878468899548513111176913082797912919750461042960710866654549;
B[10]<=2560'd200401347252153635426821521885247869721169014994417274403034507028032665878386578979036299707909850187292325576579854144088095148383967359378295581048705845345020116396494520092311992684952128268779878697509572184128714380834333098873617616820789485581787406969975574094829380780850163731481632821426221550781540234728866176364885117774020693518157155250627799935863444680889722529316302252011040369345106831943559928317468771741221897736148162085805726503691686407476202725598958298212163109158488243967775710811935184690120474701793256484874935746398112285828731052845016104821247477646799918944323542828139766561809651798047173646848922910923445935859988035807433090262174233827060262281078967440503965401488499700207491575036426067945156659432444767970969109761709397;
B[11]<=2560'd200401347252153635426821521885247869721168704116762618466922543161692555101516325990059681612906655388039179250673262689354350391700186230617424902563442013915189664886328208727662100819424090694873573566948189451941303108491035728651935490557701746080962366028684961361231017024306382145665947320297731495035625210506830878010687135294246527369427453814629473511886230471316678092424421235620052025129566710308516866054826350190020636806011704493174327419315393198538797433301204105997967741069896411356220885170917441371551852210927882162288480360859155144570348361610689384647271459347149881386518771804887855085066970364956823153510684290301844039060965905995906544861056318284607826571108071313341224580525069810375376716206976106380567470036769732680881065052951893;
B[12]<=2560'd200401373085164097894249451940124897460150689080841067542559951706738176126645573368964979591303422164224614814878818623624131201402926422899814125867230128279605714292471595236597868153782055486898765624547300972611825249927490994020014772343182299470570303397204055665180171799685388300303296509941765841867075022944509537605897220829853188992873727935520040869516640546485585121326153200561229423339757705188234384476124059038579316489566555701399011888652437726590208217613777283893516889909160942604417825332305441336793727814247142241413471164802365732755834625154478490254952683415684269657634627833617829870629907267268444825546435663845700508875931234713870616659888032580854697190953585138260278735246955350419305949919497211959459033202541560378851772333380949;
B[13]<=2560'd202094365258832363251073528361014799363143616950530887857110288807834663966091138083193597066946990191871578463267022968701832068015807109584884280919909739317578598090798183344688820761532645117981504946118831304575535865765233976099462256766640087730500785862484372482381606198218629498730480819586469417992399634158113796384370088049735889404553585954725441980409548607234524515605669842498505872079197717592827615456370554513439244794165134815328969083169202305034494514275910532259257488804659124671956930612520653832901373006188431788533006333095738248298312045499898731536465704984700666702551050595464870887807329356494027898675241202229631827224046445298535942486921714078144467745907948096002678197675596354504510213157621744343169298057797645827818805584549205;
B[14]<=2560'd202206763073185489371305093129486162870557601501800149222705535682517108448561107281864280745756175391680055396128989493757594580900534050338315346559970848544348667748023639540799726465670045502851751184267890664957525892199515257516551196527524899643056374357330464072109358746362111612116079281568014287298970225226495910831112803538401510240796379905528284836214272756241785561950754318754301115628830688535656941702780118507644969951352821072585269300747905058307050200430416981087466763599360700306012654244025436695546726799652338968806209974422161016611520818507566567590683054483459967131413526901759955292818654297882723488971613554108676575268607598513890057267651957856558482615455919054659263068564389337474576637727596306669980580677242540589239192255812949;
B[15]<=2560'd202206764687354559029997197130962491672407566980473444572532818844512543757589941212313017270308280688903010896167961861455860066168196782386318519844159453468990928372821614842128235820202063424453332628564988242106833280353273575125955231951034957041091047423064649636037489819407864984288700665761011030241178655906522399880758896445113519283485912337356680142647021200959432361478234279176217197911652821479967828530579189101715582891234618343706783669906296629692526049263884411045390412684446458937390019457212138601302172663487219647942811555030115324540461768602866420492476942125204539106445328101596324141736962351746238955673486633992727167869832901456245975778796434998900687795762319488312864730884235464262036682171329586686509173173992945168765130336720213;
B[16]<=2560'd202206737347365941685899685605957172591073776685444504584833210288214858210914066515337542372412565502417851350958559882283507699191588139828183333643568712490533874942258653860139393897698628630701863617765036357778007505205712561349224253019686227270713170333263154764354692534122155497107915922153194927075589296329947938063897534414962612527759516985239531099740793274062589290158540277996437897307332900539781529133963096408373374315964172837105364718230091690635386487893593162337836689837656876811104271575888619336454546060393740424837858163081121314801275025895667964519349456220239073751254520016963306873624449186740573647459512712735619987816720904065777229479042966275933579810097780032921236735007260332520191665879902731229744490149402395420941548571153749;
B[17]<=2560'd202206324120084109060721061228016999317482614145080895029048720817383419099532580320460992100368257515426994771787732191163848546878269069067793939406647649912808583472230369950638807110736820223783885035258614210731574134397846643013524491823641745824444964019898550020586401867898657289852834028882876176651059911305392514268775602752310347677272750727951413109185771561628975058205686896011844729681908953200559720923525228897217468680072575347946794771590436476601921887815756808243744268482383368638371215839922454017771394757267705305423255447276509009955532828056531932770761522517955862976943372123188452944568065662762067883798935914999194827388742563258352982724722291309495777831575032403106623284133352117950433154864380249576961012289071741894847335916459349;
B[18]<=2560'd202206351560958293258486829253114588948932027282526915976112534571305819353022757138089513017754034093741259564706164884778867412575659955293866130895869457351930922656246318575721110895216713829077962143564624404635498852409837494098054978440190736244286042557996443369338924625398384984569869729330489674239173271176522646432866741892358088985202647757932559934202085578838754395451275041778213624459564497273561746363141413671098419350851606650353048708027381340957057759640130847916057294620059215699304593902319918021900731090296526066067036559906073602319307829993319763627810157248838193244718200566278376384604870941332758534442272165186126955934511966195006730139200857082555259288020798676368239021752894463366630436765006350024286643359996807042552678455792981;
B[19]<=2560'd175118476681380480695633350018783887950929558524776234231894537431184475367025408469812162459021116732112717143580285115201097254154848005280688238998408248568423468841338721919793969202370220774733761781794183382357003400368443615747345358218398541415002977642448147077732231713832540602676411810443149010067134536949470612430438066018421386515043266520442073764958201940866943727558161088570910737346880461952890440172135653560172563418394921972207376528270247058555125971726133459232373049095511527692009481752472396303097634409812499401259470557914518048104058512393722064865843901428793838377174694046191855776601470545267135212469055366654915482407861601612175177247890701693148897339815065731130264824658820623814201281290944507971528269658646724500390381272520021;
B[20]<=2560'd202206764694053991205341683005793479875459109213430060727411215688381484612609884477987386441629398044502355649380423635405478018602645723838911606854817536817329337720388405143486161979589542139904129652882540907520770572637658056528524314642042892891435524465793640685370907487424294218667439723534803943268947631329664347493410101994414941626008864884574299818506554944998757993747670464676526470674161380259422748542126063957337412118369106094211525816821038706566314138864469801971237294042151526000276970526397135236039400994350840431269910851869011263352905363054412063272284714088710293490814023622819219093177618246858020805923398232478744037206505032737992562325449327666449942547360492531787923646444870511415478074741448799766363770693485727181275154091431253;
B[21]<=2560'd202206764694053991203873604789173079222985986987585854055255089095592199791430278830818902151814537576878727521313985029475803010124289924853140585069521477706288710074053131494632428631665105079220670715839372924464720931389669166952089435577870249618830015167341466263656367559991908467413600550835202379388925741608553279222086267917995224565795708690032966632344435296777811478555010461982353127372284575461676076385751144909496715695198209515606172352914423227734242663258934779392837351336377744442985256590022264139356160113228077715234549007822842547060712557925925477212434114282091678926063371122536541941105193425843957854089156766850959767397497154706288464289186133830817929213386251054309430639086785965217204489750712846956248562338787830556024092486882645;
B[22]<=2560'd202206764794965728113788340927746986965382194277223847735606686154726963563255220994637680592777097684954723693382267542578554674840752744378565152296970299621213076697571808874515081038200299721388278563663137476146874947485663393385114219548720171247574482142569800588378933873500812740211976226985512617187903710375853244335017827776961126508720211990463897735632064993783188647781265172240412747813132158850730427654488433852176465804226992112594936285154241850730623649240432388810211419579477238225779938276315040888029441610404090970245083238822309590635654704350162971763593888950654696306075679081211599926320235918414065265943940748175030656295548194024966569710666216905819798992186936125830428696820616239046504844924781348009259917091051955607843548014400853;
B[23]<=2560'd202206764794965734127042450885099919034897806209601908361349453718964527138527363265189991015946043781111017212354796297537408602033559673564186141583754985253857896408074285929575477353009722076008238936701384860367253412781098669415457664699690478265904892605798215559855025211420753152755611755628082349472137811925362943202852346180256662406524262717458043773939506482581346934047468536047903344918378679771571789138995596070934624406640735750757768988530810790233666094930716894138192658868384524814830822870103456850532737093536859659168927090711733833398542927331332716321739737361880205073231105952745620602865607005344533886878776446440130749050324879329112641417106140466549904084416160730281289247994535301181180683518392850707807324178164674988815093549323605;
B[24]<=2560'd202206764794965830340570577627524862807700386753436559830869444351888922235728940854246943591064520341447639407484166105069219431530596737258412150665335256816557608880501721021828903202387510441557485899136405817262231570953321771895396441720414081917989661528706580537535656163681205155116752504050138833743682147015053961855077979923660597533547544181638884091998165869819108385769310406394684260334803115093977926627886539109217493606946686852757798455024279994650879596241943477767998902669254053867672475793670607298689713119459177745169207425461480662379367042629441290941137361996982688743183589473246123318401541688344963275248531647822267966647235040492227713120546332116961558487916964539054526607400262859806800077443944528801702331321555504773540849112143189;
B[25]<=2560'd202206764794965830340570935957553853322601790277296203371776383871900720459248542889614029063245474688875311723092753928932254175627724874092570825664657921074681759501732290115082860000243993441314899111402999150496556188635124026097305460020028803532727478693206965746321796346844925332987136869101002265586296130548585475817388437254897696916794353549029135714401804179261043389002552546069574638987198511199598921257176545515434262717188868714260105344919822839657070608945028974326551732390730314830884211630905859682056255887339743098552116950054220018891911476380546698041359633642632381868468936806026801790459476912576652940948432033087352922194132975483131839226758415199107992724552270557490861174935824116083463743601360707331154236173683949920796649935164757;
B[26]<=2560'd202206764794965734128602666296483752766366803903774546222643735983062346572858974301194829319971448700548002944202058768914177453150338067526843225742171867010760695139250985796606159536333124743625967887506081590291271935802424719878624629321553472685386126957589277424149966746432682914826379078891143934143439778031849931356727965261192341556723641922084361525496492125164067753240125285073127034084115579500696540761645100115898184053640165585328784464815051609751244108515907473351336186574387875141115690563520253825054563716691427445518434562208130556235162728648198877875361861649334503627788448173918299239648563382259346077991975820128398327655253884374972611176627506818134981335603257297916130770428114335539203580184694523270810904994328964617988365379523925;
B[27]<=2560'd202206764794965830340576670731060913570883865082425131680936667570128431678221175530117082635184321444780559148209091299416894870318126751443907622535346349964817798734555331478869865150276534151446570702692783486264305194151045933944099535702226510203383096796437737327804431472149728330472144097131353790859964460315548570611650782519219413007089245395744156433699349077555362081459978430349115773779527857492892782307206290949670138646331355281108117219912587955770384592638408496799553671064692727958010609436615500598751889366416468500196983956401558096516500101125188143473007404457973989104062070782812452367217137384591555664417254131963385356885616686276129843240083483056741094870207726725196971270209981276738586552686648779818022213005794160374977727084975445;
B[28]<=2560'd202206764794965830340576670731060913592530898012365232526868639179977409166464439254870778110385053655797597082796584845005721252703445465551153204053571054089714574508283436158879835631019559602425181104980860615405224781934325348713103867546291861009811291322806813114855110943273492806527181764764905434357920709418518517769558304326401953102116859643409362578452588026595706710942032734249723449001175896057252967822103421969666749045574487650026941014798927657020532599165085098748110987687867481494969022877689796183309514247941313560394538030041156742851246474179770973639329785808174482890467058475752895118185395573392808231972880972120342541495303342000159059480876993391254933349839636810786122285437943644144434577009684200582372923805503081230418330535679317;
B[29]<=2560'd202206764794965830340576670731060913592530898012365232526873223117485759416612622059346957163770798462417627511728926167378575235605039908410909435594837030679680986503069922038905299165546631543222101430470105585024950752339979648966796385251896490791037316745935241842490651940632084298690969182316416078264323164128548019720021715262012125931187434062114871188753234892551914103078541358103546074968225734236864893725398763788765315613439081033969371865917055886317976096728497421095516406277859829814961429258650433347458759985973617785837061480923673498490389396799569230088741626687341659444501643934643458636416918759444514994834027042873021619311522247676210550226909769310470175123349851565439961475116151363684044197666582997357209151332647594557944750551684437;
B[30]<=2560'd202206764794965830340576670731060913592530898007325139935443594837432993897933044017075550681153738200387221787310719327124664086131399251798035867033545295956260494446326997196117426185885165705508143178075239182915128762006991837379391038493029871809979577489362686211634537428642843000349930161369367177879480807798087603210784546718074296865267501992341836029346632952365900241824905118126348511171821763304799846863398027741420544974128410004060098165479100269918056024530108742621364446193330022942513456422985273224008790725666692880762712706251524814083057952415116830229772829791947419692477775454901458593935128456877189484404712797446220118323095897850467188381902405401703784264351199286480321734134813965198742092174661365016470492814146265905209088803165525;
B[31]<=2560'd202206764794965830340576670725591896054771962012341924175949154301503570762962878126581705134155171928672319628189072367984495784412902991321456192369254596988583303997151455282670754393415962740980741037093507627515194375265405715629119149619081126933992012454429566675914136784868623683933898878564751620546530199142432362173094383893560279321979098737451197976410850770553472775251910618231413291801315393978908397388633883256414265374682598855871562385904556441652726399479385908630208439989405720441913928630974519077991888697202802762228340581734348657870651058656452717536910705317476914416353845892746584151485677628348141032842758520247594028341001189776050297759876293938563009737646402560951945718599410091148084601906348502872726078786843762935389831260624213;
B[32]<=2560'd202213789659151069214043671894458574850299041947223890957517075325885562316819695036295687403170701507946964831661644084765093600632223112209280227071536599368361606593020745126396409256131875673116298634078449586968116131091854380126297541181744894425584005961812060909182442945051012356216173133745064654503290772782761131551111630007125715798879559217626349418720312975978694303552364830223540226375051660545646430762588009038301138116014239842354612581144271439274220886179249564387558826081831805300574573828097467740571700953521940627962754089094834528454696441610047269878608928985971761931539671115560358045147851073939454698939413018137894930655570304365546149288705804023426174116947507037947635395526980159855296356602101728665142828668168073249983076133852501;
B[33]<=2560'd202206764794965830340576670731060913592530898012384997294337231972585323167483170307173062653365130216640577863230090429368438819591775249374909354139588700211729936549757900244436497870145546489416791395229750207099093101607983013756853022684515691154923069711448390126393938191839079101974517431611164904761606226660249537051436741065746603185263455081545838839180461095947106680490904381235921169231038267479522230580720507292987147771273382453206752173875501131326987928067372043611795385183705076781400697555543292861697869560650026492294325626321032391845269803662903391956950458900243424239623594534727015273205949978019735514774608120018018459647275290520215774056869082672609390767261323664247481656738713992716314396612377916400341039312378422184937554577806677;
B[34]<=2560'd230980606883535186778549355461206300292360907320963352522779985782207697803711283945714893626865679090884241643704347673776871908449511536959378316409430675073204144070526218839236068166454630892323787798856508054924246209913373666664508248070627767323666257530698571102257008282442187299625587086000147548714774040348043654152591978924069620623464772442745826323482850423462687549629219351507105217588569223289079479164259260357734838791930474032603988849279996390424478781149642166701438133873160990203820573824573409984687262481572543466301426045860839338029623067988978065616934535306088834234155097795905826704519525599002763896581219127013066918419361988410989756936029662133393706471540871869098075197709162859141976806307455926982653601392339528675591251134076245;
B[35]<=2560'd202206764801271178268930936762316680501913123149753827190975487463661199777358925810981294323799646496647821245805502336102308197098403639573037052433858174412324867419580473989761035607089508834678848799142084440366795484425247254948827342769353384276185530873746801658068980247358919524210748045343758908533140365148495496781036966449969948682953213311007586069015325565796775282659732185660677278706080827908704461756475339391176021313086760228806741587417008084638916283016188075463495042335019682157423707604090422032158811604674481441818377803280662080156916505608134055253266636923806462669988664126248211993916841268074257229460668187113722401259357288382057907262895418997781618551746211898712117243729262951286793220142526499899246564529312396745872021118080341;
B[36]<=2560'd202206764801271178268930936762316680501913124440036060349139015084950453745997695516994920340135407991105864857619787931895133404820962655617909399275944743160680922711826708740477261371339877461570474185886358370851010826408937795610794607904852132139239203087262847538553786868334227603944547585616971647952986107148239270808518428800636215221264455637775159704106527158459570205662549371784565474165512427778339073049455312968097079711450936914370204996981357390469665250345335503905345841466939390146343014626380696976332863074786593525553852529775006503473214588459132960444999183640317612705053755290879495441234917666080351850697480410392377392018697227101672907122626545364416306726692067097928069497723791856096873858947001493012707714931907480223917370068260181;
B[37]<=2560'd202213789658756984968613285156043859243580661198566360044121930020105273351239453361281613503872080762900394166572975866505964548482994795307459892105285897403083648388856164074261385752847214328718383534943309802127548153957709790755618343411103936613437511085524607493711202915571749267030161493495485747661818255283211955740794981478503597159908027846298782984025777353096923582212786859424668568333626706147032013930420727033378827701895238485416859337754686093826020198055328497491711486573695301462739442985238411219942746475508334506421128850078033152533258691371602090376375661631215725424820291819527572812130848981865034147882361868745772003457379375096549308594292888399398950391101934025570724823345662918211928203736409084186730615823970381730078981734356309;
B[38]<=2560'd231093443758180607991387474662494864812347729789283720307827626785656952178778992540103747384500298034675207520620816370866966858999890350640112811467236123516148452444022396529162378014451296422495308177140400693430007099062276702956735145515524177210851922739187141128428738002206390329125989313577833723460812864528269487012111160929920466227685506179728841102132281619404420106611342189476832716936683914662261136013996087633744737866010210386574151254313356318983795201497818962731922767176749275182849138740030742823516865435658504951399615892564393754344961989485418892373567456907864458645098971789329667222419604447934912279533512117232612767076321934265703365976252611311379753527145964038203909698679586148087195372319371181228736026333150833352944706666190165;
B[39]<=2560'd231086420609444089875711220739080518513263554924192661786838362990022805210938542442883197913807466674669632995953742548453919897834784732358561777578725155105267020345760119178318534472653622079522565098902111343619379540862944517161547056878624938733232330682589276390869127292863228153753553442364961974554647811975303619424732832155405655520610031648207321802112549235388675463052008983403949036751443058025307693060812957456678600393902773519766517432057715427538695761694794067099819797664480771595173423030990477410602403066234032415431520524705519013522479434266152548266888435457432765541365287298656382578546109834584079020632457070972799410049733963710784097236382323928263370557239694232462930802950514166497105806834415582887070876889268832268332650988918101;
B[40]<=2560'd230980632710240301317623020884896050788247970985722704117576476345944950044006658452649678557118560925530074299881074770088224814408817728593142648615593306364671731292765319779960336735003549097743862334973791878877948147300147231962332087808699099079922151871899606887198971237597241766381473562937172019726091161336332043772026790214325077382662751667608457016639285689497350086495637152505100349263924966207066179277861515420892382009250448056775697601503553684278090500262019160760587842937107604521581722863416469821055166964105823549997350229652997475278187776483116575653333588601006740227009043524256343504742951545457159856124876155318428501119749786167707308693565705902260588780532608505093013990530266459659637868202842913848355373898758821045194294975354197;
B[41]<=2560'd230980632710240301317623019484827561121960356270018311578662001248674074771633495217158703861449486411051716828058005454651590415676803020329043411778230256026068265646507529730496748562278470326092286013867114174379936069722939642430754501807280803335562555366453765312663308672763136632703238049617450685343334734089351234651716435292801584907022144251524680328723225547325170777627695064435851392292240077877511243273957793508396383418120173616470254918079630814309690179341147172122209228335386172453396963778756397315479674206941732991864170614273571638759088264264384599608931811933657856485159804129596059900970625083362193911975153262059963391419535592711013960125967902913815143824213484312528422232336406624951309024758903806647700118321023588865092669414921557;
B[42]<=2560'd230980632710240301317623019484827561121960356270018311578662001248690213474753987975259448740392708518328148513088837213823943627622563242392116261644552789163810261487488399961961023629096190375498949001620633265131129996540372657649903920789560426818129757043996466597533096515216931769532946169620575392726961671227914318807427582981704914807803606791241767852633910425123912004083571060279449481313494260243094160539104483774929076915417290214438869782291161699920479971712632912160641953186242298587316859246173435423224555463257868075101117198653446272802338565607541220791426890841855702876759522643748462558597805950669962638226727382401709956262843175133819348856033191731506849251416718618614742312083936495328274618395721828657245554670758375077364349430748501;
B[43]<=2560'd230980632710240301317623019484827561121960356270018311578662001248690146769683720453359121623535762570994545777749603774745696489670451793714542233074466321864946067722059195346867119807886347995008639007124777726346459113578995306720582582115158593309870308374307006506949116181517266615481418322403722724249745969183712000563364965996902692255808772122941606041395884672540070335658322667579383855163258224579554683556005543438797729538801847470369273956009950364717525989435600141153318775725433112624890342516081704579824011615859500479518872252318864798367390336429516793418685646742621458672538583163998848635857365783821035060740896640598623527728776819519511042044622194448773431508618081110179687228451164694048548081292522083113176975993261808482116289223284053;
B[44]<=2560'd230980632710240301317623019484827561121960356270037999440347273234143035056007480543284574342029287443019963185656516617056429547182668116251109140540236566212629350042480703419611187790602650981444967870301378774377207752845990956028513650860992018988266716279780253780830475805824333249913478216518217823280258420787835889306088911403710960148891947901624716630727218995522604672980881192624464283454414131219141326380358253020795737347060975301263418128075498091728625384224734518082124860708286938287135488219114325864928763607124751434361184744033228568458240648112268109845110681468197424188348481876780860409707513951075139784741207083071518315739599442749742845744474285995979711795275386468897429520311233679407442273906461639972390464731850360279050003923948885;
B[45]<=2560'd230980632710240301317623019484827561121965330312492806556453423110115847462127980444132733763696222179599501004596644278598577028957482352110931636662271349589227513989410027895197517933609779605855678601099885232242353372253364289570531350375154051323408647353195843573588892011589698395056905990419364140532869061652728674129421484774748901868656325401622191296296765934421877802273420780113309147324957872225556060712607900057827809511956597927005161158665666693205145285011169722598719963628622598465679271862868227508940635864242777815737655094648476924426511265417274596858741686218755069953119739697911929252896933060651471367056391724285309725159911999871415926021725353732732234202744980873929468969972427539788805025597208223587889512425359280864975577773593941;
B[46]<=2560'd230980632710240301317623019484827561121965660700938835986305444039093455807109537437885590747866579962162314825146821041641674505677533985680697217271022959768652509860879536415161015532482302750315562330487548065557828443363543324846092413848003406914705825907711566482091675490910804232076195023598757137261234857991267307215422600797731177226789551140029880191588511045810798646583713217883850457446887953966224549649420439107868549445413373474661385999657222268057076400996077034166229018022522345851609777725599310800701280040321789602336945353214678377732068368577771770444510533554066651537916047419077215487575926974023281994782874470863022585005072024450514749811323484688914622561576681478389725226000648475004023599918560269217480368029558864239760306129425749;
B[47]<=2560'd202206764794965830340576670731060913592530898017444778048969537987518775954198568010997369232298517219129125398362372040699510355613824157315323684431830756980173069550102410701758112125518452707074888861589083841454384496379692798126584658267710178255934486994261553582137075283732759088694268521159480133645728574117466279527669143093731681854619862241472110640869980080815547627551025687672730570796558651974695413432585215913781087848957429450802956254472211023799962844887274872182401761057986875284894342821708492379002884956240866123357756095204702571287153553405511927669739591049845499812711416152270734907626887616124234894202979859555631810871344606934341698231870515756323207490528041751611315230833784325845125113578357874229339861191224463619830845191574869;
B[48]<=2560'd202206764794965830340576670731060913592530898012385074785479413626993933146218396321194082688850437600159446028679498895092464519855123157665711361162644968895105445251082620276088619585228094307185425194836824922966512466252160153216188918966386296654840379422636668713890354214967188512825363196894544096548915105099455897490781808721958369883962842386188108965089803171645015133494468806291513113561391204460890729449936907577730025338922383983209062073117158699893512110248335752183044048786815023316681391378454242359677815384104758447955781616618131810987291511861688609214512217465870746890208027131165394850635969739932057159641607314299577423680272322555729993028704921773163122812439375631510322866249457327938450800617094820076529757337639202572805405865760085;
B[49]<=2560'd202206764801271178268930936762316680501913124440036142363115609127410755432806889857121526695194547413906578374319053867981428627721656597191257775938024876113785604589550235934005740269950326636327314670623364822917491556992716089047571980248684903817494900789977207132821474356278465096413115667744287253610766683817828996404147919284040483711481526916355412525342573626879967154656140822034710545079891761011609181204330524044316675684887065220371966973206162078050597367995118230933084172973692718725445201488866245882635873157549753972196668473462120073959375930951024619074898693220411097598976683054588190780723024487638834454733378316222376957956155740866954953858166377325738855623212890844128696765679908243315541913117954048042121075924133659729616311575467349;
B[50]<=2560'd229288027943454101998747420915437413802551520895326069903936811990357442384865484037152244408839607673113144789934235207007144393645427337639002946648870077974099110006020047318177330981258249790651309000920836558330084584380546307970500945797686901646094806059863782516055469868486117829841571202518779462662109491113194285352646588351057988702303774222377749512776327184201129234286914906740559998307227660611505983979670900480851775213516951581796893338932008905202875226035757601703244666905912811771481796916630693398546972045898374450772817596011378221415318101947841539868729567904683886787400649029320038878602853300129447286552286831495776137510369104825307112309444810992782551535750510391697329698022640392593963979762541840835657279053832898117577036990338389;
B[51]<=2560'd230980606990727737164129953287392767745106125707382919191740582820729121618546105376986743069132494567031022494040271328051426868643440665413682785767594642028286979060289820475927926609151319568806564074670805416347648395654785027719189655560240088649122411341944172081364967152423849030692340671426105004079520416642522587671402925682320577682791435371138035481832020690240695163022980285497964255572911316504242833454190973344630190971585327475347740477125614125565845705895939041623069831504262671716323456075709446425573687138536339747649681104306713116245718679254253521212852297823648681441784750016499081095553988425907551883291247157284422701779767692215517694925425353177520667179313477852337987659190980764914394905587656276441621565505854602049877022111782229;
B[52]<=2560'd230980606984422389235775687256137000835723899279751539493465591981346537249068140399313399381580108569425400925073263112000330453995111805915179495076087088856269624787971414221836502329228877153346054272695624083436098237569305586385910496473501135802503112147005526969601598939085710536659573795437487835832629956626727472224327728586365109396423043757442642108031959174051914568214208290681468255590221778715019273559329257087066094060933592662246142599537019577909192500849789341470005522524881929245530661896586007522725448519434464568656391707817821519614285815804036579591626012978468304842851170484014072070191586256977045622200989597401953172902246368587601465635729777233445413068332603169343701282680387019475229661686739638575442342967927869844151956548179285;
B[53]<=2560'd230980606883536822382107430756044730285608276437334530914845942572104947793965555610226676041627655062009812826874019089776404817108810093283421527553156630463492160591405456178143686066747700312124510584964101614082191253497677076411625453396904388377204674715594786287726219795607507102439706146097591198228262945902747582427228061225393339171862063103047959460478605111157563427685006649006116885776558365399739051894928374336664218065669167935420109128653329514022700346423603621567629942823746611159673407828639179793211159994631326825697085636472771373949945788881087180581782737354918085050766181989739500926804082712365995943574548276566322970662639180983452735911030596441488519558963985383804074674471166032894693421321545199585361688338825494635347784278299989;
B[54]<=2560'd202206764801271178268930936762316680501913124440036142061524895140989611232867655298730268878461102922901801102325947517107756277168514450111170827601597863755433876773673563346799430448234039377166300988894633329498904782732620811765099220952143312264896645207508129481721297482830160081064188700325344500146935530448100279020107757157443421640191213654899850410233183720269370271140749671829842967914405703844911698375694380524034678268417760772442819739736232013889157772255054436752868422555627658168538799949568453758449359159981264111149628959793400976851807620938947608192318656828898876524019318673762300181620292199572868252490524975109001149679091479447832869131037153021382190525849711541620067463777388853579707358834303919157088917696335837913540454258136405;
B[55]<=2560'd202213376437780500295278178275284528109581876271628051508310261159263380567411882798633883634330854010958532646856250895254075285986904922440539630553314258195116651566365310300407500279195864767771949733965019921459950482687030373295862292084019017086862764536429122901483966736348157771955918210308420871015641964114698061784970747544162252813305969409959938157399827956249625253882687357494088592225505378331752660411076643004780042525667553887472754064812857772716236175229541230001423100944119491264455899150551021219003482919664541533925877237538542383422564907210164626477515796533866906624660026534752067526916192243448968986955091146323152806380809062900263893621833851380776108241251507749472665088800443391394152998815423015553246487877607448778966279069717845;
B[56]<=2560'd202319601675916605894340440841684455983341094859630466043351556822502660137891323271203431391660550918490901504971255263809120320389377304575640501143006740314362209937992572785449357437256268099496464309137222316035416244929452282277449485917868749046613997580887508311100291333932280128355543825544643854550159614324454283876331259988928849641945766401472536126279496353212503908414659084576074658938301919562360173081909369830792865695495546059030793983262889791558216840170918772522722512573613163294543382854441694864359098361313050784754935568383511436914682158309363431959569833705080159573521032971094827879647718731964117432480542613332209624861043323112482127331731514884579153693199458797271720517459192998180707415152453796937785717948317480513518936738059605;
B[57]<=2560'd230980608598591464907716166534432588571372568316589224563879358805705756541983582606164723057758177837458478456764092297487094574500051614640926987511686537004044512989973759103444137839167146439138454419476105596589200456023699641851767175788910084086057955772472534487338548046905876163721882353199572253067878455972815390186586308075703466129037823282900873231784392315245881267283950061031457173787061911801578802095817445921140105808109195445425474106612264509516690205785143726371594757561297739985099356866815911723160085273398519659820599060205021420280334853718958436036642449274330359741740195026607601456164839796840910022568517753298743467456180921892131128746340690863054572671972477106532427538765025382399942186429775076639456901539288613749878357103039829;
B[58]<=2560'd230980608598591458894467791257613329637573864758405146680090501810612808658750375894476632701453344129012727127574455216952898108306121757566607261681325372929265171712312067310352764578748399346222088057839052100487415785001381005381072916230023580905598120231264770762734598173727835411881492228867589669498346142183135346256075760644598696362785567183085029018343634561576793816069259515855597241024226468217470026755904647254870431050768697739466641518461112453604825477799114667848786540996882030182178730062532695131632187702908479393817371560785427056596299295860733589770327579283367573239346076461457331723493300408109418262548740077245469434095785099030135027017296472815768830644060448721573153329477295344097567642072939128642339654517410319128450770696229973;
B[59]<=2560'd230980608598615992949306998896810096738172516598553797306828942122360662742263172349441006147291038512609108879952437725225553654060177019037811341771548266207249367615189612786410701795448121080464254096625020955783441251022747261782061618968041778872697293466464501989287474948228441983844644008227048856708373734187731207784735787873766350232194676168384738152415871890209986639183115611159026655664559242736280371254399445690828784161071215529187041177580273269840220720429496716864369602788851673534200093712535388837265680115044335910419286191873295903498155575217705294638089957803234272316500830397483905952734852062895394306999905933805822380723724701071926687702760252676483522794220896217302419345871595097865450257837461599814587936043493470027846211060716885;
B[60]<=2560'd231093445479959306944437454890577626546909842460847252666772871579134047783225627660134201728198309388593888739323707678532131948851220249503961741020036471198354127141592256919453495707627869552096088678368541453349613294546872686050646349823008846421523158881523319897491106015467194279998769668150386756356454054213303272406635839586842242742222881575757622257678158593789154659440678925785059501408837493572396844448099719152934567996252980967573809687304052185869443839535321488005657717853160182693033806969755907844829366289134717441819283213202538654737030402366400709967218827953634189236283361384649561104527434737753912379623539364789612383241648944023671633785738905682237504714582414086930633637210294150460529210989317126990965575677856401698269068300473685;
B[61]<=2560'd204012182236866186518414106772331384000448770185091973254420410939643722216880615351593929768923123632673950781154866876698012645637243405531424017814605470569879817117507928966565010121666996387261355905440656624401988027058958463967356679505639532558054139212143112508916433180380186844930086966643836222856030361562614172621301587163987916842898044624665022461962125144534811841139298512378397026244831831671134276903638260328858524821697422462876711848017278231427712218457374071660244034307237624236076999997599842155232024133851123850228439759047946649827286437939417935133561992308832274036408358415958470230247552442969272713781546270525774241090321557352552782814816476065315677954421426407114523124325684832071052589856109503397961440545605003010606148974105940;
B[62]<=2560'd231093445479934677076941517742998995419104503847914017321446981694205820477650025680859945715074566725052583833341905823496657995274662374502075169198101967055786404443137015169203096377248720563503843655491664574784751706499802274760608973023436184716959438822507306986054060622532506193391189673642489142820460021350663893412463525729557905077694038777752281406533350878347211222358771272023781452575185101430749076318275817240251631207838408166050699296554710923858488205896732216738202014365639733290420717330368259368586763157410240566329534540282202624051516374014440083447808833945375638709931095072169102389036577843106701866049352071199991372298309793859975204216934423045559636887453201127543548817264019027467583404194473217974930751332181403187542240338990421;
B[63]<=2560'd231086394782738975336637556715459257683664107265420008571446264668341044791656985341242791861694071283765550980591474089182737416324035678242718398831105017845825659662326318637629873413218346406582462915703363112918236593694625571497941223235518502469555773165685869166869206619951520573359603415953158808530857724396262418056813440393329349940743919186237451472140702350151067180101650603570315153423327619338663638995010591757819806498007667438665122247233302690358308331015159477730075872245446733085262158719758849748924590011540004185494498906090640157019338077008969281547683085746598477326690104214080358464834027097904367786646876514247094861297585370946457660957394601144865674592677778154093000709923537802102405835374449023918369038850437140728726428975453525;
B[64]<=2560'd202312550979114982409793762949670346862078659531243200430921791033906496229995249703646306373799402472056572873820239422886419341773191574560447245661040154152568805839708130314232835962448878506965880733900069299259403913087631297329224514593736792964385024903803085136968182644899128093530119159141281339531746491851511199716100732820037282076065574030598096191572169461253687809877344215643777775979088212099903931366103365814168104517241554900772391387862742637924698939572768494635509663030497076962216556885572202978205974782945508524836395939638581500983352162688640009853301776630629920578712798055356454470099986160213027938742801022966259774802274183602886435843355014022198800367740431144125817901248966838357335116224549121307346229459575362063081902219547989;
B[65]<=2560'd202206764794965830340576670731060913592530898012384997595854637721978910296941106314967173762525340324870452338729731005851848696378710119314738700498663353194420763755957829354920473500845357271366154682848518692273244535802196999585553984543803702689044481288420423668962980405286542599862742370402059525254979351202934188869796435053257293442151122831462123712977375429159092276509685997472687449915095849869803913347713017206827275984061819819422688790816791222886127849494938357616492025010311816444311183107886012597023690407944484818143768914138668349655708274136632272139822098257574017248699484868195482963575306638382109748629689166445861891961634253960214333221720176514154647483055410017403226730659962274880519489738145494045281675839165924219030103802598741;
B[66]<=2560'd202206764794965830340576670731060913592530898012384997595854637721978906372155741008905860611891326562185876198699608708893977439210593341345117282028249267554743787855396228451864840130608996421622380648411853673506974561355258387314437386796042842784646910007145879514333480831891088593447677591476827562773786298821183714662891788503947480800499719863354982905790351143572752288230907561961468034155994710153872022485910901519943928120792197753114171035384132527418474661296414131202382469058572679203834952894975000242403093792075411235454725853822607717366889941599497002694274518684448964298399505223893161353863197890821180577404280575734462758741461544379182629484204048884282936058814882682712231455030641042551216038944386057884392714193178287294282674145154133;
B[67]<=2560'd202206764794965830340576670731060913592530898012384997595854637721994978370146327264807275263785789640441805224141483895259364224667125479240919553429889596500854043831630903898058014500483087465359994464079494799123449145754203587058856778721717528106490591896969257097751597986351792216023905669235869634909191014536355128191034422706999549381085235777639063579396600435793526750460935793008934041034163463173727802532746101457428076471497764874080064372413802136431124659725209229656518921844793226189709037447123640689930103794894193383470396976252255250225994027039901911008720432963701590587492960290369894060192363917999789837187130390437449614612911701662666139095107901086818393072843891533771154934143261418081039639305500718781153495523934780546351083017295189;
B[68]<=2560'd202206764794965830340576670731060913592530898012384997595854637721979910626734559901916279644091768637006198086995792373741421417444834333590283242240725929010682485707843218093741606074095455134455834250108112431571276795433196389451551542865660011810048577006888513478972618460192087410254651286866499520415345747683070436986325815631224115299327633773222715677252048549151480270681934627124026147684010295447767378364623413688853520327323954264330487904453822478071501088726142347759281712088924835997087022669742330559512689011218864776631288688052169388783977415492522060558094638696551581177665432432990065098805279417580655208115042292073287839765138601942382285696096566210705648501972447646136306739118081448280548960975363373656627476205102250570652415110174037;
B[69]<=2560'd202206764895851397194244927231153184142646520854802078555218860891441421341334396618649488370822874438669164793392295005024788699370720554325683942788056978349820898136096055716029589901109407724792682618737973007778258695475638297631781236902360225673631772890986781566749070310913774367951500227892492026418447712714863415587953842367487951713883002941209674326162426012112336770794160600681505817381145028733017622124517719463325107104900218448353787998814067730812180959792665001536290543111719315520639718526225255638059048865106802744409288084237116512908064287137068958746193843317991726576404290815791047676923477444735512904311977295459694074749877058302223690979827277953906159562699873030030318402652062998738152657852079306164077413970190119836239975405671764;
B[70]<=2560'd202206764794965830340576670731060913592530898012384997595854655627985802619839562260935171341937229663991544496816260050654688739696126329011252236061622842553891107807120563987035457370746537322086197541545674998088329315751658519690720169920461139072660513618847236033674611231983213799198559915990582278633219682450794053877317242910263147657258320881032670298445864693372260621815908274539177717216558960634352402259213661402570682625252127326508261931594390887107056810059426581977759598476405470150506877860161991123482887182208084053261186866269875324370252302925299754159111155873939775924046838793167587359885347579126642189123012005984759897962585518959637852105197645414247363877812079470453120774771641160644629892026797541025426131717357219150090924396467541;
B[71]<=2560'd202206764794965830364065922196985988822741049198159154150092756144458000176596689666025015955148226635962754718559531934074121838469615693724613709349946388133269805948914810095611413099700030295411951985447935667863957786137383061178307164448082756101720654355074327705859773764625005211181331062864893138736144302005402489077377673485995315752044344990124055283749048976708662501700488355894455378796547503265454981366808997444817294428274440790498591738641286125299475377321873513953105664700722213159898817497734606824844311483359035931637113970793679303304304989650756302421727853149045926736996000397057301022818005199560721035180701003201486994558239583041082794047606442733826038309171067878397988741439555967102743571471083523119700959603928308922468989341619285;
B[72]<=2560'd202206766409134900000736852949157559596268997940169177730321516789285017078057356772879547744522999664338424041156566181750606315378563203174890135855589316169502623942354776470110557124439747029231032841946615177544935417384247159765547409622337786650578184126367666539912491769735608097504232100205440743150441862074065548227775391942665464365841113446420157516581802760573051685759832471599547276263106533858876300647474228150499392908848993791175775679994839592550346756285887203807730699519379283970554984816623452413314380387289288607803315740552518416688847021896505623653061878437530456183780472819338737104181157104294194804765371746382673475033970568552560206282173480510610490566748291532379564063616768736198723248386844127489202545208549812565526705075475797;
B[73]<=2560'd202206764794965830340576670731060913592530898012384997595854637722252134263798912229243451348782273007743352953949952991597205927122738239190780443209914631415371520663885026512818232384731214596912268356844203549601454104840493760690142578705903248975877343219110476383002958128669601217002459327580007554399044847771281909070089652299697884454628119785972284259578382557836844342040921091388330722556529798787014454804556271201582174875708705522073684966124262403566493350903812681116911776731924661709419942092954143496294487745717783764357872891669693965811161776374288637520617616413437409971077681219582099438317025802338249831226849959976730222064280681651633315395058937261049830841197146670673253437050773412786224699320063787817922015403448022980335239509136725;
B[74]<=2560'd202206764794965830340576670731059578383171093584651847395594461016702750544318898403920394065847544434288252144454275005407125911815455186777218800621312801129766795969743310009447397634297796867485895892818419375071845854967012223765671899916582766410164768484734314187881519494650861768808326838641137598777886929124463577911353788133778832283280959450938844854203482353225516980038940154238716764874485921483180919939548630507859024069835907232662419539447884070238099071035387326228097584063533560971544088963008695329515476211271280777846068513308971286621392006261190973929586776212157813027546345060256763047303693671605665555766465466239388783239423337533759884126582309214274437009512440930057748235867568020414801750057738473106893119214751100561510581784630596;
B[75]<=2560'd202206764794965830340576670731060913592530898012384997595854637726367632784312820614950777208689931040768098431370730021813517141137678407427129257416701015567049489594560314940602195357008769499505688877666399956781602239726190182177724978960596776824598294948252383684907746354212328595357336455182983873143707088064259857605198450558665627848730433390436327567374460092388128237625265223048444478623758941202614978535555641397423468272004083276940870778990644566775007826090478788447089352910144511920595850429039890984216489929113870951459911810092491179739589854984821419298934750413541833847079371595589980127817942838661301594038881033954203541958700459720755398789524925332576536753635601669378648313298039524096453534597381573691279433019325533477657349310469461;
B[76]<=2560'd202206764794965830340576670731060913592530896722121294189869816004423232044226069424106195617983435662061550161763143224220827508807754742451471207263673630967657511052127502717626796142721339568677861510901601941809424738919244215865033681322414622243796338765533129999687442865160692289347387842588433199742035457240041980762816154590583170140660463985901787974581616238352054931359944581626323940686630580454730668961101929834655398476529122324784175282637856068708877559381727356790644793750085146586132428366260611431666210941841185573868059489156826896656051896249776399252019108589630159593333612458511118347641263833507561406335862834320951567264358328669647474315456124513304864273859772766176366885811598056994077840161452197155063800169132604223336334744704341;
B[77]<=2560'd202206764794965830342044748947681230794419032385598017474259849268568588290595947563929945307087012941798044703134536723688660720720887558901316893826781357646244489635702713455919197634080780522910084411134053481527985451890952343449652388959139695229065746375247667097025836591603913665993428990325485473301763653901832884671892564221049360743342655774174410482806586224459936749210300766953967252432341982528624108443943227722902716360803373251413130453902095711942768828798212504335868939053147034196353569591573005517599091846530515573117472912411870319969513899035793240441133506283496926039152885678328856093673457609581451380135926747675575963568725171856085880505857580230603114386540954582973812758599783297320133345780554178825590595065010242638931325655274837;
B[78]<=2560'd202206764794965830340576670731060913592530898012384997595854638845491934014285742993883823598941110873652919928175889228139690395345165876462492024844954849986599374493841992265334069287337641133051493811589642337837488755321775295725507969046164759339282438185862760930885139218360625372958346227774978389735729147261443966173478367165206352495444017793718061975529970144491554136660377242291315037044483523859445628983865152080628884787168401090323344814725598233093079568597397364443663921272995621222586239386449578922663679415764646920379508680826070604682951303914085626316855698335697222106686920684515229214046899065688121389534585439422793776153635214772666821943198867399086501183007182616961789608991031893970823791126463864578321356398652415198694072540026197;
B[79]<=2560'd202206764794965830340576670731060913592530898012384997595854637726367633045837232290147021387774268478005619948431922039417856361272436659775403293167635104963370749095715089232749949601042670545470553793861211591909180831063764301770363174378328029794476302067125338780190126096658332790785092952159977162103525012660397794746800403517890843573627633552327613606788925337421748485828940771501141979147225622737574570032665871472173814141648032508154441370369793763241772673963387021908181123986288725752921546609648964172839105539370702430174295708514558470030138135284525441455256740173660959707910904553133673770352528121964540459363378668751307529800725512142890901247581569469814969846881657173290236061368776194931830409274805481805437731296571594270711399979504981;
B[80]<=2560'd202206764794965830342044748947681230794419032461495882663240397374238141333166200706719790326868698720611738576497770095921473829299028031513413006645764871893367863088042429704935927876509725256772224683015953744086483624018218240229256948735736918358525350726093634749105879349689580996615730561013265983968118882800122217030814891178993010049156962528440796376728654965849605731236799163401636189987269175442327764830120518118463557315327093395572056987847487506759620530978933039017791868504568024724032156490737483537627734442145763447259713069972647288251239363324506669653778365535098671857889127229607876920281208440920899008399210680076333257567087534312240429566899362141553633206124846264860428264473369864138045089097321223586946457586211369352727283142772053;
B[81]<=2560'd202206764794965830340576670731060913592530898012384997595854637792198537045190312773154113844896053552007135093365975377327305546189331985775914560053431020455283826852136288516408162972912611055874047011630931259749371162108174465313306023878024121872785284031448883748488676811528153996904984212265859677314945461342700136970364048556581943504526807680477155005047329215258780503459700744403536108741537826235089013875886949707797692222885679785536472316164746859810040947828952011517481886073898611450872581718196224345959708189091408260820053407752203538463837426561328195285892225407998195469255661158906449469101911235961556416445597419697561086433912828263111807936480483727488962079486494112696615030940519353320390568239718954750513158588954476782362095351256405;
B[82]<=2560'd202206764794965830340576670731060913592530898012384997595854655698204428793055853188952968160732771098970021185552956260785102791074728162302233348022058440095128124815143729094862814421376585025085429969764960695283908956631255436595842814162110989788929275920096320359742872375009745318814186560834563940435473962280241370857649443934021647612981697690013974304637164934429330275235045804674926086082143669930657060046354774707008170795037613324934091456490540338310595515453500595993482376127998160652319877602222400136620992154317832219603686973267667136796017821253829238512320601912761390539705665102167141328334178522526146286774284589905013044094857421495268324879424636282155326277891278142200041607587525172909723089809978090455636699267199215931814261393015893;
B[83]<=2560'd202206764794965830340576670731060913592530898012384997595854655698204429053622533007888865662261863778393165313169068052940333381531757860547800474117381209402874357779698554152906462961803491885427853569176016013549535480590632106444907097106125243495314448308765692597680238742245510081167393944664735515892733155303069910672330991777563751065265087311411178005199394506523132768988450622134695256417300239643484676217558298075031569197991131107678463863328994082734779579754029332584006124347797660187670227778029390992115698299389397205547907534133859832729661348510788516840089770480265926665602799324871936752372506631226798210182159517324252700321711177587423215901945617821342000804780714059912009837531588591184691454269955710642972290536359925170371312452195413;
B[84]<=2560'd202206764794965830340576670731060913592530897936487132972361815196491881199985789068025924443017771143103056843417760489205605538637468709623776308902875697069172294899932349868970704689995300187659476920293278382979681672191791229529583459381802211347104778435534355456552437516439892919669350396994934250507920952360107217577969498662461184305435250741050502041072570407947158239490524830467848106324245122420932024157139904765945277288740759706193616593354917873969327401993706385220171401314900825109141105497333337113114212775999778391787625386809618405130793309059199567925346076731200838117246427474121553494951659057523894070065087979565237774269009681104684601921449968561635066522569428718383632560324665460766306103643075923719445671816084440319986484087444548;
B[85]<=2560'd202206764794965830340576670731060913592530898012384997878600801468929541625792308152201288971991041343696397082731022670453743661721557474623393080403659845950761162119162933770507756404435756517923682707053922838257168290093584969126610704753826025165383803420836475416974893197693502366481616117231893486686599147088882958949204751889377565897540305768822254610849962412071499723595447801851602236633372337228309835763999574126579370700137680681078620199303924739842993551719704787005944051171385116376824483058886586909478343198903972064014560730731982934010730846688510634685650027599669845868299186169614150635365711745306553559509102945854899342575211468175934385608214656690316067465251977396241585288436349719348571499958527254582810878057802070985950949077767253;
B[86]<=2560'd202206764794965830340576670731060913592530898012384997595859221659761551779740181583586004108030895607377326779628517216311277106303548711148683231463376492351956102776698963585098283273700317748336446589545448775108312060181745422311428718143816213407922610998283152184914323751334311407109193042307105663891788773393194139001140862088800946465505094440256785988654784053702723022257901510535737765500010623674504938122155222066093672047933858241676983769932263242576416285299589393010971866404081737628915835628545620020793475966479724901531275074012052769392387433873883566486750822535186112290529297194607431067374843927465636880942987514253494521489461674825387027900437845433622439717662251720108197185048105993764167146828516332242715138470145324313949408769360981;
B[87]<=2560'd202206764794965830340576670731060913592530898088282862502162670676648178133443753462056840007227527426644919510674020699198870664914689047836204272473376120800888626465439576212486150279535065103293440355836600010503913938543348549681195122319043883970125373493289453377764997385780734165516053045621091304917292867022012242470490478874061704876871538270154809183301421821197428343975833287667111486919811621706045109781509603754288515315042223176932595356684196427891556536888670203479226400096275241516817877476385847985709018508158597354703048294089569771275296918101645701245100613878144152154055335592058907903910167131137418033443797493007054470789995902336817360380328319208013505110540712369908188466654469960450145656724308028643907279411916112459345216337626197;
B[88]<=2560'd202206764801271178268930936762316680501913105010182726066691368544398003195479530109402487350825684630660239371341385180504179611787483282523056614502123027619720247932146980586007747923718765191111821137203599005543491778306096798423165773893477337173848176261807441799334141584922186629784460976109990923129348547035759139886366675383707884949739100749460081772705465501090728218069681781364638585831806017306197985299861723366611806499790064721487182372391733705242282986998283537249397618436413436247264201390001089548311586937412314297262429349874030722101228556615438964052654108079472821861254114477294640889938257066047170090916685694276974248589129076729018723673603593104465913931070144972085630582321714798144677241013596380147624911198604398099217844759970884;
B[89]<=2560'd202206764794965830340576670731060913592530898012385069978872826584450213428629785370814497431690131340677385492186005028396450865621262608296182911718893481778656433722860693240620575980811605541969278264872839383959189251741328634687347518084482858822189205580774886880851405212591437157909263494370239858756124835905244547047431467144893712234317520125368721068191878721973287128615160971639094014410455341864953156798761041731362647907023117957927852386580453365100877063801391561910118034987184684108453798482913081676047785193863035285442650477296170053949546084291361837265302556209286640976667466781136558592785042685053953898001801809764465135302531056515259715407689342984630567488899782859327514246142714529349835977196566755550317512221633782204452564949550148;
B[90]<=2560'd202206764794965830340576670731060830141945910235651675708407422306564074021230163750085512775189196217252258494722770552093038679978375356664724411529381032865940742001969673098025689740193363736172428825756537044154948370635186637685423765521410925841714473850975463890855336999074571090335847641779777676808391766912301446319076848589525218145941648850658612217907761169973903396741656922099346512179414948648960895116580392397326254657273870028687606086084807502430027768092621749500679952827180659950964283138705874270071025295774225873249421693984308623060342199726091433822923873417714951787582510090023538776191573975879043280764164410747614363178579591354469717970898953088199500168126423016425729950375267850139708104974112148717815707859064839760146746756580420;
B[91]<=2560'd202206764794965830340576670725591896054771962017698253347358797513110318207619419555246234318052091438749856916171836955275211391138086725260615799568793540272687091911854108980143551768175169709590341027420801522925245078553261118595040305882763665716184456483753176108828549657457568607187346422962877129086257348228579551203347706735557072525468862572371012916411569244540324305510825257868966439021367629653922212425917711433129298842553795813862974037065316425021654249097666179509892872714970646146373135990888944996151122459329437568978345340309441831743928981646417702635459437006229177122353285305529652783868193281161936351370990889976283890229867186895715811901031977927579200023329011528533650403431261399161489801301378825287008955847835368386154094692484165;
B[92]<=2560'd202206764794965830339016479208026658399785454440490222142601687528058808453330635950368559662037469210342469952859116835506284878333488997445368663403439173625857639071419154684632338333011226537077498856338182964362303021756003381451572574531042169631934232095190277030513865002918812411049126881832634769992353924451058421874367855507756642743805782022050762102328282748371017566044822957332292865037350543032610622093233218796283833497150659231857475613769769519971741160481355346774372762325631796246155019035969561025086708813070357906382251890452139583921598829673154804436441109860113785283664467530640039246112676050000657955249600617346944390658282356692478392956343168992366875536054836484835064605237582215570598394255912522489666432889718318239587998538941525;
B[93]<=2560'd202206764794965830339016479208368471995895389154246035875271842669561675979679488525283689050874782466219875419232693353452676814611056480659852182768864090696909280891965779335848677306281415999452887309832303128682126101392944356898958692566797113318181257706981688913757874381709186635250654479370703529252423966968159140169273291830042606662609954860235130130535701497575309154518487281678776562119224492992634089774778400333930080161964754703387769597393352220422419749535182939323153980371810381320294598459282703016984990348460565329851510292263746554467675934062848607412300364398518395528166374759278405252953958371800535088814877630945790565104243831144921455623863687592341709564044285657547516992720573823630239481362192300418209711316847408305071014165103701;
B[94]<=2560'd202206764794965830340576289906962706824540759345807011553145211095224259209581517301470426085182507919217441008976879517304841328486843877801125495319024532948352774842583333754280696995584213549246737519049697864041973669861460279934945519795010299105008931598863239710947181867857744509549748361473086484569719591039565725511741887909028695429942038410171826237432392210927692086881238642287438467797621675747180707997237958025854526301636781077477837331748013713326519801216229542614292142144651608600876501307473710571653243744515953440063445779256091857975812952272928433370607755750346561127755476896802020422416093408070007240323511874635444623463096918157810084115962403216156306434166136178588467591065273746232132998933508293080736000550151540317573218904065109;
B[95]<=2560'd203899343741352263072221764351008270114544360126718504178865927068436273559235142245842278714728663140811036145239240287713803579078041342365570022727114574085588796085513999587257153002094976851606412643975974664283753382162980501145578349761069623871941513166309218480655311986944721441953254545691334132463868207098736200797304161844734126011868268899167301430988443551650187916472126258071535154201092490103141346507579563847603929607191644525633307894873083925881000016154412953935068809585340338566482466378722851904955251096241666393129645237169937744168508018059973619856247356329570589478564440217439898112557449768553455429015789185371275118058221841212546888892024628480398395899600115301975569620205348970112864652706152288444977662403786286790927225922536517;
B[96]<=2560'd202206764902130575465669988539525048080671537370330085879916097088269475521809930605250559632088705953930462963837193302357157471924500725711846602266508794480311536234004314500492047320376562061260557833789702991114465513244072790922065787545724500530921891832686534793360738457744468818937939643667519165173895318170997912068676503254196662789029994787620288463071752119037121133351278863530191412402323320500172782291602193229239291750966632844673129749931855553923722709037885336446400827968386478031202671565266084109825509759071482274946502166139739991356840826300126661843977814170177091445084780194288772824854281654423931944456409616753583911046672260755796038102587830854360113115320407239933012168683675139425821939949674990377648188387348928988413240935728196;
B[97]<=2560'd202206764794939564471673461584537890759793757078698644247341000957097508367962944319064029299203453146888311419372215503952844645316541222026074219827012885081059603405766158870581824154233311454678917117446591304245587356159585718265306222134753116040907850565695558581202193725437057920899855867509440466299638753168672297091490914165379752626534739612000127917427998279637398590756547008460090380015070609636894649182015403463308529031770700062440624739085894667067988778327375488687794541250999336116643958529717259818105941580152184505526995441154244912277251202288063867253769089590084258540924059690874387693275479285333933202031218102772407191789632347122249783325771547190992950937161788043139267588550601041569779681074851564075787757734066559124739284760020036;
B[98]<=2560'd202206764794965830340576670731060913592530898012384997595854655627984798120915398368914754059672542473744149221693957551767302839864577607833536788818574816965839387167301586597938325230579037692354095786206011033353561952696509672303846310745681846050141218965206493273912993822028983194186555884693879090800604762661898787785876157992165104427582930357461203134698473216445905341442579042739468016099309129683806460426459316195539828519697690679735822151951609536370228020507533378900939817060538966189884691004726062839702929547721005850699552703049822489313121489285233663575719067721927077059492014551144016270339894333319143229995612766807080844745050593532238131166287106438382052485238108573394631991587159916945073057802318229890042040560822656772542946808710212;
B[99]<=2560'd202199739931174675712540056306077967941486419826974267524295755979782113472810276544349651623582024024389181838621985849164315662585394003875553537854797876059452404313972673356813803710685407044629450749202143551140953949485657162345536673458971073368124930704732912953820791390265320640317419400913151724435589319863580941190238760512171888063472519605678206765134912289413136209839765753986578517463183200012667606465467042334346451985959557703821317774928447324296372611794029495816152214779819510055784538321718192560827195425146598777044736669066691012870060683506661878340644593178473246832047960890670926270186625700482907396343421837879249977316434524024825339577645445895498437680120160264876538941608430683449761928050198206566415031472124346295117036262802500;
B[100]<=2560'd202199739931174675712540056306077967941486419746332786080197510479828886251506830040526317467541238089454557133634960923331958848785975402087783780610534247542886236866993421673027416386309254063077926771884591143770308191455050854157725479749314591865925641748941978606499572361004048762419915692435423131200383019082038577804667114739702958649789682067144289779769554671692751370413817660182355541137844561197050760833154926662187118837097323509309954589897420020247113655444864325262932743448115432475820000177346196279744642936251442516048032698696922227846571970023815467298758940760109078674345774185334214659333989193496758960720397556562602504988768415400755205604687809869030477638761387231723404210968688070424986952453190405416531150021167762049092987572732996;
B[101]<=2560'd175125501652782906634249438043865255522107626785343644700119907208430641369966504948532731022855657542688312717140404161575249566483868244511417282323034242844312799407921441442351256483835966830757441210239248785379278567890066690038908453050651602538293920893389661233745470611360893901558852543223074953106020752180902944740285714911038952814517637273811390226596516131372225489434211502097361033156241123324599728406175864011039065691358128266977779619212756982025076750857882109473569399724465259685633616703589267596530246600715595051514895338308002059551777231472976885275296126652936334391078695630623981849551938144760634881602909980665334024577946772954825858246592365134033747459699051496577423242122516565320738608575234271021254450252728428875223421306618948;
B[102]<=2560'd202206764794965830340576670731060913592530917442238413610637443497844801359684540215483627553652845517043624649839008395154394273246671942269912695857391818587623945308127898773125246357098525102613562482910956543505538790812567559089530175651631780406437486130054937818602164469708830489809756033715047400617523256792397036448438471087799365000995741980704407285172704694463678529486151417538660915985841410961387514174477335777716236879080269130762667595102842375185870039854852752538222781956972758187366576260228755807371989511684145121611107677926805278454054406682309378120057048425580657748188028293908008777058273257005824812318797688609835703584717947454667936382713765225056758453006196805783960977018013400873089152850656536713271890917355968948972322180842564;
B[103]<=2560'd202206764788660476398974029422644074153240366049033787368730864220654613847216434482823260611575771796182070809092122032312918948013597162711700715414819892588296203415592039814367397457480263287174859670390777920190982704556749769293974430440915256727887346249302329205495452802887045778427742633608183197170645084245926954977243981291963986749973290624984933977030517494129321040547827678299590576052686510787214707342634667001421521834378411118612498816671298688154294439471148570056935854865275034732428283735678855148316973678921958606239047723444894997633021699197208085486566564082200506343258831258306233362312034417031663227364255075545277210833651704904133404675777958035650898244060720305427259999892000996893527312678197650580833181081235358730459603284542532;
B[104]<=2560'd202206764794939660683647466013646033700573012795278047364282823522244966119141856923032498465193704699800913241733543053481870619535907662523072646853065825567596734511220692078595445487949394048398958682984071541986737829900180665249623673538445274003049912167742627209496455028641026619397922676890163663336268753278177917496536296515900426632575498837030656341933315464470848299174319384737461559367739146169726704201614155252287880825116983996131018340811209274217003219864473829463375895754110208735887063288955839670298516195063499422038231322125099645589773003989486722202338470809812821344052266295419724547774739777651126185689183837896251922035523071678125733939021283596195216120432957729056233737262802275621481866133844565264023211838197594142117829105960004;
B[105]<=2560'd202206764794965830340576670731060913614257515540979060588785616053402267156764594366870351912319402093463128333234556962720344142346608205233058974317650422503794430372832060886989962813391971714973859139451229070581096197048399597740182836709623386214464272722832389032406601269497884471481152405593896848048169749255255876934318490669158450006701229195172356541184613614273930381525879333434943615359536407970568702255865223869901796468553095572834187188979566157894957377054275875928870585712727784715360108525012001934035115361669088606174488716874269458936085123352416087627693924267957291081623256106092779935383018158160211413604432249680946252223607353886946697723790932524088155607822735470596818681550525979986249358715633369469975662027428446860918544450995268;
B[106]<=2560'd202206764794965830340576670731060913592610482691976917240517388624189772780638517362897100563845810483779150960035245292650159065318203698532369005930498524339653585970367381843400871589553653355259772763129872951785559190069895719075038720775549186498193910072490263815406234776491468675482021658265209216306489266061003296092472313842628480214947686017767472960833938193132556280008901408660991788367349501021981352444948278178905843256252253942230890629417000928627708449885945780395283986175509324696852863866176344391175613209202520410365176560982836674899757978144410139864272683278372217442860710232212462118237283061632982049711236980214560748551618140801558637742845062554968197187980214482054578741099211455619491508253167431899929282310651332121563798039708740;
B[107]<=2560'd202206764794965830340484915842522143767413221131189477728684063063878826320874941562260425074083700142981326533581392082888843874010923008457328817716963607242766776267970011202373341107310564060296907113871883410293428616051950105042093218849495184856531658558203243891131085198251417008836993927686201525171155341455996927430431057669268764063704784739988796688321989182278078499838890598942665995057758215797761814429080337764573388989162398961620352831770525221979078147322244720064641390663159389775182739102037362059975665851012647945262347868375335049932295903590109361590572185257125720076445921419562274291216503287127747800376944448494372678477988708025595056713104398299424153937189752572270616066751630668161996123132020535716655399625518736329672744096777284;
B[108]<=2560'd202206764794965830340576670736188117535453276025371735421865823450585829665443754361464027045777998716415728395250713974030539064396598163478362147480860475792964911251595735664444911317857889134643316312256769061147357468458240704910474362684871001217791938533634407233770110571649804322727108694340620193072354676825428352549267868086277397666054788908225164239252404232148484876909076765678296246798195330071045717362639790841948455420074520820079016349133477111328033117339483895925786706071515918047467200251283775770171139602034659623190609212834478523108340369937215137681268626056807031801006625973611712055999295199371686700496686653413025535965066230194885966151536059378986393146927178787342018463104681698303490291063896182510780017389878659260919692059231300;
B[109]<=2560'd202206764788660482412222404704933769286095405837559805098592183491809490189028236701848300896126836671669747348638254727931379379872464655788261237051560332057101812643292840366609746078085052944208712731879805017179095504636583684604682109617499829526585115094989145330616559977091550977659334126656800393715644173226458854616894950351025286478688511265204206675212130802553379676914035182442404260404498322573963967342127906832315951733404926613420117781015588167886801570657050544007832141592976829066989421997887870436509705109817229841072733901189272997430505041253924308895415229681172035995803280745937231477278350982810927875688496577291263466065891598735463661982920863891572561200766932647057788682664852743309497496385780657593813632452248327588570870352987204;
B[110]<=2560'd202206764794965830340576670731060913592615767612402544189211038986557324464889377499643471155655223985232345405834233866276738073264782901724452957440954182476432989623489570383859280695827288233405912566611018362131713440679944327167689499450363155007219980173886742440974039346572044291462742451373942755343866134641538664640798698810191909530947442691225269896843849103533945156120716486725945881587159149142682854125518053392159054882093860895436838035025642565157630917114391073891681944193059147558821172277890863129566896318759202229487068025647589981077609390215220347111939004490453438613031217215152893931624769572669337958845787466815511984985040111176989809967942859680204728297378521199598756859484095590617322142376001507173877087837196953812600645218485316;
B[111]<=2560'd202206764794965830340576670731060913614262821181225330904680839282458587896329593061362364304126094005050455586261423677979979942372363929931768625765591074334895770175248388713913963837812734854579936018049553826710393194811978799651334138457926069751336862351071255708973795694079711419927314223683463168721673227881223109404562857200982267566519827301315416465715639464267114373995460847344055116414007019757268707930930678948887973778518266870592286659148108166029968697211479529637142463147863895878678583282213210659691679731042475443780035471351010060215668122245313699594191292878524171782460088263846582862069614260329274275298435380433253173993374279135166474567543622631820163721362747107817107210646826637448505964713457907232523714823541292557636711506789444;
B[112]<=2560'd202206764794965824327328295454583473818134855148208843861417797286039665294172956497470163624253976182937086736170997724216245079745241468367143941087693861997037985959805045191221641319321699826943139889442799751882024922370192648791405741207176436970659609728142450215619080271622860746895719991276440569646106068465328047374227893651979952908154813102535604543512764647150002964191314870034883310323987150883504142282568172979796132138344857655113819856164627632577773903466594156095992637149910941703493218099972059923837641737216667047876395110598387085480309303470193121710774722268543421605799235288972360130159086623365638898578163513757736212900975906711481761670905629875988626896700188076775251033082914774400452068580001633878666496660353461290470617244779588;
B[113]<=2560'd202206764794965830340576670731060913614262801756115531465313222043362502268480838274623210820961801949630154334846564959949802259666540341430978887394902253512480789749306407446708515324497231098282774448437246375091916194765915222544825080273447146178834598522439327434537804041744488484155331744000389778798953549925237395271153676413486214859919656919172423663325255478202802368938056789714346527014650577078117527729185927182153398637077820494089264284772475170869592096341845287105878985551842986944011243335236401463204702545088351658818157053662240868148029975260681107419525548107708175672415702785434263256499720512739426472587583101711985966424506379156145103539778943020863596682070008537479378132065583395720784560019636210086461280815107135541361456581985348;
B[114]<=2560'd202206764794965830317087419265137257023623453916878145472449734705315829271463294912353371407709098253557324416111136614802362516891564747503310106380026464605561562783584477910891413449411096850628447188172431805128200193918419537911541290721185100025187954521835307083652006022884100497874357457913173517355758699122240535458617232817423443992056362552960412720230685800952137610036353426551896367630076347842676894765340516279548575104826485375240806583938897052359737508206152711667562067436731501269858654839296094506383254072760758698362984335642137797287541505255375367215704210147083782931927095094684991870150758167710466658206861772382995542710204683853172018644775971715763742949389830218261324953705663478271950949772203286931373095845937556860102682192659524;
B[115]<=2560'd202206764794965830317087419265137257043992177279788495524329255051020186749320974312857088352281870541030914749533913272767171387019936590028576953390253970500522294718050430972382633384675105674708701734946433362749975320419115307805729027202033296871546715598356093686908838955208964868884285642640213087401763727581629660712699557749806162346413650648247974841769706926981310104193459105005421053647981631482628436128596870071243640538238193103919247988127135806874781563267676161113406678281100932361340162787645483888317424572845470531110412699529702804217613135551071471865102442410072541018356594246397729969876197353283500029203046175571840351188354415407971876705531893057357847942480519965360634016455365357564314157008411667907610789137732102737654904942511172;
B[116]<=2560'd231086393067684338824277196213890658679329704966183045558806936150022843396048172425392151143559047750400996672090792883321346378304879083076228629869227568261068147231016615363257653640316748966648145532918157840582866426730107987793221248582280667436439824589944731744128789907964944018909298529171302664767531412945173610183636350908175991268884877674891155994910320132590470982648911057121507233770517720135228460938594988542922957040671403087896859539334595352471770025626542200230961276138372830309981161947474284469667496730548809890616684480590778504157928050187582706928328966236950279782904076913688672574345000188516717422212596268017383488015478016565830230143551734536112308084119174651557395226989331750732218967914881754662871476497442892334076257003390021;
B[117]<=2560'd229288028038034320900572159918712024722313901691156584013686590980392806895628196861397220743475981022301422325356159372278078513497889796242965915366842163740115020242966835178470980962309380422210646242891659756648273733705121615469597676403496700741300541747029775984086828673738541468957232588599655312815498357775141119837083042342902951713986247798447043653933354170332172789381181327519730053652661736354620409134132498898372975811197611601229612676578610759191050719779254331805040294094943541721703309778036171163693164180753537044328600356246855652637442719543187559410795378743627139615468441719450397632166527040576446234895015178130357765820317106031046097093628433965867131418108344861754524568320879517697467820049498215659532656849096874782596740700980292;
B[118]<=2560'd202206766510020466852937031232994114113680415319146342058743371660349955918399213733006719379526936955853404695512845237806607831299570315569672819916137334316312674200571582610573441880236400140824948171267818719228425160350476453409487454746236477271539571975464541695440623963317444516885116369999499838623315507966540528685076421730883833384080682354284840922762166175134857006327050614846348193429839190356255837694535229772425987481951073182760962030194781202937227736853221560968307984678867837120126210830583379941307724941204855785940956162156633582421784981953005714281198256032996811369997869405565742814173000004295436809411093438162388121804338630115493239826840922144602011765442567216543165340430287270607363687873147551300420298747822600415710602932274244;
B[119]<=2560'd202319162616043018900035513183366184372176188285575388987605479389755792348615697396260602049074580871240226282378716853102453661742596058542582573610284961758306756140153809811505644117713639538337779334878449298805872771553347066254308879285800580128495332218245549847593436553345574893015987127177039540646339211273525760984827778950201891192745683763903318766371573123571608169962371709899669906609079970157622802590339594094189212692102102084577145643225578926072042459343968752376058173602416247237295072098666868200710482626301005233568466983844906027720186015048771566196958743514841859005194058151790352073076714836915917536696674093310367399522625595387292896681499589193554515363222059282337459879026301672002591591761547798057471126362152362414344530714444868;
B[120]<=2560'd202206766510020466876426282791892487485872063175143557733085721258593969019847109956077072555407729876722627378878710693315807591124462253073512891979647950788780181582879940422416556735904868851894263882506791857182017192608347983657514642995987776415026732362856693368844715138152926618335607845357987927541090772384527810373368058992445889758069998946707696034841582520250397297348425043257968546016498016771824166423568255130738581589241334253470325454963064584315972038435651552634480771248297244230822895875828511713290743100371737682769244224312241679209859180186500335957826247599844111428445208112806791378494393694289190098364858536425223626370308307590786167001984967782882849506742308120284897646228264183023358598379301303856915134050902703358904026750272580;
B[121]<=2560'd231086394782738975338197389826451963417613115178895993555052266922179401634466028608874508236513314155117172951486386023759971165587087349455480542164770533668901741906368945371729115291198588651544590082383152331612615300088785342137715602326766842734887891274304239668160982166643357898103022721483709939444449134416281086228700353753130794189228189534360676013877483264210241398716295739299425914479173615750669601128782795164508676085525012278439606617448744443962684166579859738797530717002486993098008015894555934711664851194624589029551053372068209584140824983245757098187303740017323946923804606042290975097000147786052686430242196326840409580661256463573371482175623103333873388101177541740597529249232215452122602292750890871587740495043029520566675925161493572;
B[122]<=2560'd231086393175295507510310898288104047779141058704535216436222878583140824010026811446391847355864126111033640517762922009755861481273174725269307896857799760231463757241917129603032548838731364593424640435965794312852529133911001331925441539707206621101639949288889049626503701739113830645739743934116264808769118988601667678724258294030680759598023540862697366913370903794674167558753903538819353313197955414462747145530701106606572575917768509835183215986028415079819168628943886856379732164037644509834171856174315294309743201743102402080655811183118297884743962614584030382219527018989899761063054833227995414692442043130803760896786253758952365130725364484744919795701046350720441573386584895716722318339028325850197852358469648789278091693996190532613925829364433988;
B[123]<=2560'd202319575950517408323360766403667552522472544017166111354454291289442527168463126335066849368055958269920479223561568874525718932727001604708446819578002545987936846410704862202404467069976760487048827341424846639331610401964488468232232078757593703623890014111693238849119827022921546104259473315249817523825493764970224033237075015397194879836150173859977321956021725016532844414450084630664049682472817368783935998204754298947594379679965715629373212175968591371224690613633899742239098100738798252764449949048685957971187252666102610139885741688969949220321595609531229071964307946523910685817829148215318912405249176354556662634385908116754962408790546435845145120812713604705553652883054832333578804470796628487684539309258682238712289620983568947261595328721470532;
B[124]<=2560'd204012182337778025254331819483900659668427953421422443043757911105776322406571123387326258878299337136898582329861796625770056436684855117243489143165986553135209290247355600072261023504311670476446608978137281609289482276996819301936276544713843150470332007819304110493423613153184525655284886195171212663937968525122467407021810138351019499731585844897850449626738184033429792095990778887931778344675464243880036475082254501913266137813214375482375389884056227205855480399525075981196363363147088858446588482190116248203833155716796745052800713339447179549789972996526313626403747739389736346908421859504446093226268469276757478881549711390545131049529470835823051272383654963690752839967350661672997274912172383443455942277154161690757207024677518193988528806692144196;
B[125]<=2560'd231093445479960948960659052264069615880753136563475016810091384945074129662697942470485194130403685528927679711826238416191460782623660492179434630645152334038503527639494624991376154131685710409122233915826862476893753057375073097415782086816092357933591280256992913827923125032797824279949685254219723707774839895151792120159003887368023107310581656274813317056485671403754381908178573158600454174091460191021579564843225657930360489016009157094235310206659115906934217694442629573601036669628131900449560261370572116386366610762079820195397671647358585742806266801825492047742719929616620594477137747130407943910235874548702504993897142514423737164295626702551637163270490720645458929533411633387165478136304727516670339767566074328203709899044869421308495722522625092;
B[126]<=2560'd231093445479960948960659052264411434692524651229060716709448940866424040803493380939371417673893569642127142228954286174467607344434464665205102779488619397475185137728170416814715613210279604075383662419193031680845027917722604478967564776028604578938215903539546969229000702920105982380856586821082817185019435102519842274333504444417835331881607301236057090726006697745889014667182304723146661001518183326583194357462063569900958190250649196298986287861323046433782981442821532069447472109187034207366435314359906270912192977501083572820911742635454512132470992580349284617135589945927561823374369823560223363891046388013341089170520365973872462940079882514207878252396281712856143493264450262121659712950606488130002385914397551785581036743048389203709585899525522500;
B[127]<=2560'd231093445479960948960659052258942416808418474569875877734098229817627350825640948460940348124831669638473860314303829260606340092757759494983414345379631084928415382536254288055303113457892003178479053759285609448831022174069540938262598391751486957553197199142909752553748589121249306250484961180878438934967700222637491210717301935330866087054684936243356416719324352537869517264390763379841158594959397996297162303557053895561606409737318604556639363727884780089066157838638997674181057864698645446378411669658572715738169862964575817636272271559553505052942594794059884691991129770562083029443944090981407480676180242486796234189800840463585684249112191775887440229732978620946058142313789887684125813567181555090538700668513154788458674634132388225851130008509367364;
B[128]<=2560'd258174708622143872668454363261200791536959537583456522181027942787084062188777254891896497535669429113574804430638266301748606041029172437542453989302472389385018581237579841565641807414206625599047023816234554551850020354996964747005258918829067461398507936536662490023688288666449946908170498955908422997898937894820760932671422790019293594542837528233130665218520548006179370234696006448891831064567283571008344703035410342208332446936582814021346267417246324426481769965110285703707311922951884611834976980323075923444603977280236052130534080501408490912704457548225689921301102820756582520946683988622027264607556683762240195117032481018835125067982512818517174224539287334525464805213467379321970048171179686288447596013759671269003110309737628730359997547849991236;
B[129]<=2560'd231100496177182922584674811638740000307407044082658022540316033277909814932133586013201142388306546002740699750864097460324611406771946055022092718860270262980351184090252131481702266129369676704094084066383981078635495694310896806094537318243106965099677083674384346341700849197818185086914756375931764587484745319744240028230889177207684692749717818392555542649310457902438047260025932319844080847981210935941993530409503784735773454185227748063323555999422082295803311129022166254193137486842835398268098335146382977290756297709933865393462605556583911361781743311054186645462302803554748305597630182336854125703226599827855520750033165986420944726514794371495445301162441051842493917919648687187453567682243889486800358266405342440279295976630572160392742846576477252;
B[130]<=2560'd231206284076386711141203181275407976151574390504770143562668098936577289361837003245375866856386120392244208567815469272660499607696027360741564100323172462785259153711387178163990171094867719521735829324390140664880856901378435846017490262284928470551105892270669838941037590705608031900709521272512555315705085831950304551258786156094745024858596794299762765588365902317069185860955294087301808437748985143932237210346349225314841830202460819889159754324664746707582116159242489245456317812076629256950373105479641001811763070267140797158360521508925126838892147923826322604969572157630863054912232480015799321017990722291597252219120502028266186166905646888221479767280819750563053206213144126325612028012120185569921339092063154523834853201495163161211064672676234308;
B[131]<=2560'd259980126164956067579175866011385552119373573178312884776618091139451296512242817726436728471695424265072914316600719448958874793868186053452550786616474891670712628460096205628211107755225906018475468323998677113658584896160384973028343336722418238927874135834085708351907535744285251262006847703999532921130130343252810132272047810234915516898863203648898876848134105604284696276300864815125976391580717318570039981545746570557733390869555680483368568602134745785125864863908758962667464894134129354831692033494289199107847495717886214660478503040455938917347690849715162134313884471440059563644272625831545043611057275881526951610167483149007704918167242774470523886094279266200859713621338014228023583106783271360770653188176054395377560438312211957129605955017000004;
B[132]<=2560'd259980100439136519895336026273207424934186286741139678349359620902005624919491385028715332418332110428036705276030615589236880796143422724291280152749927952995816419986343113697100440502767672870875297301586608699747077627601077246680085787532845849612814723122959106448243551077603975878705034932828164417860574896529171059319187563409289952178295382373457413668666842557610312904557810575001880125276802038472607648022041737465088162321504787680359044887062801405505560648275416149128185711778218707123318508831284273723655479114363028637521330547205521204596432872927097363204872981431428032521712076063685119196358618328413317283584534851995939467282818062395900874743897116925151102109207856172534435052981891695610368527823962428014564513041617177770917815895999556;
B[133]<=2560'd261785103039585973388517356996529198139529199916141566720812637190013834239014287562690534827351607798468015391591748693935495686741702611586544057786700363014373082513202375005516824038263877858097653748333141882540106437108793592095832626603053652323330433688925904141660137781597314166353632374823381753404520374900969926521536131761554503112738478835631339003072468153569018783362168042882265274668246373616093946280622383062749721903997158729605827396869618225635903384121114940144842580447561419512324565164743345633388678772356076755029319150969306464640441072473781912202516565017229579901311282602325253311175426580254539484737899956707485517717487093444226497446965860713942109055652214283360510435484026662425052030110261747138887348772312720685352232899855428;
B[134]<=2560'd261785517874337443498511679118168114465612038118963650705002689526320897010525254100433615721794965737272311649783359369079278377276930820110919393440690313026138279757837597726197435348021742140873712940214145214526831334733959129713154026366480015759128496981690123919970739828825872323449365020318776147323588823933818931591003225609846833925652073575664906966063300744358415788835284046089498579139974776746984515982044633607360207297302963626000425229222564757416396312864473514810897597270712627982530439796029994878229501793106047113036256044486977523463429481214706366150645396645881403705050015740721236197798184003123638801093798433504956576394168701567855553498203610082341958336519842083335677920460043491770515482173090730664327648769150819166466952399176772;
B[135]<=2560'd259980127880431060621652628369359032429184194769396325124805854537805047158525742161268043990474207438424179095789668820797559275100495404124439456497279663276563131308818517652900640309137904779085723407887910730615607091900577197216750809154727300777992983928277310197556715905926695743028946305245358516213725977182842236995760256675526791982469041886205171966021304853017263805591312806169112247143816266205580006983727595856241854417252116610788563927177616554120292127165216573170507730401474728592455243361575433434646952452965568519614746322807201025694785255058975955514512592784163717816957532840231229773929030743205689909521526567352075549575671997502566312551355082231731592412440601860570137397741143404557996792823935361553188891702747577788562779060585540;
B[136]<=2560'd287061416855204096657401432588891892790243330480824807083203673050849225369293592001423585544542623815338529400230919827664842558358386970398614298899225494128541858572619275779908718084752670429645444714210786753128820536411863750685724216052835914764325328734610369110249066075022435339232156789064585820663550933990281724829299335069404305864011072637079587791885770993143997071033956340511875478536685894576872041010593001290308828669940981647699084781558375198616551569802356992122164416907739519169484924728787437660923654236543804569720856476800884574822870160370386764711689859978202455854637466571096487683268903654081487181072419197943990781129013862625544107926630827065455633677125648685923574634960464131632362089952174270790432224868889944380717583527330884;
B[137]<=2560'd287068441618530028157216591942312906255340128845130840377365442162651510817281739877147384422907943298762522336640392676580213942949859830521149215016010755404260927681212118795854241522830648172067463787757459788305762665574244168219010668222375143164529039549210756463387767823566012780219950725972290377183786230498887445328751112713672768823491537316268506547436609311060019222935082092861206649183151889784136310608339893013562601876280174213037131592843011925834658968190998216480586081956596372420201990126373485040056925636898503758458061502035549641740430999585406168334649062422609900068025014505011712397647216908973800730057692396352381880176342606880294286028348126065316881313057197151114326746186520330431369105210833936971667032162473347295818004562199620;
B[138]<=2560'd259987178476347110861986931236063832181504812519506235015580238160866353878942202988207514032108519531411116948017913631132596389304902931689384196047002435766404908506551845786953555457418097569805117438874423373264730440353847568124171896913363287614458290056873492367070435743460629224059724063687444223280345908999629870243780912906777147460089343964010082508555256023929150089477835892067205375843038111867423419932345758573545435991904924943917227449451406471149720613537298198565492409013485586408105579212805826906617885957799764473437645642382181362414207235552197397180905071201140444991153506766690826127384728831941685992278722104044107778789205253378556323370199956516518755859575141032109529122187901826581563776568224719993496577905278919039913970907759684;
B[139]<=2560'd259980153612161872011917428050462774049506365558621064423128853801869253523363350297014480138089806621996169797203363665524471993887054260561508591790480777947882428869591177786615146597640915549899032879511326374812649933704315872637504963554212241762345817716649791785893376335299332637750072767091991403407529324610496869601108644717671848131906165304530143066346297848850220648208444704992787526557161213576750662279444808964082715093421935936280345769178291278734387394908547750319412729940649249713784814923431184529575702040665058928423435329311570318384505806931677718100489374301165934522105670151408328659600511683500693555578275365793387486701186042482808230690195090432101944179340991532508140118236307439154788181642978607763511605177445453856358860681659460;
B[140]<=2560'd287061391028919331880511839719103132604223263806420906471353049728689558398395404260948301201712390775858606834605739995597456812229259065079433749044915410317112568245453552498973813998483169887338858584353314634701428591365715160978736003931467257176016908122089672026106267281212701594490354229876872554985633282105309947284241979957803878099783793774846196883429754826951045940809333599998115974596947062826866670652947127504187474854427723250026143923274842675142792455273609581530646772636816235718074282832200651800957597326342475655107554123314286765439748571887923893333820661952248522126658581849745457032824846552684859436429655011270733070497358885057017626644800479994702409194612559528947051111372941271164068413779994027873759988537048707312699111459013700;
B[141]<=2560'd260092525707394882598592749094480976447470788662984165781832793530026782027571985535011570224144194191599050882982958399889401312330818728340741138040252789032000767131611199624328446937270880484818878957212950269764002790262736725523633162545099378523721681341643397649779153367660036822389569559344494056649135052006656766456900294594874815438958762571936685735387963346165211365717078004165916763523637244723731743748970287853927488619923733073476055776306672786535613788112868713266693103881872702616766830753774749347176648262729344027259935049118433865243685728546483986089379915150912904136631473205761790454068360921347566286092894542741737903556952180543630520411115568287653455884679134832512342024337148405951924993505563638203561980646592379393605749411431492;
B[142]<=2560'd287173788843272458376571808853978276179731857093802827670182831998900968651111002260546749402262081977242630349798431349030220507157417802584168259888602315513912892482273467942565512630029219321573348645906459980660987040171401549210570967886557933478243421981468950726983554917860628165390647178856128241078590530722466564639257178010749898295615145001365881285373315270939073552085371303082090808164415025319641244665676471912984120714174115240131912732053761158297111531511272225072253069281812972589158331381831361356107117874147321940654587618849718152086519206627465380710596095387373327845573670903993351394111867052292206381578309947697522842968382509969585841931261990319089088400794160065490543021703415556519708947297562522406483844269552140424665934592230468;
B[143]<=2560'd287061390921728321262344074142857326994928616960924069430865418273694102195319973591087557799960308452098233804197850211970789407908596238893202315297664630855085675946602725979548550428189709947881350309486865834788289887759235175298078792573392750378744173732730554965414286924693126147088223508547105127860832229015768926812544694075842983692135779936776383582967391670941792221929115555294133888172788268191839949362392927331514585048472501147400171435930549523516093840332288537264622339116158112320134484894585208923268282661073943442364048329933483382126862872476604638130441166978059896725453078686610268238492815298480389742964728808764318805907846257368352546298261597741338968735072663711180812651320549450581867967504416175407847940164889117616629519401370692;
B[144]<=2560'd259980126272148624356964380452613585894698170878839134890101542188257481570563840234491530462125206398790466363588229128508376867665327020036137338911099931792400430692520537433524514425787450610875379757434858505500420345705932054611616005222031352462361392099015864985503890556258005567692257808755844884962226321155816281635531053227486519707644859663244113093101332766205605869468252565664306330361752109490407635930201844090463949276090573731117559389931324339041381018587851125649225312106932938388150146923182454416303370125751424447186432882546648662094629861673794901504159638974453524877593806923095793475898797668381618990306164509628067892943237623980373710949035171905488422151148915860425151575211029682812941169352371466883011676079281288687320865572148548;
B[145]<=2560'd259980126265843276452099007469749539645896728492517073900607709638599451537337914714631216536097406040889351596641739462116611171514915560060787834785757043006464795282605159264445405141305610244463496871093737012504758853550033324671330686226989334973496226769642684471914104483052501434188824140146576682603811266075196576221691496821302893807815732148193315141517245940257951750892666885114444504225713591256078275213519088746137742659779456668699305786720308192179091806561663771874996373300781232441534374876194657639887491759574392621641013596175972968929901639196688627207304573628145134364163809698333036393484449545033204100451275696219500273712209231096121469839991892413736645257664236257892566239787878735263258164199687827097854620186156089314287320217961796;
B[146]<=2560'd259980126164956073994872675674818833886792570768916260222837396721187379350623494133824421308960765240747373588035855065590135607542905550314568065323527069380083288715373202278835758756884807817920138083581122806830263034068343276577877762173612466705946817905897993611090282193244660230840082178960371468861629172327017526042520310116002282203592524219650990610570905715437476897245504532268178229177986990586815135708827385400667382579857600572469252231924731565212194216617987106881968296830786769766281967843348806761392883878077793133084311887001377502712955154261099623234144008925083739921209094308693920519553064950186489993786462178426148331784211967464947930134776111532526447879693637697133114627302925464405297054116049742802246485762648321095972116526023748;
B[147]<=2560'd259874338366637845877887080723112614413890308934386674754478033709363556416856322623716047019715499712508261079545755147003151433690595969508986771828278478960268837189390817742587837096140728061887963499817965687266441716232942746088264780200884659208002323762821019958931898066367838089399929690814521663174495877815251779589069597501556984777891883779565463209214220902829385476217871560162749439383624680539557669588090961190198678152998252900407701629345901125298493583389102325134661546608932138554439068469260865744374712618706419773700778855115052453452540987204909058963885601602862911224955050441198267388936259949834484557506276092495607760083346181073303148868366332056648548153521686760844942879150752867786727404371574875346858595835028562781297885874242629;
B[148]<=2560'd259980126164956067582301290703766329651480216768090942824715571697438831733394791437367857154058102708772754109000297202469800508964413625357489338324428601981701853144285161051549086402222040734812126404804653485385570372887161286930883398622802973512270991284234434466259004952782770513791609224499780351256914828938930978429266577561597265959745663882885108561044641457773059635862313986722094310974839010631202322164742195163550838087325526151437571692620669479025629502684387288712306857798649585126400956113248297223578776985084440622622029148279869423459995251052773255393275375983763593352965459351938594940734813870188037227566012713136756284707407338994071561474594033698579317071624229854429191003442031061089873204704662456862574350983671681896512818712495173;
B[149]<=2560'd259980126158650719652387191659961597237105491790405659429022208802335262944039319533136930897362512625118502350603787738300067188682241385784630467636911958633716828080036274592203716825335103339833761172570867799732297382529774304299993843160679072729562480571331262691097035669269604031885711896405966303261712937596411054963076934192376952619106471721117566385073417448267853497230641750708163003372685422322368902243112038544106130788292755008965697722653650675479349206504357268677296978602426083451809278784598572964718467808036248471277336879177146600573189236178966204582525835875256866047047732183207662269384801177827502368584498614185170294060289012563258458038820689578511180657354500197442676612551895923456282756091699406534083598592983503212121165642679365;
B[150]<=2560'd258174708622170144950021118199695519713927916187244008983524714844065013505233553951714388220503958511084608056146799340085923997213162668522661890152970358453778390585648364187511682223426867604965488258532701439477015757826361467130014014256049623781794893018807355756109163778273822225444603434692963141626943440661465328437696492188406986158134882314527526615493627251729608589693805263304911950748809259169949751187806426880805915434943078596167112246162316291048999334364938519873839663342827364973187752253405130859464347358447309086289400620522964884934225221547922585097257810970807431625258677932962529234284596245381225910056088479147222240568254423093517655479311992886837124971342157819469004490890584883007144704612348886844773108214310462428992530002822212;
B[151]<=2560'd258174708622170042348970691232675380671787523541776671414264421696984608343731671853021996890288639052427079659314026640997316501420686603693888201947388426389730302637885900481808021267801488134125721663262558176810215200451873672905135509585625685214055601986402081680386783470004666130100322236345492507654962569876329569411697220401200151343527307530492189249015471340295219011471404646390708779849004367920807527599164697373108422419040906884156359304690846422622068144667026979450542798314176503490838382774061646072842032938200003928911438841627190142246313232986070496322255819011799478815886130580848591411632744141745831605305798428166311368188725813860901173023472189223113426777110089429928191489517483260440320574076714561088544591176000087991668177673409604;
B[152]<=2560'd231093445486266393126042524288450115909240141933374170793957431628438635185375402780015313565933279309492646613976902686203188318111648991450768899805521461764420346621476312908139338815592890999757468109067095001283799755051202575058672427725879415358239130023876469088510268813900340718631634016421508823223922700574788914166426554507926830231898443596639710442022943450767849328586350632971480972085667476629962285144588348373707001934990107915029632448370482440634174091745129330898897477276465379892764535681012858947338163740857823398662502247976576020447753353037062283459150048923179595035978886118322742350245788324827626203670339391854244543114984694116059535154921173239251944440525281771302701614588936222024087917836546971389193934371631665882807625907000661;
B[153]<=2560'd231093445479960948984154420722563942086205711379180687255077232915947715675317099938376386260844100209795899203511461101891972252941401107108099785721353949085360683539535843721894570717776293326560641187111912211377290757399698733955793414210354789200521219007236622257587191388672584696949310931443037037928164538067809702255723933792706588682144264783448551030113128543497703804445148215702517138787726554457358710446093000919263870284951288834607049134342727402398608674103220292349440084710005080976966877964084525248555705175442032336588142224215364961619880770361115144244913813596013000156777703527845477273296027516355776923521274066964971156290933386470338780342794242583051255418900686909779657268450797765292962099446397791500461986355217009035904421916398660;
B[154]<=2560'd231093445379075382106991178075649746245943257482380751350947235367856467324626677827632520246790517267069349961030075328033810116606086542333844867255636692911596509564816473031289762101840348451220889680554196220489491645267692443842707069581222416768920191407545499332212869574089794733983211206954857731286734883954199965027686827959618361707953753885337633183190959024154668269344331570016662826271357185714439306879221887501544182543074892579106925398143147624858410835392803243323748183818634943696074130277182469115775842502168391000731535584880122882237960294247901348741049288932545430893600570136614805223579710629363159404257375389250778721343441208869446468421791592851465703447489947721959282778611652760826885597164659925649639152506332888863784384639358276;
B[155]<=2560'd231093032246373768407126185749375898989322909050022103407978373577886040093297546766988601857626576011298084919628429112917414959851352427114854377224542155950648720095392688280270834651972440196693964630100170559264491253045730116331632942531904856126803424163253921774463813952811979364027708544667026209834499060063162669132132524863913823261143158390009753202684119388370673992018572834370316600858932149821542735584789354856280617509011977582366776715123318507345401833524591532479684609192615362690664345509374062305074318273272003833645644388529852992868146957378007424016157933792370464313586416645135304534373881357823271566446542575930027718709037084121044214022272258476278498068349119611176740574852521498269280365759654027240471360160339743547356327381914965;
B[156]<=2560'd231086420609470362158746030186711036248990207031256369550028166403822757724820330142826154151778953564350078846742303074063015043411753683659803852270704770296177490993725164629421271405546054983717114300804323152607572885957657408562425603586087686550050745744600196706214544888120921018755156403883044750934318088742244862665365375566648312283768889939919005119902871818223817680200678572974708667105114388160980825202482234183014078153209775849606409704636900534789537120998713648130808371249598885073047780760941099346917105009093556933021046173369803361720631233276553873126746018224620238185435065403580235914431780634704774719477811559212885975321322710417851646850145981403937361233764275267582305749894749273283934504539207469337105883735405676951514619637486933;
B[157]<=2560'd231093032145488201529968653888856418583621269922350012844018871892275489125470728225850012407562360972956678124124488372360397364932676287033317314492592524772932236915163246634041974484616511219765841883327981701098528726533414497010140970365046357513824250809789829431471031642476940317076350791267136404606592525959200546961161992904866627549895004085670150595374555803391746067691473543444328063669991105834490053319478832864918670110199314118343753965424668150365316219243119268988673799129388904024235164899812678332924239999020737262597850854069484258676750262124621259616320965000314236156097485367871670591015215968874570062514805859171804969997635693834563527839014349015493401921356615218381440045537631628849125922345604474422456319411377909214741499473122645;
B[158]<=2560'd204005155758907597436024060601092282099995229093256095281359347897471581186378038629636723589106737007612409009616327691705025366887207108726267877292837062505989600577175180622691690372842416823891414332562906603732203417953351056477115307249961465070447997610471170457779039065888692938817567410728625518888494240854125568340711201363296040125424338930045201703848282167213888264954570979108056697913955935974392085466420356158771818247906157421307718991415584096615744886976984855700741050515636625657588010715884312746233303879719180288403038168731552440922564735243958162290899855142710648568312847995390365593834238274008661157401084561053945706146465883653572625303028190397882305907188301367854609455758828765764205073865407395640691471688554764453342730427651412;
B[159]<=2560'd231086420609444192500348747246842220448286212547682031861375549175913763493666281389324725570743847492978046120475118866192311467493283521978761691203214750357606079899560829138871682083376038156423723964454080553795410042624888034245659516154591273451752053819385293674925658390581062055611373754413404419401814659029457672486622020922201924154565559365774535974942387050669068141347440563953546196506310419955029218687125220002257567765657544091352895115212408693742158378243658464134833387302716855052045047906843269405837972179769244895427994248136668724741039706736962646527500920601618759943042641930207758857791486478537858113408546534247849183611581431030718361639804121759291537014212257469256316092537397159810870443683503961929157131902333250712042141170095445;
B[160]<=2560'd231093006419248303753535392169235801223970200415968911707512963942306570666408524184209936850976219818237261049543098908689062223071092294189196170128172047299113934439181497094432878674402921668306722535774058138019775089028104764131336087913599942222035513609191376924498360182371407562036996424138711674062129594114459013263208196215566456087622927303892985168619323150440042261358533863019080332940555000491436958200876340225759749520144246178945618071701112250423616727031156806394968565776563015620740930727239362675910191793917488147911468841662725623823247196848903466857702953894603557229450094189043295455384356601727473731294704511782695507735543432877614014345758655915916993917118386470538278100661106963520876310873701455312103621205480550362902547964187989;
B[161]<=2560'd204012154789292576160026423358413057498915540655738089530575258585660961489704757200453283848314746330446796490160488180039206620010527063816623541353382358349136598851130904895704902438175289528865409307168332694153229601203820264853013819831792374656770326703695054597897892243043538994683595994555138828434126863638195579827228874427523825649424737755812819593187932185461657969197583025653378486265052072789090834798507357316865003436668617116911066176859547670830920485337779901871476650245541821353354859321773620778655410849424108177411357433216074142922908562372388309847722786576688539422920920380508081955491393126317165547244673929566018863612605228399256694391935238854086833731812015433946129299163705135039337074193205395329228182064915379682749105204188501;
B[162]<=2560'd202319575843300227673903089141252489974460714311146939962430908176120128393784599257861181650423306959535593001152743704727771515753825194125088596106109685374049535566397966351880234311970525676297096780362146254963201892339553507960879955117249466800961575048649154975535014740150791261210881285972823241187730489895926222375880997568488398454093922406051414906270691187110237988493698616560694215295096884881086802899407019718482091491988610600976861621306449102331786432000813646642832025443552301121101037732830559510993677044241592339687646236301577704540389501949431851265749164918356165077520028445318511172471504428694614456635228139556773936630654115241218513132339362236203894849763128751409597855117449166475014838667690234849313406907743100851190341760800085;
B[163]<=2560'd229294639681267711357368503479596289788917138323781661056907854972223647482476618928250349452152109612550769890593079790032675939013147891929689968600806730716313798877535588440380893097131731440698181576704571319891952088946899529154307109285846362624287104174979963406825146183517772223174986449524695116541459017704312285205246070367473581677636941158242008787236773254550503923680672296627345997438355538586119074693241015946021217865912090260726175688863631136850839343590535936469643355227331404641198686532728078783113446134531305654447166736497286389150060851256711316055979204623734611156154491526515645045263865175694684599530280877122511251580496095522499913609719783342559133111353183891263416578979924597268722502326434160808749716851401847437461353022182724;
B[164]<=2560'd229288028038454677028245886056513491186047260841816845959775659174474491155253241395049846761528679387069517747759210278648432013597318421671170723855764334798342502900990924012980016077831628024761228503223427439620646356547005836103887315947249079011804049855490644166499418963703032995662095556318162639664996734510083787082177544386189689435475972744043220738543020391253512559590634682938742378368642854670390535435693475756481890502527013074466090145746027951240038831884341546574586561622020029849450857745467454584068433091223792840489328520872253521093903577439511730715127016175006939102957628433798036130210956300497474822034569126990300764302458007624183123179178844823719568286907206925370924879318415070336522788787932442590128184194579448203047650364577092;
B[165]<=2560'd229295052801360265178448360533930584056580189850438400410513529700037394486742326249030750532125898490406146154845861746389974443262786792394023512949960356749995769425336642408270495539285062708454722990917164414080802956354366214121575045160002462786174120602926295174229339647104110302372869171394309043364566840544260228865962991965512699171092115696287169671010981166899860302217186411603883848645263165875689893004794728193222620142529289872770175814408933947612083904365181797708293406846744526109316986225524846668888507358198113240288259333600424927853595315947913388767821480346747016231589076993743997162961187126936857238941574869610536573018504307964590749061221428458887708978214414530833889915997661511878843983296117609762336038872790538127191417917101380;
B[166]<=2560'd202213815485880916619604627906558872079663623278646930155399220419448701997387949725761355385419449133603388076505384434125285028317541567714220613093559587660162167850511508416740730455888302335443864193673344797832109048854727073099041144843919410792473661019095303896743798279530432965189053412829792653486292193782055656733610201236696498033986248258773233200581303766011197148082496075809381860505470893856764556202332598472631405545345151996169309400798851505741020631504283991787031760248847496970342037061272130352766868968265394415724740441393159123362241741179317249875964636862387552191405383035029748161336565238476954667774735907252983690462150115477969699090252236127185687343143260265519459098205126416921678432244380755094544448431105777482526836433179988;
B[167]<=2560'd229295078728924674313204580081775326906661853341544142142789100985555397197149698026858219826187179828892149952494704072935382444123159284203518725449112732593245504108768778716383585806579829770251559307226604680015415586285168576553120876423198120351829017843507102816577386578467481180083815984527357786481838094664014172582301734935844232850612727135782806409886597959649212886669265291151095419573221800068597431844868590823878079000373765866672182864553048505291999274221470226558917139051379477657888839495254635818517146506340824975422345555348481219572441347959235918113155631085491724882736947415382351806228586650185788552925413639767407793207115869618364754110684258002969764214823090970054271294152267813311760700371769955462237453822442458785544324718613844;
B[168]<=2560'd204005131646862938950248660925251077798403324041593296192609332811564018150838678913566825595399964116836556909715541458515235569212514191750655957344842325271637031430366714543932303655377154123347836294336575281208365873934835037032465392886100316971122273369932907060356598840167210082697675463147733353547105911894086236450923115232065854239002724946928667042119758103487515043007954852149810233681221625654190578067223640992567890497591882705286540072059542872582721653900416973770201800375249201596503726949085161948630037875916062339882684593509512091503583271859512228680496419365984075915046185091123793308504470061572440910690525083341975638720915136225760480777080242322113794815378478812169049995328904162035566172636733841784073625751044323204881196720149572;
B[169]<=2560'd204012180615997684660888265430101834648599028215049972427965307213678254102643189961334378091195194526037623462667330206424467315151873394876426159380685623841334068470535108598613238652663228077402975682762137404899438704201533833504333200839729825557514244668564445414648028382124171095863239967203495421111337961139406794641100921879633871236942544697751337933984976294628666285698880204545835312363065148350581140108196860671963706576470107381758451068028685840108068234462637301081936268384192700597599297623390011340678082640718202610686153273785346424360304399464447479934789907991784051803192366185388430436338517275411280167014020762895932026355543593183788895783008688039057381990658638503109361953362342397768564585293774964657846455838051546624410008153314628;
B[170]<=2560'd203906394431874702272089629394832350959578873029663443282255214919409125864416460737021532813126728757282682741389046894501673742635206142761407950299040144733240850050115038230324001297702061127560174048898674857519299774410698497599485545029705908568181716794415045445609528667620968198666373614102438669573506912369676457953932635695126130655914360087368664575307674568843073781386689205340563488512637347650255037302353715183296943243227395948570729802254234629477074984786508926146710617926101536422419532872188525762739877937813426085159141788209276381182577516544680997613530270187738064081441139878577030946336132123128655081100085501566141782895500834883426188986379849882416517963653880594907231103683386087471649729950600988174865265999090851376711538324030533;
B[171]<=2560'd229288441171156188502888140171820960621670018868972247372223703998761363201495464537855320645469461203983283157311820410740272761221641659050507280080171700029880321123211751724543254448947906053844739767876089782835603543543195760163694095611512528901985593802299674857238013804073295105421817997383370678981004245799928017084769679094465626710518590317742217787640231579044337017812689228193009880275510484073634368381946728664485073927033276751547800347099292665113677239497968827239935772904507465139241147308692519772065898225499843634192033496623375960290484979024611829834794391821683445144228754383917567913486119574594223837100196851400901580508658279183983930805499411545434189198076515361476033970782547182799551986264226288009333037110150778023470665766880324;
B[172]<=2560'd229288441271647671111034255044959667831004694847297155226592520416017893323272231084011713468823555516968615830573767644616351548093770861428868218147058375792111022390056719790295208386779706293726152632315582800814410802438590250554773908754819483196874572272752438357284853424013626091111013367201764354672471411360921162934906033433650086698723281806026916456033373382938280485563689807427249900015429077918051248495490682633745214478458771075590354085004345399229876234542491421581520461638913418157029236461559082151763566780003707841672182927867983086350765343713401674343904609391678465142656438386337656776179926102976718786671343823965757141581704920654788098474814069244544591811085954189713848398863496227144109766860555158021639342043449546685812608773477444;
B[173]<=2560'd202207203949838344734325239087857724517619770967131578848353508908116324990527042726427776921623077412619650237427015522432933512601198155223870733609656883595927074611856620386770200851263534616308693717834719552190158178637763588703241096048737647493221820381840500871159900496617264101863317484693391556302059796931489886752671459760100890616633777319733256701695089178046530636396115968984291588385413585295533022692378110108128543042800968749139403613983023999687886486871832745374828684352777425399432727457743546813419288176261036858814854498998390021297788298471025886516898222797810992504972767307314721064188087458894418279061906795437957052221988903822868022452092158989252251540149732782379140395293026186184017274090429164219193860235610850964975044206613828;
B[174]<=2560'd204012180723188605456159163238609525978060722333482085419500018779946675248705412331746682320259134895389396180391526969224671210239248234158717470605524989825040294221837496467448413711046347419223425229358534411627301126422751550073465017323023681564452021458508055105737160979343032853370309120582093433508118790517383335333478255109655283564899496111120311380453014911421383867243230804679720220238206296835849118489721086104250113581298936130031191350976565722117229068067596524759846480712248317109771428880081833280033646123223595684489477441228254521146134011915327834141536189696906089225847096015365922681621203509931886635730218947118642822052405437135016798384261333884333894636125012910609325165115703096740948385114038036274391599089251171731693616462386516;
B[175]<=2560'd204005155859399086431680624108465004758243909345781709238261153380122067882238798154142358482610003434051779268922557122696613722133857271370084197260520027620491745304958789902219510676460745684988940012430070211607565095246307446781893723622514773707181599770585492513726573612628914154785489580056456446441220402755148998845656813562482425693164897604413222220721652290530497333910643897926892442643771980108405056373078958991491487258522790987463590426175095245321762023071869864935826070634613004708435602757659963364956983325487273786435416170187133807655452848295432083640984017600895308341620462339128103880287662051338479536237001316676543824401016322588285487846670892372781730579976787712469793593141329874538204894174721557300385844236020332133194509204145237;
B[176]<=2560'd202206792242145464691919084493683485604134991503026590533149267839165011993375495863734624521592314341368664553791305841300752924662060917812686672898534626929165048064288278375344275684374442227285706745570562853155958962975152428390891444953978885945185661942235602991257108330496154003779819970210025996737157427202437853559381208235397293106555055739107419944744729138700334853331095888691164780515312289037984041470131452813833534204304214839965491430080468492093567006396943973438363335742544451732993338045796006830527123738326872166908980944883285031520028802527648974233958935502344013455581870165281067885230000063247134040858602703165137903605780613236240646184497730387134997394841197176671897060969455996278626318824535038563775385903276804342293320405701701;
B[177]<=2560'd203899343747657617389652787630201983486567463038163758606927486331640787550287914722830173139967864032664390289105698408951405554383175166374943124567204033182983390331994087123899628678642117638766986999448408064154362184768998135374106930802784943819878800650417743383064202050598678759221265793615912567063358966265122650754146939222900309526777620443170818258463833616640741916052991775850317498184171818680639429323340684408804012845823147262740859889671188165426284357362606534867024221022807893145905745852493598872328320351438718396764837236837799445222689386291114328375556187646259938898184256511939550192313228684533999341031044772954940161102591453711205458494083285148997729957412380216754010251151493294746739267408225381908126612036390819444665638802773333;
B[178]<=2560'd231086394688552847070971191269254245942904791780026747027870077453794436114624368044094205509272725064374093293443819884111957328842521220959957052239850965555558310946735754769025911596232550093639962830471264650425834026553570468925223645152955172345968444327180983835080663129466133371399140339169606020624330478358169149128020622841241673466875357884385374730175091783847503380170730715176506645029544057258235529102036688875725691920024467554936711479544766418290949637441197962021378582105383666797028636848970257247672220834791877149454234639499288352712056361159112484589228818412329270622053132512894786718695826244743181180528203825731622244890134495735095142989071429594319601669787087805831977544705071182090708729507165138424203822026942664428516093795325269;
B[179]<=2560'd204005157467681522697940939114803044857820652799427711030475962856484107502182786352411361912397702809899606738210514812367829310336980462555694302595795299095119161508192861977961414822878392529415552103602389885088292381821638046619863163009991634643836684213088180994988231872305597520882376851284342474036438644777106434972735536041368260357164960173028223854786200114878572865040469503302691572067693343133107459308191960712346649703396612923333022528971737402766963516281510760991720720938282103514921043938405346361863413341113001463734091796281394179003726947806975335590761512429235030100526619702228228371730701006690155240552098172592704465807492046821948389714540217459866395602295615586844607509728491707493227889738057181135016811930949027318814398261581141;
B[180]<=2560'd204012182230587110470841218828563783643104136616849517406134776960094829013695663626532229783445402437641132122188823400878668352625308241428239795812365640555235267140004643557308795705430889577245716819988651727391602172326360935075387284437232824742562263700431536007705272290284912631874005691334736639241403938806648841911510726575438963346777407611495905356759887136083183344093132047316814985795452245897026605888242486115330183792906814610526341299358183270196915290786638753085523999247201592700854965327038938723951058600487724192964324027742285712767214155673553490663396253771648884599632904091495761217216649525329815993877358371422712818167014684374370092386977612651778693337127547086497196884269503415008394043684658280830904636768317308568961919338501461;
B[181]<=2560'd204012182236892458400565692688738152134290838513328052847322557997202108113243857546196014052352059248702007731655049115923833295918930858110329236800829591310913148788111096792117548170864206292894961387696655146788104910257437023824604790965819374871901190081823402639313240031318116274046243445120689672832101845220893024379844844091479651651493737209827845266858982398054297158748293700489737700047571869736153054339070204944422024998268123423228731938506764848688244297899900110805380204938209844512563690988654805929620384351687506411330957111520740803586789069926036334914482545012450659229650631598933628249776971744576866445277912093252791355074129267674464212715939133171515432253311870414788675900192313006252743771172030891834591552368053451920369181424702805;
B[182]<=2560'd202319603290506025669017752615956701451031318071651291335463600531560195020227301216754526755671694136420828907192981835835398713832165169829276281112654789128265017578877300711504213615018225065233465295069623226086240203447495844128024278553311457124980883027076312151525269242135013691391408619882223012946484375544122639629665469439022048048831138368529209442833426290039295364016301965207810777434515521612931844380759816903876325142059541858040829052867416271644057035448768366656270380771806757682513949201677847909389754833068516848933739391691962955692720193955710276043257091149459266465717384390875920712954523162291233355919251706283771262648205133118494589331440546616611369434419422705494733443916282006193866293791220887253769519504284522649342170358961493;
B[183]<=2560'd202206792343425116191992707545525509637253871138459865520885564683096329742258182385945962268783544339208591168133695709657823650393984986107462656223107924547475001390410438439496363215232280597974601669136944159576092176707894670587410340068783597708882435729431035547857700813810657600976252106068281554247985219491622946562173138851324102314713104094048187666287410521202007060964586593390587908257870320720891702476214332513060919632287694384668316210913292980944291096423533702456495255312328259869961703980617105595752082959328978546421866772746415703327665936326986139674835600069495623223065530556235031935242548395597619391880513762287357154673293947002344835848424012645209850891375808645234309806072711863627576062272815218127566901981306626286058415125321045;
B[184]<=2560'd202213817207242440453469275314972981622396236295701371164441063911520131673201084317815815769170032886201655413063677829399098684388769962949011107718637096562415614193698458471947377393125741140679428304426649767105688587501992339488684695777108097819050742023662243512347583431373808965832784018285271849887994540384822252615562335909633806077485200091256251575464916504704135553079530320219267973717621787358704067707014064007778020923099071533499985688058745885123669091302603388372881773719665994184361899709135857532249922819058318702656067340086946672577712915728018258148856920040307580766327125206380975238041624543359130911452739428150312627396991995699240375726211565688144583729417012083247036512519631921621817253186456059938272058258005973077444328919749973;
B[185]<=2560'd231093445479960948960659052264069526542095629097925303103829162582666042702565092374677295022478505297210687648746155497755920751920079141952836221126230829329243762039410338893429924501636590644685703155094843368190394008104632488549542849510154795381325102936525729927083518831111636633668837289315355747520897661731071389115704390474505736761672824367934824868609668465153427744911803794043727165566658689835377087574819991560682865128413038869548364653256536962837030050021619263473912494196160419692729662310085985914059480753758845532289268133202186000265121610066334632119940990447218819873839707301755361923348535277439997707608194936985498281921568817595786767260908920840046931261995243161049355411761588010804687570874487843063874212094013949605489271306016085;
B[186]<=2560'd231093445580846515814327308764161797092211252020983865527240908263289742304002972782585757079272058413132502992745774652562778564912653038350971905278903564075840542873203152641722790750096078601396602894013218107178985456542487326075110580073634871567947564810027839662616074280312347165174652160690323577669945824881331302787576537028397800692393100150692702066048432043216435279353470271829441613064853165449463318806357672317665560005344650485318032798511618996662291008227394861699358041377186877089981333824357633398031487821875798510203921457647751830721999382548948826579510713169846325011808398783909915136553379784927368057808719818099684765005915696072942220642978668172424663743148540645550427434349458323674227884248556727196942958070107622816210619639092565;
B[187]<=2560'd231093445580846515814327308763820072487053360769108718688623712578016000007204839846303735333882843903749197390456465427033236712370223393101219737228886657105439511744689511379153566964207427902725174592270916541936136012722593463809134406900216932096096751933272228890702392322893363682712709510483283116765684068975588607919690886855253254248775620645032238214715310150541336373474563540919602347006802945420087835718031310064774711835725308193828044653087328190093173333035443927897884084333894732602762716045996419898544988924252951073696562007499058785710031422429169455840306147244657308010653644595013109131506324702016696801357503436236673237096950033288080168195619135184278740137113922555255043228262963688591732307698812638089604984523753929197405022530655573;
B[188]<=2560'd258174708622143872666986284950923460007365983196207485620461322783193176972719014845787027202845195668528917523666892030254966492999944649378929836450597124499254639124176113356440670662814331184027927719105119068882836140838020342871480773881408443869714044053924702564490999873814844543925842354274989176350500612177562953233055887383075563446662474823579729348820519345886091711036318966611306926827096443722552015726644336276283090882771351504751011321179009871976787995986309659602029576589261641628023927635271321114009267536194043050130141460454594695142633203026519101655451904805145916026515239304279405333731939803733357866382235441614681471142504998762630192878424910151929583766280260595962872047547156796512248104814609790729644231560592106028865438984000853;
B[189]<=2560'd231093884533974065781840545383045929529469521716111776839424268314853153918447622526947557851493012790777955130927641667791618502179268417303713773985655968532955280611835971411148869758435432473552324117847653609642025563507892430604861010167411417041231132627436040041314810370953002646068607073453115047809205955824143771667955551778497234418187494543155426857504722979429955076416838047340835424546533171543280992536052879446519366798253672580660034303966730747560673474191153472440367350610850984689535408443928682503515264886591560478662969606896978074232407282904380538767984687399137636267609343474920283060380799495800449549073234996034322984101311706857444820426099482427815202623830238122343980708778788200285247593166523272884440161216508984094653315923924309;
B[190]<=2560'd231093886148141596048948578518791971278851376299661133959111083948498666869811669109495222692690861221798641756323864768619258979279904876306826468164707575156101419150469367626500118870090283431613053577807861494284342750143111786032960741952941746280365948418545292684329272615622202579517642594671878846025015784520334347608681730177384383508516040877650726020600337539760143246371759343852476053783080709985322844769562302880832244993022920938584811006422755889213016469441087243062530099994663984869988482647972213299087776195005294225142319586586662242021924310231548566299694115715544953052829502967162274034828031592628296373352076912205041105057202539036884729750769855396853150396269746892740656892383976791729962806485098232784467500907397884900641704571655509;
B[191]<=2560'd259973073752679457445827655963519677475377092639220148323701751918222085479367868052017441496065238148452689512621578598880483357328343018115077382680027416268553927407117160037116041640775158385944775855010324327658614804595301008106810271830512566667461049855013598283606334928189627967068486301226788916855944344942571115070706471488292804464298065585089625469314677116358723771562777051165411786784276629081458327913889708017917640244110852836587579709472106122015013622260956578973377142576160374825546282004374486679065741295171132050491487908837948959256916455737805533386705569551853325227169621956857654287718964387164924124410347898841959924314853816691792464628856969635499596966265843171646292430843715152279174266292044483702017323987155183696356985657447765;
B[192]<=2560'd259979685389188785460465944470829881251033567446823222641193030391338596905849906426165817340056798564659926024115606990065087675140418621059920547563856732221260095854362408488011835433524179357552371018206268320990577465685935519256813958346716293237095602948881705585139549002564334763394784958295877470633007843120718281826078371490815575014188417025608803929451407680455485781209676463347201261877109850540597810674232174119887751190583045971142348901276349963368843404178069967481590829956946147217991929599633121521185737855847936648699512499022167437068307022824069255022917270469797920517007918390074804587386035095132864204008609158225427920926727227267627043602643423181099936342657659176705251235357115410550046793741113624307001803528834959293964561092531541;
B[193]<=2560'd258287106442802353104648515970185636909137197009596511266601284505061462866756043543414069350054084050126161629167320455628365574249596699078782953634400132352074467540817923671307378425004715739852885011802251500193922337972881648259705831655520479745073293209384172756902351747929833691335159979816864253626835870551302851275602270082325147178150509003482435258718068595280742476545158153144853621527547227204100740681679538101405285328962876353044987137958481893727509028809007260668002780328803088251467968885782586090195441098784217624828886086366402103113261689800169714950461432621127188672371590501153155874055575861454397906499089818373159381429593064965038207847294854010519706942837027042777308287657975602086999994946115707308699793356695350371703184906605909;
B[194]<=2560'd258287106442802347092959973804359083687640467220601009073327065326845475626394445539600563585555040323008596319458301129903318498194030206856091979426716540384625195106513894410182753334308710607218273949566339394749793208510508154779006313436799035623025910993687568525442822484934825794760277443543952012127868781764234873969977301211360279927813129226827514185195780445299492355316188180835669732524666638201582576066274528109418728315411457329710730224336326677376695036545236327634892113544114241907842798408034470352934856915986108866396908286519249720169261493440159463880080113513023826392245072728803989310534128161867300855686288756886355108226001734984108560260170358037506435618266849859917340077821704957061555633647971332991191254417071723295251675785549141;
B[195]<=2560'd258181320258653194671404109596873521986587470764132601274133609325462630827126687821089832159064473320056280550127378223504774198442872022470294174447568387561472023038045122767087036544823792132611904809364207782793361937851668199140986077252361682032764015155691550543794696271108778147863416677861616715541118739182269272851259827632214307126451372149597538785135601259805048461342880180416582454674734774718502918110458006823110626656412332272267420248609589454965934622688474554287639914163327240798726075191973055927944487341280256981549281106798034349216415802477483327847453062295522728924261127844762191789641857135901060329217467971044432154803375788767765076999388709226434841763541753552093511175604245174858836015293403905851623148670418157835335890237740373;
B[196]<=2560'd231093445486660483361323408907305418868567076442482128452815906386632134958442105404111689040411425722662186234352272490219805697340870619165045251549003167520049291350940752458518924051592747049797826643309254769074816385405321966080865407748735900997772487813619131705889776919860707296194903978186353022871313286554947489925847636651578283126572053282729549530915544437269473829033362998371265302112535034814184804477228603084402285584372260049554570444440527813193554387535431201908877953491767001626492979168151067885483375616975686578862492680359130384228064695203326150130168679634556518262331922018919047962420482359565968614893770749102905324090413552297333149439043443338912377978533436198479189220253433925757993053878234748808259011984575741726509610428618069;
B[197]<=2560'd258280494812598475267173996459587417690300315723127788138539678053347877603257977512590516085036657767246050518593975174897650388608703943824954639211815733562599369495248878340129981438664666918954382401783194470650753165811961514039500194204581429909353656817307384976005672249192400932691941566557197094195248434263181020385614099604104502261876462651470078503059509438790367439777990104516856939345503033373432915602979517081177683313583793313237737571766523464737418804610773310629505434503571277919268997634988396684729919014844298640565487429587832622672369369945782499523197356238742176856260961514477290148499511145920192264012533110478631820770332918796275284174951188973312539907491955382750824055214424442890970557205756223197432088158927650774446749041120597;
B[198]<=2560'd259979712930950166503092892632425040089291559025261300485193886471615729424100191793072430631581059391653504185977102655344500137951262154708447329188569284663730776951683772121517133612259725573701038117912890291199788501386819611396515611367599635822733761871927868865622779327266473789628655582294091296282387618603366691082751724257720513113956663640150743747774709936385973915488170274891552806914568948832631926425442824555219691523029215313723489722840635581281833790799563890951546189762671807145863932270066179501957573698271989349661564801967975293210272320968308163627762183577880205689099859450844762853288116197520130642011025999305688596957195189071211054842234466653309433572317874989191210210675389600626128186366498307898892889183490266788831502835995989;
B[199]<=2560'd259980127772819789334666012802296397538061819072247983763413673389767414601292390416745377655103722312110495504047717834711412764023051359911741956702512948636862647858976351132981254032174688194364143711071080590741820050827925818042183247336868008414416117948762720935981948571923932268999919537821164229588608290124169704226283892093887364025716796193960389306933391587251092585550864200320730318169756084841289657175959269931942020168627753213156073011117916725274250862343081879946283590625979756323734224512223723301972372247645120158052968430438985534750376241428384874944493370836899986430177133498396244369945026727415611453339954229182621010888340681257067680376682690526420481636035395005170749334976845427837578061487547189564420078804732133571085997897504085;
B[200]<=2560'd259980126272146982763647181253543161900733419197463580281873068431241415111530978691414741208516491512519267083863018017232791167123513018469653607592648977166631525703508174532820577648609687312475323389661296189693850264107467841967395396333183561508889657604384544057584395781436388491489599992291009406882277276681537246060517581765537465266734455367331176273740833186978097880549416088673327242889442010122186952519309338807181684791450943630188527868479433781973619449657555096435433494214151455341054290357418361003859602148373051511094320658736853072652529533108850171764993458082022599646512558000255783143714443248745698896022388156573331946793079603587534343912187294828144447929650310720991109083387715455605779478036085094190395357239199022357697586517071189;
B[201]<=2560'd259980126171681772037652650891592752749243251510398602825393040470329483131730834746157949127703716791592374447343334013299633312441018741165196967807012883381207120711528831215692229211409338738435861770660791400557755981963024287575553750454815429643452118582572794411024981121997467934411025395171554578443022108514241903540274966667185630095970874627718075153056486524748646009994773428972178390510837866521366108990713421679167299642088139587070323517955804214975064529266436791969585375525616010873178611582457229529519894843249886299281894059484792029545973576528936674376284872041396946154443663008854315127084361957266523359336617504014231337500385069688068743627499219672203498978228651353590123079178741824271017064255729682523696467510650826742649005748344166;
B[202]<=2560'd260092964660497802300766944965579649220423760328681902547901152265724909774748694845540659911515519657591280354180290840887413383578734995647263063262261250122154131952050794893235665578284854830256355229730834889179374987480007018665965213250189368128116178622736060137168851882274595091999261105690377672658928611058704194762615470955884938146202996985780860805650582971623918495987449836972590122689113083905738590788302238800480831085795472335294757658266426026664481481521290036238382042657623629466445267746449057528990090440873988064666794169769543214104317182087316057295359997152857562230487890184630634201286054677890889033146122579711259046338743320741197495264299984764085732480694178979533252549850839204704663090383945769466706556682332673222615156921816405;
B[203]<=2560'd288866806849951186600238962038583420167180865226211456200228340452686447674645293307380886145096012935149995709219763281223247647130002731165852719570368344036352923692505860485913073375177790107814886393867175989426075888632022594704669622288666097759427772676282731704933309193834700152559176352806281196980927999296091501775457702733753552779271774636313853669597613163031506443786585975670571768422044267896760577374223341613186983951469157148872927802640875109748960633975208618970842224186245424793479853686855247830184859526748919573946602410360612787379693324820061618891427694736875635005749122825843843114709737234720903953037426919696639416759189937121674070395644184578152257553052669818611090164881971037029807725517357940412108953312182016119649867762390357;
B[204]<=2560'd288866806856650618775583446513344500044000000538997212252276535365081895784780608878867104731789378591831995874442097696956408009124004058832771355105374232412206275449086736207799689019181983451765596492108702817960191189782542915618894494177746615119496332626774388437835940155273703540808316959186591702252610603796992883076159925577920206106352318494685813057726754879116556612723029732148600667386847807454258669661862119608574323772729537007769433751450457651165387971210731382329891064143708073916255349167125213239831697435993030545112283531930172442467210886203162754079803990475991162180987440101328234334246441575213276060404832718104254649417350875276903831103939063522663509335801537170040086849436115674508098602903760360809411055649078054051269627795035477;
B[205]<=2560'd288866806856676890657735030936709480369657514989024951186898409798406408095087937088400401916713173314221632562771981635168039152223989305773671834137393653740661635271682733352214533025647238442362744224464978974839330044551608979196696921396050132928578076495466523007690643050790518153435852199056627438086555920010449017951126735358216343779528275942631553999604143657737718152056858516189745959447696477409594726247563318284119140654792818177134893176824552497426143720235402854994271575482052369339702546762629278561604900895600130942529626755754670326344957899952009873379264470398311657584413385570464070563003729250402268377878792308653409873340212798920440911183511352915504561432580736210052503109457186010285942917855179004519290092613845702511804280907060565;
B[206]<=2560'd288866806856676890657735032430093170787908991064330105707877798154434324320729625532675356647882755162054774547836133280664155019744255242535077418500462561072109461855633692295957705004850618438938077978394181928150207436747476227907511088296932626290888222160138389456272771633323418061728949832051294372289018141940621273094283985936319247222420380608983382189000974312118337561353989277125341811702820765322887707661965466121418696091877330242415622796587308735870068303225090084582718502814634033614941106617068584034852879518294733970514966788417964149300865343929116098845736481896754223868001616713757526766984595462123695766433061990979437369348217368646373979766635264205483738860598955664195484215006572043058493432954332600078639140252851395810557652515505493;
B[207]<=2560'd288979645446376948782250787053676613573433970721619354671151236981127051155654612681091900152609337817320080245804243963583288008309633358573434220063891169298141863684777260365975544591404126846064038574524684742344288065639713769712327454256125468121935992062892012478387913762972926729387975737975775954233864052808523962969962344275342987173326325801570471792593649340780186341307466677798721929001691901382249471881441685078509511901353222297058098983987093897491484985632311806567497859270474067493335383736774573947539285663039324757288071509907615008838494445848423801214831629486613994209088103787706270610527904408867756731932689532141450702485910174304095160167322050247526283544163523739885913465126188332584490755289035805230987262744864354186352061435958613;
B[208]<=2560'd317753487534946311211450673811336501178740668142000749471325906007583308668155569843060116207753066410580689844617308627063740443956541971191833205583084608508930536666632353460091601069110986544617238798933080515543521383874085912558385283006525077725229907907675670080648486685870647332687802115549480522615283633691680576580666535154119034186527521918711209114429612342808605626755323719154670405583934994304083592927233365588730171978363413149896513531804687293115598979982103536584115421528209954503091971352490760725248911078625146299030530164184103037062147926967081882775801678030478855948317420054906627471870285507141280959414207980072205211840668995424824289466773470267149748951763634776134929783075639173801574481080239429104468419088705498630764478638413141;
B[209]<=2560'd317753487534946311209982595594716183976852533692889864687860067747810280704524917586462861309326762004703813195715582899459322543244993610742587592176739796376817150292471483796645886801345314022984208880948044525734244852516731849382292867069807211703841372496672064443053106779724022099382643704214074653582774347487029384915337669806806377318259512341097019152848102889169611476893738795429127660186103397267830220438939977432135537300877211515693239872610501046820911807037360737081966391703985368372292311428392883313958123031360346989741680362587410878397308362842847216456392174471038596810101102828181715001501406469531565628472308199654837966091751573165320898268550198159350394348181886876070378347783586605867500014936808409792979079209227556416457151297705301;
B[210]<=2560'd317753487534946304820906196863095721359691411162635445832818251135002682591219075400115264831622535140738190654121764484758236878841507698454855227054542408534774081095729097755631209910170316665560443438341029837154093533502535486691687926421622309502085328409574856191293180093272565569145469402183897939233998661858531309315645378843836159112545565242390278046872565031236307580437001803271609446122915152055490891568849581598716441889662448898359550545549636085044844580717417834426529280577824212738516982485089583031098199140716891728239765400834157344587201616879087485422191274297596562876522295967009632411438891097924162909891482179326198848644058195195818004930539379618556827579420599151859427806376441581523205484543765763288701319477878415393508529089631573;
B[211]<=2560'd317753487534946304820906220664260045686581172212007233377605044567919655095232610825752140666375270787058827220199340651108750139254471911028184933166696195649675789263286456676502212875145979102898219523924572521050334449094524428018419035532860247058653738701806150498558323116079668317865634879295570375916493363616688418522804095330959660455159086578899042140192752593670844125193121953032203406860716186036366445805106850741311332137903203490282357573101049119809124305750436150061336943369553884578436641323087842626250353607659267172752088525894238640839842181566961173129212514072607683037148997530118171540552597793181497792163520923177584089490668253712853829950506727806425496633632186695944747278430865923236241638204599730044911970595658857301786039143454037;
B[212]<=2560'd317753487534946304820906220664260045708312784502877904963354642874947490554836252843386770692744085491694874768517753901972865991619148624032181610235341486892060822392004691867298208151617104896210370391647846473919098822231475410435862679853341438281443853705467653491569992914567349669771492699747504412023112460360477523634902761612372843261253637354609188199166421747741948485795122558692683568783857652637450164263496253705758408166404820298688202809236807812493043802665378332636012939259469742303044739178864601335868193119264720972195590990561845927914557877338119839895674439177387077381564111170760317772541364399178174838837410822417107166227556969926465171634987017753874125380129716224751060816739579654904102660347239061654401342614652295661731470093145429;
B[213]<=2560'd317753487534946304844395089911488860701948910505839135531854074237262826465370810543843036022416109970361866605461582573962712924814271881684174045776611385924293830595331525657709007616393128147947770855880367852678853519140424961698500837061819335830840499020121043063404430259692638858884993290827005561124040341560053389342556181789480008259896073672471504696733239393693570720733817030399124434725310755423014180733197871515470086986551680138109395478358582772942297890468293767197678273983520194819649371091235199354911162065911217279975074978802495140700087949364259812697226013284987067922222016434046368640902959074457673110328236513497804023520497761890981511763175658880408604848924617523260721078430739531722108270930198061374312722455772210091685221787587925;
B[214]<=2560'd317753487528639321288993855542493329567894748470228013670436266589678419718534776473588637085289086982827995142077738900464698257640735745864555664780197548410393441233719560548993367631896476572559860120015579144487220626654717440702619225588949504570612655437231576996069497307528746824121177753348617126175180475093622912002720540758889327887859298131238284725783129240897720589582731239077295012938809831243027289808539520482194689388102331730517421580862278371915275120737713039722634653376812491855065870283411785482486923701505951466897098566378117731547153663876874002259683605613209240576439344145203708377333146425621626435351753167698286840467583118457800879582810726546080172668968534694646296782764009071457654749000831601335490309380737385472162991246234965;
B[215]<=2560'd317746435123088415608060873056233879647461691594630337918283153718068934005903215028873022541615844149216952068049476716587426842962640428744350090481921638557382243245852302310963186418855755890611586293023093860030391246335499133785978351685811734957196247375624818223345779058840459532067440259048802537476309521670914823340292631873092909862537441637579339507179979432541831889870716291661151057797961914512582649888485704887167419443189100884436636996870847891364823714420627974020418091490907525768538968346615324558706727767108419018223597642283775328512879705486623158028553623892065845886229068766285591452783632060055481028810873774258102137017673605114927235681335448517553684362437245033977397067714873397627887467163411531560990797812734669039782221053252949;
B[216]<=2560'd317746460949374809223695876718010647302645154426264453457498676725077972171348150998760707991291382951926540229882765458957271869987473630411777349444189417592718688631130869171533272935608604091185271952661239965566016053903248008326799016497767422341688876153923060034723397936967055761088766569055616624068649572910264616710797805077058394490828205768111883708195897138309442352967198269487801135511481987125824614877821062807851596971053250436490292132220458169261683630819471232205847607245067925189972294180455266234339856954185308135978222301066193834460216153551367576958486929428375572664872411093944829925973614913665671991175542678444245790043218795649964707002090949715097302200398622509751741799287302688136240907306231079390883804167748815285318085974971733;
B[217]<=2560'd317753487433640381438687106292655936377567726233049000725506697465330629285878245126730620841494811414987087637511811607461268417208125988862885696425782239821821339591102645794263777361205721240886932623527820421352164417639600600343241601409693702861732114672273603901328443822033740786285724392140325304030657348741942762412951256455345466168671937793711974333871216886367167972520423687009153808437821687974344719501276438244029382615199411344529106100076171099875400346631171755639177054285560841481429864287045065966801765768755266913524395965147375429639496408147168129729752716509544760128189497221791959925264534780801831810662012826704559048564320886642832565449897664577829247529093851259619992986527836379915941570236682779700292343894037444351750785325090133;
B[218]<=2560'd317753513361231062855010033258337593438400965091796374155645766186621910720505916099077251538865969733214346337012529509896737253669670955995792394299429917999217482767858669240911993472913157882052081684758776850220384655758754416259700741826598343460467106735188346002794115347354772178941812509621888203163242546677844173682098876684885345349012894666613329537630682102205734086808859855112356286987800078289985584342811021261167501777318977183328376033385372616179234558604905615528944639287157273211380385046266016261340030658635128244445482934907154778273816681029832032360335455667923357779719831706082305162206047042220723675498769441957126891310511083421532497164413549169273997823664233137665336300088760415285282393769243290670084618986787510809559636485817669;
B[219]<=2560'd317753900762203500791669405650300090499659171021887104730574228384353512586878366574029379147478782401654763411407986549920248501722363883466245803280078716703975684723812193587500809552776888396699485518073685469831444462346690059224996138197052731743673534470150148741722829448508426892653026251991798708380288505841335885996695992426582456469786400390297575850254764594208748954283229266311869195689826721405445461583018094255999341326331120193345774475696456225325555599517034524532907794035335404731128157283639130796688592795673435810319417834517169274234011027696634268527984861965018048909981961167283839433829327691839906592430258759757630146628099444753981954277272854616833972483905170063857543714782550548882912449842546143590155603221573964650682754318808405;
B[220]<=2560'd317753487534946304820906196956433620670857168425789794063270040846701652017769724453531738360291821491403685266793418234590373798842274890490015354196256493107038258628659750616329340587569398035916452406042317049750221389987875068870100122949188143992959802954019316534425107481668094507862735770599496940651878257344216767077520218264412520175262643907821597121546985174592520021836645682781160147905668402386747707610678889779520297790370737753240801623899821176466294142174757372550380526360018383350074593270641778213969426009836965700437136585156210392040961546371579196663565023611412529536877007032027653023579145894702389516287875532139891005487527527824744174475087977430962469893889769421305476778537248442376956757905328759546295387790426703248345191960429653;
B[221]<=2560'd344834750784320143710133060200862682141366950018189261976008896771490081605139322872044652538720941162129714263788340078943467626347391695668831841211004199228198216831955914674358447746275440463255261211047362541588134527965947295551169565742335177695787439158755400462799924022112292708231943344335545714512355047647639471190950235256766375101058015504387725290253517347390662815506416684021938844047397836738691788534263153717096240700517256892493128747581199666686256004603612469174259508045160409655966280175149346438835701936177423549190826629448620328692904368063135690240578403165317901872247691089434340458225927495765552830538915274704522461198120841639534762736470946170102737575450104511751138927469074366444866775596008975460328799874473170538745330556879701;
B[222]<=2560'd344947148605397338284308736871898818975764855390588230041483256077008911515121434374652215549535348699199024953969072804776178656964560633807509520476628144408208333719801872054585330453133932006885499837695410812427906788607256882258803195622893723792404335917607507716413041289873817644217983563942139753152203139629965185863875789171864983078479424693776054757184351965773829856618360700512605402943880402454187042556135668288932856405258659997100765163023000170747541700462992643717980153048861330760523430919156979918419827977178219436868061097298798823242388467161903232954801872060832649954698848537176104114590267906541114817429290539390020086223747798168093138909071335917359784505434248787928905274670269334474018498246793235544841651578372087874144026260492869;
B[223]<=2560'd317866298684192534876895883411111818309883010885907212717722667510842571941640277807161912600611137615071003936691053438512831634053375969953628531153461021878711957807163459323787615638592705684153971978463942886727180866335555453240287829797885937860176202281633575810962797570613106683708835554045326041083337132049319297208796994610532663370773026755959248854373683675944124401359492165331430455556684125161137047296212644510339895518308131724201405152306382436223818445098638417151597499745417268823367808207740728760565373156480130093314226234524386228135497618540423910759058182622294513152629926407095093451519631769830063428141612550814345227556453703874474461668772654815618436522417062733110011342193302617245203036884820270140890872142473394088955152114606901;
B[224]<=2560'd319558491749591100255814464918723839484564017355805357056730105981304556636412406966110438320042409095602766051221902135651701573072300300676005514654836507094204436978614204553154734719452631864329058275691203531673634832694856435778229140342350659555657954825280259620029808996689203565480743974315960103560310958796605413327916804998743531760317326893091246558438831718951158834574808803183707927088417022584829031553061192006043594857828634286459305138938379590640540768600905460654591017811463325143050013479926059468205787662404959884833735397012956970437195444609425961142861116928240036087407692721388760946485150761366693058899277891207422355242479491710383574364138321560506683069534973472967757586435990458569459573408675252119298538427618552561039459298333462;
B[225]<=2560'd319551880213967345106624731377263718891089371975152602183421110093948483774549082444430329020965382200792441636413191199689953789754433649128276574779808146189069199143072707462127380622230812914204221272597237136273578392728236113088957573260373179460942503897884219791461611010605492366137801602465655111031207508662039668389607548490269096322830217151792359350057613163865986212293403145582662353719396725449475190528530245135328632729798389768259172799320899408722323959919794416336681523430951365470618654760803972621075361086475287262561076271897435161512365716041557695852323553038046322540157248305844604063344869462803922242897923418933714425277298687666746255458696530717318317787601393548511607098601322898417941419964019716720909410973256521783597792383747109;
B[226]<=2560'd346640168219941423464477829955346034493020660772893565874061069997431982315691149280420370861846522151625845347123132853513944221517901208313429728005304722751265541952525663160756734001249940883927525913628241082094896861488891034830449874208485141000083846758760318865525908114811112509104950383241285712759577523580980489736443604398594081380813979248523129217675697091452837900881193273730553394309811283549261731141612089594893120304256774098313897586276121011462980191697559437179342197584019266330425212601301551996810527034323784775537056304523536864599271749640025215667488907766388799420949977732540009354478580223127313575439400028074433077175545052656926622879692650614322103684918693320233944249643506176712265836373877502741411118641971921943015401711748130;
B[227]<=2560'd346640140779067239244690912482129374509895551909489349523181250312541859976647720316090396308476776598563861433690269136018792627657727806734290383381061697943618874538505130320524471102850133194499444014313683238254146923703419649339128372561794051425893031272286800934026824450934277881741943526257143748193489505873318041827436443404171261916844712045195380131287349617290490416463390171695930950077739754977104289558349209216843282312384222685462912662100294322794051185199166827154828600208466690398626991445927630529156398997834876693874224899372054696169182213736166416470556859612302066626673864347984080062714731409128633670780323002002672663959764440771390990547890765887583820718115452770188656303304513232378036036210199525820524347802381959296103859323487009;
B[228]<=2560'd346640166605773995400577120175475351950240313698031666749471488739164795146366890767761068194522842541184046489410612626116054951748253519243129502205524781668783827490051340218437546688243042096719044542295920287582176722628571168992069516020655067868310742575843102444994260653411768095490577146796054307292569135322466209195070355796160993104790493615971755233870860345334836450059729129028596344464864065703262903411110766133458975679825616625319163213211766117152372555870826453938377130587122135579858418383319684296272277614564436502295722400168273569049397036852418947649362112787964783762193286858382413160409145459935379642945320283221377843823072602886502861014253282097173515758402236062488109953926212004440233157504179902816894205775963801181838184362164771;
B[229]<=2560'd346640581447224898058807793793072740507155726240344191738180217225941747177515652468349893351572172027521720550372284966593755404032109702131296086973305866797806934349559891642626190863114213543624547008952028738337542644164981248017768791913635724190550754190924978359727518731785572448039835051222694186272329942844251884613774661347598793205527710217811338463657724079442122321614682480345060505354948254166888973664307283888568679531064221514440762800554996073395370143653562556427412395651992980450795368639280192223022271444890352826801552586935644935197097797481528444391983912687346511206172644303682317668160105226032724571558421151765278821077628517298984466990380633467491105892351307131022080188625976048616053671916553717757331995905945036363101806966161955;
B[230]<=2560'd346746367631374050104535634545757098546493336573428238019009521758790159691176133945053408406139428924666421182125905512590384017277091603052695089134101520721689842267219940752740056286863479084275863744886598139197619916206297373613741972468308882747849330101309682794038826351451687196154868943617089792159743671404954984048050657856635876613420881642674347451842623231369989432504175004485631456545839564919794100041038250816920468758408474070121998194954039794772801852411863744161331447353024731098128933284535626046423404230969529607262219214399710955686145490004050603495939798160056168126411679929086836376459981076084538034527800523958384359154379013495161776647682393284471119698471368736628416779251418700280941747112521557885704434018090969799426140479439395;
B[231]<=2560'd348438560798050727214549818494268200602129020593151545603816495688678818942391565334955496041169708739326811574299255193776599156366353518892181859037612668069204103306547781247382186367387092528428296334747811452979639673957241733765491541039296591991520604922075717760850493551896591202388124473018852335316079313814206597687291070585322006442470566795636383242393378423810607267432671200411762530544290369329023551146946872261681136461372073066045980664797981020611260332399400079240966698653544616028508649454495264258699102308411181713960945850883443351549830849818210172062295574155895478487469560834508374324837169333016557512568009695271038187898685806414224362130837083656766272852025948170427899872506517875952676168420762014448390178763272299702945810184684578;
B[232]<=2560'd346746395173158431446363877493715713824764440913228823546006740621325900786032161230622558371788813326266536091235484637729409306425495493839010914757911587768214489993476875436272171477685123029214958415003379387980359829128234653650461901524404419139857941372375209024945350696093749786507121452861102796641256510494364716345817334460163458165320476066657741905229417802945178248391575008747601202842085296469830207398580562325691900322178075997058584810469053768899192277974733009602949375963454379542437533194218048429740864885162846077088655957087816711317988928435263064261016056718376972620325327411759137029058115285726819266262466423095006940207359834312585729916982967070090879025570186673776499064201535404490630261660533058534676849673169462511906554414195217;
B[233]<=2560'd375526848904936542061070959929113125243271667737286424106587184340816897287884321018682404583038688497474496600670968909641825473591671096277592919903791576646957258051225206793961829304774546844670120019493760386984052185708891484277362100407589682637653277717346496146810548544009824612270058248286372098989818877841497087570824039293966533758001788895373380840000353724977572619037934065362357427638447253421253658753731621358400572408364987610715172669099995748533554132734088022356704118114523695010730775159108430492949097120704774204569264780213042785462255677950249991769570534624251839000571528975950912203019908855245059323381839549820257636986015484887620478753041468212510139495200920463923975296883195987739186756469209095346691412697819916325456925506569474;
B[234]<=2560'd375526848904936542061070959929113125243271667737286424106587183217577097276830811409139238257516951203291836064484757142687559043215647500987580016606826223074385296081427298989594665763744279236783027958726943990402912178642325174589532731208525984819564109345152335012335878394360226019080044297850670145358207469182218174440562903255075764007569151464676304564970463757146673245500652823688967332522762833562655129110319034005267381757097741286180593749127498713123369124302337052545942414450924643879649283965274951085153889757604229128833714867817210069011448216889001148191084272576286519495915764844516352728058836625466942866043382304633793982580544540505187417160108750159532144584169608083703995976705410992343453129944346456269637545599960543138908589530302242;
B[235]<=2560'd375526848904936542061070959929113125243271667737286424106587166364608517810373892650432926272866024106750870103817540589983406331161243904371592544153885203362254178399033415398741013035459189054297657797071113162856239639124156268141609397695753260015939463661983524486981713203845592121057715876933663972241280925511187378916563770147155631379817585754988556812014989252272252655773197743984844620412475057748193472091797636094259717386247891300557827244828006293541380756025014660577372947972120992726507117743228521027438555951966555828850890500126186803637324429652710848663494882406763292734255124596271882108047191485457219589401028333542609753799829499042212989946071086947336727731420291073602387718125204162892796394846400439265576559996272283867269545747154273;
B[236]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832258886869673310431100258640998040429416015997903057993074754280482346248922696337973779821212970557860488402507349841757119310624957708119858621097214295903699702266843323291668067703625866008239076434578836714428849002314881897016297375674406521832111652826269318714133765465357524619520004863246920096353775303352978116474151411073838229168623502355668871801861853778853879917754565443318732874302237248606364074868640440437391894170010232245528501382430270194484291125693713961352356234866533908844761976061245276713073864109834761974279956871385728780356650982452811926552159169609177036279348983214491867954869500779488148941792958295716782705573386637481986143034129943946947096034349426;
B[237]<=2560'd375526848904936542061070959923644107705512731742303203823232049672469254136235936305915870408881441797364496215658123751459240287415337224147228511381156317510458263156382430335043416499600032328796514562688409386773118000187241906447279308219007635879059696510540250491020928841366234131277684148590469514739011458788449435271516909298095720567715508399966967826171071772121370420137597293145710387137432676231215976827986551157178045497404293598957515410928540181044170042767376950664001223214396101324404114478547168935944303722705205364757155664475383831758931719874228078907702730019990059568603086398582176786257646519023734965396344817625094540880840239711761682456860503125656536071314824241783066228392963407920817223610077560527725055278096461150975991519326788;
B[238]<=2560'd375526848904936542061065225155606153640862795991279131701118668999103513027127945150200232793292397927528232038559664546697083024715379447025610833725195491180412960697295406806542588213746075533204453409409289416994395075410361372166369086339266880301548227257275540919535136028230867464189756934782589101822709985485632424413213420652174975715815845539446486876661475292543572927512279327793077888241347237409218980310167769905459517662979893027429860390277394660564310217187923862229494771793989755901938163516799975844653310305844076760150781352546058475151102564731028546353355423401661733428628892044592273682879724453322148975736695956987686856026379378924062950071669979999805597867409874475930830492311653601957653538311886358197324473101043739270403823819183139;
B[239]<=2560'd375526848904936542037483836582080028866268975550228436299778143311619006558016560733946595097244295695416156657526104402214709960678569788449602372304373203126333876510934196553254711838007589491830867943358748854804954613856315752791597049006922004796781796669782237813716727368077278028832102545794743000001630000549333573315327361710252013912280721171458629306392416220604064234680630423037612808281985670038805103337069915463406462060173759553405885143820089126510373891156857038473137758536670074976556576094943061442034994280127504671619922439288081782851013128771167609395306862821696563868110113981168567389617052184183384375925360760197876921696784544971066848403709079032532802376980676143411379482208188612990335652455712739134067247236761346319464843621532706;
B[240]<=2560'd375526848904936542036015758365459711664380839805793990750324498497261492383932042403718780954331924348499398207725062316205806947845091146586758844827770456663936173677946673000297634828208998078025408202130556652138790226120548222543092999005849299534105518538254891891506103792761431433715839547615838998417869557273573012899169746383219983638363838790302774489161716313421525830713629022209992975503409723281290193676886105811699150673185171942895590379946744255356390829115594837123396886576833946252029788336239589330068406050250345470855792060279546281128700179951127996245069234916702187968585913441026860739964247079499391001733990364986967246608137925792689987753620678465189856828226377012420656518527727303538154520726069405516664144942866714236635253182649667;
B[241]<=2560'd375414037856996234986423279732991204290631047314142076851835903593959168892061348054767653219263854623092258318270815478844302380713898963758472236421186900519131395017076807677827932339621186557555041191414956319132589406271856179910708165228087578225461237246339849303415168704156143722981745160492301932475570833299141840480114631584124005958843565516990106423094263180850202069909591222872260967278060832913837534585473662290470843665226108173731370990224456827208800063007842871614343144617037560009490882510986016918077278331468463692462692265157034250034796927931413452162318204950757069705689309585123637256186341201046642149014697652737719134256730789705575260690623609243395531005385165469875703239261259749307805061870048713350524727889289896274518525566138418;
B[242]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614622124380461241603259487782026270908880245333760961523792132117959449857122259533857685058446761548919465169024989514712398533613874737171230756027686782001497455119413036999171814375630130917216007485386761298368565355964560149939384333140213185399858955652518080017576109400628748841091811875007553059424405750788299137498186145298696496119261213504572170792061612076173465158938218688011945827998939961827694843302689917888204100760676165003058633850918635557221192133479277743977019789042122989486603468771707245588399053983992643521599186490576843575486245128928077853974945123793535955357398998895981375000083298873077323319236299178965065714700789191681360555543257841747359176685987636;
B[243]<=2560'd346640168219941423440988578396104423301481539449802853021465093237677057481490341770169542899668185228165494510238214200130854131177838460475687306015035367302581079600765322852436566792766418560816994918393087691534223884020803199982925848298410194537915174998667607576025243539516726217358353394702121031339709976418577233019387387754705472310054085902973301808985870190293251893555346474593976776471973363285817903726620716917291433392816112257225333535405205742913322119456706253779968928693446902432705976891389746890320014454358571740892989342883845176236738217605792043928921910107960537427927507355999103058618143259751981595087276179784125322939923224811091800526526701827325696151978347535134670112836714329435787295946799484590760200082760292482796657516414546;
B[244]<=2560'd346640168219941423440988578396104423301481539449802853021465093237677057481494084737407752145437816989657727544201946775909660888584263196277420567322311011164378463993401962793826185909111462371734585381543380586674414099616499268701791345407287040475115265389760129862581422728466415151001055006297904993898482580698615278852753778953155158565306449599997916693967888872718978869601499333011149074474462848517136848327086498175332635657178277184185926054068223441740061943164970404985659234664811224060035235407884093120669914400469176896686048796862162218333022573761748118679281927866087477757562120067971689717400136283079203129708795272770957051368405849783996172385493499443533996399232137170389875884623401692458420412347154575679708126450816654680846838996861764;
B[245]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678120577262328507216558830889170960411062017429977315742325748140102296565952025269758298173451307609662457239316892253008357956010901981309524699231321763160493566363708552960276293053628135015390752986947499590559639591865261317392409283085498302946279738693600482909909014733131751870608170753874164531192886354650925846202453215730970720880816365767058057208832481392587033977868236681830004619803987516130463255629144290971988899528505084492175998247173591925748425906291541246246537153417582279824737649211701654168663196856271375622283284900307861262616414624800744047840508403763636941038741012085097204283949016927637999181065601336773443197801845846422576969705874674899962128059176266771014258;
B[246]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678120577202207092384122363244393354859957961174077426843592624528780686369552787049578794974109402036775105773813043744821634662209189267653718553731705964654562810821678943016508606357582083799046190438258552788687994192528359560124341806109868253723116081168981557012534267056869958271286763882624228395069932824276320587478336458435507674037621177037922400765509738578327790640205147240564064760742051369749899853093504070928023980478872049194337506716815986629614127046609084361477134512647139247143281478726708708526709682444494101306766994214382029972433547034246192811757956345122580340894204768552474729142511448521547327932311959783838528145699737517886535736074524467092041118187737513842794836;
B[247]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124761592792981936654258000149534298776743685578558186338270770453701531871653285071117251617746249766163187269480896490586979654411262479207146885212629187275377841838186899014085678872432916561406082151351011127897300916067600298782581716155711781773442425357061993699730005819895246546540230040069242322016611521857823063205158710768559288486147679000433080183290778126588907468705880405432679969570449514825594351140806768544565409836541008650073912939803704373779495978359642365401635024435202619793467931369448540726229480339158340161416992241526471061102377705669596167963251846797833454293875148428708187126114683746125798973339741540211452282505542159291193131949783683228303140262381098267685;
B[248]<=2560'd346640168213217361001767036793235861318926445428962888816742912050459026503596158548661284612785513517658078154462401016708088993077968046411266986956965313678782596179367223357261760837883817230148473737526577354354743838206805649231495288192107985194109683551779313713705952014269452336639905635892902974325001472710644921094990975472671831186968987508984941394431507230352258339580537987167578559388963728515609109121530752819159798696653834481098075808016215481114257534582292881365225694067015105343296202985360047266946053144374333989776715723144399881758059459757203514541696045641122191967643190563229681845406141858857695773397535983016582884540270138649386227094908362691808163081220957957641102438555463493320057647940461784835440956155123457887021429509395237;
B[249]<=2560'd317865885463189880523142295052122792400353607825920095277807794088524890073498937879676361192741804417124751480357271885740877786854255052162998501851799253588048610746728661866679453653984884113869048128385741261357074654699847841474589412644917014621635965867621651735990231193162707951876754619903434759833510070972851448402769311070411860655383490812714056193507150743070206046779788576981057465177208805553131077071978249225101122490774824372612953534868699475504184235115574103416361100293055480002342096773155242824749515577167341346870056575324036419616303014831786156586847748494267308821857434824969540656850248368245074767964419968040720609617301883729823062171760849264716019318076014323593265190843998433326073592875845126272191313593155176582894269085725250;
B[250]<=2560'd317753487541645736996250682737925379915482126612520921702187059209468758938248417646943767798981289366275724915521607092738893091407762582841677087600349068637708941448363728032058593069849282667554713097397839024174385243574972749767967322915827814580037218434005264284499344805618023991698059656713722655580511533035262379220135660027206763635511278973449569830753544691880832617924223734101092984451980751853594031348135803783683398989287785262397149703889607122002552548057907917048136242297733413647380709598243816151939255466621034393092976393908450998351766358886070394775018926117589332485335411631798336973967400577474954101953246418092901350284258409832572612322357762011704778116906836894055832246007914936478010205042723776554707441251789568355167622805136225;
B[251]<=2560'd317753487534946304820906196863095726923063743680768170062177437513702521606788544526213491805190418630894751109832841492482971257229186401292355738089994048471958939027254271005835556542869894541819889533395090256047242675813776787367718528410176160352136365820006748993607147186763980934980563035201831054132241731035430427953385944381740832085875699300926530189590820302802000955886418866472215723545216231572953335201088492093484381420480812231475664550452355884427481139358841575577066775600237689167817697673959422699419535835257323794456566939321174234799516207027228709591738490910447454826794140234328855197904935627019353291709774301103545727481240476779353674050571802207564572669125573222134027393505903564031147703407567893556013033388408832381712875025076486;
B[252]<=2560'd317753487534946304820906196863095721359696716807625409912653852119802880690799373662587476914451193911069090657235558802773175249536716861414030401232827051479331585043098328861983708387681547237162220619851243703499833848121001588698698574868815668521482947101516986040194711235476494607223389168897026312520117188451888660080942948598964476933847193012112477514110831317449827631881228070828024826140830603853786552729259967072351974694874307182301665652172643862167597573106044820819081941609452060278399706047989360874155534905970288641783805043858337945112575578335276244935972738192142270713437006592724408859899041340073713947213202372323753906831222748318179649938582446356837646786443572317099552213125468266466614686873166380263841452438106302684835788971139347;
B[253]<=2560'd317753487534946304820906196863437534955801364096919006860475322615284882130558772921061936531771964149498239087358683892985132801107621303565988932806907136315936699173659033249280240823133525981680933232940087509041547891055566455797844807416673505779392854715116470402391888025124742937549293780750202619379214148375914424589305097817440426180105730277795738536672105675963274704670683133631785658504056761466813609111437977329606558397407504527625875440324752505175979994586506902159899648295210591727643951373277279131092923532911878583671566720316863038683151208494081778475430661521035477474626301803758113383321636796426274786243456071670228526147787698173306613334872531942941227998871941547141404359749675999598734249090804297051970714035999596172368411639247872;
B[254]<=2560'd317753487534946304820906196863095721359611826482727362593271270814581373189530612006778407786640614623524036636879491731074137701951110001840110117449331969682376377265516321349822966292909452521695326789777601448257490522176055609980226556020868266577542436346567130628362255274296430370478115686313391509930761546868923177347200566064993635668563510257159380220150220888228154967782892758668736001409444437172794759340885018100168542483996487137043827867253232471291193409661721204373021540176521652893145623328210484829265326091996391503420564858043004714527430875472783061079327571449836737602205183568074671635355206976406741071551942751740347445908107920231573313804134206260225859575715318793706065700426868426779395989941618764418820403795334320840927449453692210;
B[255]<=2560'd317753487434060641755263935933895307868796531313059089930187144231763934164371817129561989796683938614790182166885878142471101065892971203068214657749223324431057810301013757059473716911923396574019963457614687666403249228370821482309789919522480709426397511804535509392089910967023842643245027209655869606386647736993820500381010236694956629021739611745064116360280182854979087744184978902509717441961488198015972670143276177261186774049359643195815100197226968018953729722957974679415620587972239133221594889776149852659779830205547207992227827872720124388949037416627106204230733155117632335097877434432192115065154479196743758535169274916679600063717368394324642621971564207604498073565344585229463518056587762707153876834736600178658413332786480041350741906269995795;
B[256]<=2560'd317753487534946202194898462619753233703360157226781801623213405266558199262983318982201916308312192467711884515274402954650849681600911788892671269558688947624160616311952300110787878275071936145524861655826653338256357640526119665185905788969294804522962848504610132575852147097616828638513821089138756932435131808761503298783044285502605188652555261599433508543090052083526733211585715261997246010881563831466811632626534942983262638043171104321295821273786910741196323249555350930986435395696934440547358885790853404719436966776449326313505140214513603159410946704190837071379559624151715991949353300647868849262584847548222386471275484133997817493437191740264518537299440681985551917497087308838049904723684748564328596292818141858676524833300023960721209169011613745;
B[257]<=2560'd315948069992134110306566171017952653200152872582352403335571963721639733422862072878105258022466719086022385607464785338101195530181815128585024054453450441709179915046548598042130341875904147094789919676476551520221686997657480973017669973429498865264785104111077684962399937920984427541982556652191421250309980204428879478003039184523832463844681795149441292882822751509662997531687372923241746954110908086029894591913370972622391570348866833074468104983018145722738572916322284374505950245374984185596212384689758108775964041093343165108415183998789318664379023217707120727705831129591313633122753354258571277059399344698016746526281015759229346405459611425321474695111043085386159041137295227812197289231133170963473805805481745413634068853962932749350753881127321715;
B[258]<=2560'd317640648938520543038119868084517517824557377420521907459635320501792548689885034053218025983056347544922876349951534495809463591875530969732852019603696663676028638305090009942927721402839944540731652706185809235227954561496081439588167072894643005750060354482095381311666890724525911088253798137661423101224216584636558871415788346058860322578747677624665432740880874587317731115799805246107256898797239582087323195967300578620997892272686846148027904891071193806772707979665270658617882956121089172954114990722200913647528594459238256269123052089577235850820278227095273675754221120869562235214321509549110168294967485052841179022246610653234673433979258832471549347132598639596593591711753683698953013598060624580883802102663538416720078741371317471182282849666605329;
B[259]<=2560'd317640648938520542638894370453404480048226440710511727196753897772337056549868125820559187826078180402939622526852819024378787780626670746720939668131716435308219781089605299173362043784022211890016275587635441865529936667090792723012192292540975421048673083144242408062303625554727345328194392727825270849929470542516724228321016288569852987190144505166444184223698476351320207893434286676576029036582667034321539991612328771221669418452915945744339424574316928277517662466884599393089299676198424297263580925506721499577278522839304187310615640230434718070432569993248133075022646706327015975422298499301802563301249948009389834180965739156232430267195176485274148743223822997859446598549161936338222599939804669292153057222965737361192387898302173394937701629474189329;
B[260]<=2560'd317640648938520542640362450157960744466411970214354718679991686109502669626095932683589427949689659253161371866911967538513882402716763941640675223694047219217752622437587855730411486761041105534912382521920247227322858488637361059342928780987344905929949643532059647168841269967307293714084409164966271752363475307778117107273646096179561744738958536682847222736869622733477339246749182134750883775996060587482986141409333594593836986849399331973222119788354941298463563690817123122948339654369826681736307203212505559414996842750401362289975679469082904844484324245074694362590931238748717255318162830402690066461153946404708471841232424932969141694696776648696993766201985573709599443256928337424998845944083537381391737262923463468468544309961916108539040237814284544;
B[261]<=2560'd317746435122669694684622212694024785303861446098327880176112366031032375778795317006913245828696099607160884624684899505231830267737235391468697234972848144148376248303854337497334648950681380644977968991447831884273811966555673463470213911254298498898607490126233912958956281381448451966960286257250506777727700329534336249118534417358775988563595062324776791249004042743676828993382016718337845579639882584018324163237636701085447851822498230420984829515945017806981288636609039660075112267526224750022982793358392158758896496890434669480302512039108785664283379328646956192580730984644776827127231742798101815903825897296764273129140273876442461833290667925479076168577594154596146024518992188020476071223495883978467591851379352872619392464056390611460882734107619586;
B[262]<=2560'd317753459986460849312560956725472569092506888800918249883062862634991083163969174093271217195096721335843334880969806623357156754529479641609411789761931153319318258634991674486683656301903345059137721112144552962039608367829453151261823566700707603283610218172830254166446365316343256110070804933214335255735180100948571636889518731204288686673401071910766731876641707256784688532844218416892718204366223312698731384503266573817377934971120121651026536422691090361723874596825748083791703571581706664109805182918569269998851316754917591363772215336432033750764649842442778637998101423852697728143810485193524996717534378924091172027051314314037948615651712901313980372391334116459344051555583171207093818831445929087759148091396139735624100005849230490243760530354444051;
B[263]<=2560'd317753459986460849312560956637990987047485562195439779218219900017315703987777361350898064867256965483236729602048058731730113008879076056412011633032633159317246611694014461795018754136283181353071922724564729801050891401036120747041598603959548158197031179645510987879763193018873934680232688260078707380685442739611357615812234783566352598227142944687225602343081362019965457761602687409365228438689952964482789351474279392916411941546689405777274795728180230226493357274175921571096872690886895724867278274697298143545555459123539941351034703310452349979329371413816018465127876979546135543276598703749636433085014000399067050595629629498253150843820459708698959814318972002007879906422816845123001066793849315102733820571602562998696870892886219671496049095098058002;
B[264]<=2560'd317753487534525948292349245794709938068249858466808087292372734227895761474912745898135216077055611002415837104828962115118744433188610474897626997064593823169306585898925531106887730188413709353089954064780979547499877691830050619940766871684166005525451645815778197329614794542465214946200545434754086186804680848326934576591804295242590237633243085912725574550973414825586983666680314280941971427209708624020303831655522382098316003232308610572729801830508922321858975062638718133613990481557864091301345777251531235502677349347441056339887165860646970423341797032257295623400782526491743440368301474768895949899530094990803500107915295633829514968362260614996947320577959015037480947063301858386023620820950218843253767139988907850271204377897525890533205784333202740;
B[265]<=2560'd317753487534920032537871387421663423500086247618536283839222068791894257653588148754663485809209020426233263820413083636101253994494812841258117961721460968507375335185209177797297582487991533302604905080050048954147067143934727940374627895903327492794619976395927464580170065104162939639647166888377222210324001161791925879851943714501209422854799571734830576928994329481439722313358953279883620668263759864751925410072612236653919443632103550715041939527270090426247205519427290971393015052946631228718079090989357874748899874564172709199758086362016020705753618783663600545403099882025371061945747425299286598980535824904037597675220417023634567597174654758557892878775610590983892911129561561724585958486328216339641475859017441964374170031467526155432170630492197431;
B[266]<=2560'd288979645446376941970361744943200146659999522019908206910638247492810100740838637370338268729188677087330656798637929021678140513235706014973759812029069409711592971367387808465447127931092489062694752313907268847624446285830897836673711123412120858947424263569100658654720867866223042708730378420998022025886042342827829266536545814963746888725749657401356415135536908967296217174234150112036986982377506376055219300730793233487905288182591325081499201897511315084913665882300485795404385126621583990756757442604016050773297334317389311892891185523089636851253787250434144163863594734439724758391586784324082065864951633260840872781368521044988165509227081054367259524566157964207550846326122444771054311393266226796502154398073457186355259705058960307448737094792917042;
B[267]<=2560'd288866806849977458483858624771883918446695681130237286540045596898709761482966975056288394160891480090463410409086245711880041422386743170415642274764497860817481281934374654262979126551741319786079972786087461784827060591061555919407263787168624956202032353540836595922501943326864180680812892046297314875485101782194377708813559786924305820215019302064383659118277112541453371223870974811430694782263009645931578054737766669351204783408077398910111070025336646132854594513644192341321596899725812023994952536759426757880512940663279683269103973959881976107062402834231850989340730088228753566455499011588223840785467330130803614928891858566154689988718303982543739709501644119916953332507308292813562535153268176764505705964703579565786456984762365349713187736209735716;
B[268]<=2560'd259980153713441625715192280146656348164599996474616019081929490646689327162569073469254301450525005956137870729411630231637117791948567878911898097014100217303164312660183367662770444908517390735257569010134985375858887701452046385940321416884065362629415008839259709034441916730449783723495757426038261345414938305972166297891714063625337560104529502103077235048308413264933588794635382190455526839960285941561047521964503493359339134252897595031067565389238109288238061959544920929130552000621764200942041974164213060858468643680010600114769383766807301647142889889749141744196470552291391395156710290472892205266391979829791626220269219128371265744056151951135535021869627987875042621422236707872206990578404854879850276257464329644252135538732357382213209350640705797;
B[269]<=2560'd259980126165376424109298767177864280144426185042439714215724752053711918711988823038828305599271269428203579734470458331702872858297478260082661441469393474001022944051984282568755502114514424877434360622529178520147997265948503179578801000242269185647900833540530496935316692594342910704381353868339700113648456034013296122846261891163609185128360983732719290222590732732034518092691645467336981095706128021511501684116217290369715576768741842489727430546313228250995454058457376275811547416137805894951257033811375145942491109039678145012796083697984210322382375139216451295066371340874240892476979712690171855283720542377430455113272753899181136870431210907312957287213714770287424056501166239955759907038936249981807910134786166907755905325898890386463450800963797250;
B[270]<=2560'd259980126164957709598431109480528522976581204176389254795563441565035817826931338618664392124133212584026236796659287452535988878703415654806503388700145241893115554280579567241610919995639880050880533018289753551938009545481786074441487136754248314826441005100224360756490886516135237018309122745417541907373350104384107151558505299980478149840639637932774267077888347627602619225000516347931746651514380885766413942714056239855867581978066393645868107720602045309979725091924103037777334902050907727053230517849335300209771384900260755633586873452307201383378908629571156007042400264727321811007717921802697677062364663611311791221079466341826934190509663112343475663606406262768955543112831184362644061140789609442469517421745580827622514659047338976529262277619389504;
B[271]<=2560'd259980126164956073994873034185690092983248946030463350693357838691612958441051328836841788657584786490717533226424112379133972763299860838236471488563311602748525007094227840998225382360134904686832881951917914218928921105396264308487979163139330391234804749014820699397178295344247931241375194128524285002533464311945704956164570845518108774451041485041521502278809590394652696540763488351274870783678694094638057351489442253662710132478479909460480940092961719020665735037888569948675613912553446728536087715234553449405550707007616147573529552668926317208690969704580749901333468381438995044340830171103888578751762598381230771214355500123035737177945579983684425360911232045763835852849839293650369188560679649517775921833579231682390608486110676164272680513841399040;
B[272]<=2560'd259980126164956170206853155514029587934616895873898364354811990626711331131052158964428370481388318118433893937909464498084430128493210363925700169671043284880409469945546266981927970355232722267633814682093530345175088222956725425070080053102197143530536911884143515275885117814778746794288566984716609681977036415366544049584639499912232977079908192658236882276823779475116632324622804080515745266285632906102107835313600530665198290214207875279265614574548262579609050088834101638240256282449951713585759625074581131759121074555666050081375154969642094753964309147820516092190827397422419081805083885543824632329594255286559081241735107460869610613246075412111206895106144123120398153836890024427982054374857713175343229929211028183829895158830908138897431325842215168;
B[273]<=2560'd259980126164956170206847420833495914820547020348726212822807264190675175790277465847679504984811791608511635586367190170538005986887603135161843274936980744967375952952811934737040793123090617924864697109154202775334160105094866109057623423245899205076014033209887130099440038993547330200651981277390392011003698660313532290335662449425160422174927987867143233078352148700015593246361599502434452505176110994569943935026678591133299570392566331304397463230727819952324471741948623895868231711027849080736289100359004653004971874584088514509659247554124557408227207096999122460822418533156645384463832742229979110533875833289820056073191083859285111728730501124557114737070950907868702654518018594025959195205189395068927861719310226246090722157368044346014003549101786145;
B[274]<=2560'd259980126164956073994873057986854417310138396197753029943385654956091821258853425432927861803567324959089846284047238692576625762355076965363395941799757801441000556862999797809798332948017222410245954266706392639349847287536744708707424059534442254094393925472518897140452094254843546396706035045936606743483131214071976138645393211654038033832309685666658284099464272615730616878656040156316842743987393563797137053066878354723191324374228050421362004497692511962645905681133348885065674352659008558387894693821421757169367405243615877179504899796006939714462879696877513864892965299435563702955857377201895019899316261486579178868542895594956631654298511974677254538949590963192738541366698740056296359643063334483713074700118707810056979806222507544511480369298893200;
B[275]<=2560'd259980126164956073994873416404387771879767763498718924179914044435435987811082233252787376235672593533905217409665704182379635889975193385881660184778961904201236497117048295849963621683012689289001650374302272993790314408452973477108800311365676977124138639756634974475658162082882831194582290826543350078866779119748773379729963895509337107858220418148910064768124673551453655771469722842197174123350614446760074602544962956868046742936030777878724529283508038782522081835110364142254400939947536724199300900174003416925636660085603311705747561638615276102241990832909705989888482768560489242641806488624259988982696347174304625108810565325963803065977313443483578508925750354462286665657974234363351518834031484115238495159842920763462020177577588735245247520168940640;
B[276]<=2560'd260092937219622078712983056172480110885186913041830297681687066764691229103699959871019440887329543248914928482219920815768014839993730613984524231882602500999002176630061301599508263083264832035420612470232752178719246358447538173955741754644179749881805646035317515385595994129567459588997629609675735605719760809339727556967298606639016686475332434340848694267788558734796399658256602763689593520352686616360053575218160633148515422605056178229304628365737131147591930703833569390760988130318311765313381578621119616941072396096185716775973963205532529764377991477183491318306794406359498705484141385698811022591500306290786083472248040540403907976443507030219044038212880948207541810496768453077173724811684252375412359319497936531847067698776776491085801510757470992;
B[277]<=2560'd288866806849951192614955415625360895613953233336898727562182412852525714902641054814026216516182792430517548265082125751717977624662277627134866922233445631902652942438028721398396469397680305840634534063190102589324432893493971521678501311218259204737815714120416390766169667264423916495622795667440620097600644174156529830698699829192951861421083069171036135894500643493472441482527676445204179873011320839893279535241723020218658947537864390061216447922077560537233217256034702925533784409385610453851222328474719633429250322030001598186275948718496421190549544599180562743635293539142949259443858219814224267701276883866290616324145945197259226061592327182494089441745685263294733160963809515421883585583989681051941582603098518813463646743535331749283544521391895376;
B[278]<=2560'd290672224392763381114578964175901481970939881190232139603399573560716973981338106464013211231137045496969994212207718179939639427800762007124333830448024633465594859214291636750237158104767421702597488431095694200327268323291451430664192274714090397666774983786449859332873228551605795513522552920007431513144197577004177773230600410105317843667617322417382930946415512105102705249204953355019820447634385979299096925306482739288523027092590782233354964768123091616844851086388976997347857899850440910475554232879589132402481644664803882275039678846180647008043835420217106147127160923039953232452806577566371501296284157612253274300852718498827585410781853707847076865990300784423193085047646391237994430722281010246461581049831895674162333474757556846988297704876194821;
B[279]<=2560'd317753487534946304820906196868929340066634276223634716905255145780776909679364960328608483517924459312074692188690964088776759290567131318327241465722876867435289462235418244624663542824719625723186667995182527045578898192552483143875733410173386853694083345118223364375487126753002149545584957962460846518977647399780734397124486382466318801168342874725174148487729458336743059851932152689271354019035519211200985445126126795974848775888861274846207330344212246224079499206530504147475114072391443252499250506356955771189448149264900794352331059558122771834987866048417287040277781078595559936933790130428293050658776020921083302548041185128218769032860031200110193334163851968339581509856762525229612601069310853293049767745787239286735436361939832114215075882812466688;
B[280]<=2560'd317753487534946304820906196868929340066634276223634716905255145780776909679364960328608483517924459312074692188690964088776759290567131318327241465722876867435289462235418244624663542824719625723186667971607344862000944512445037011847498094451764098803773510197305647386493805548129811935976402306517843613858446966056512719615342716959063443849667882784004123509082125042560032105097063045991356934863950369224972217543291943724398280603727004471444282188510069315834591044476322860867923554433690568529845116034788217711182793553707210338115266248778565344585613440524906265116284862774295606351355259534913167143613561720931857597570820524295245773872195401729103333775850295514418466259932738014075809025682897743954216714780321089653617535768852791131743749906243699;
B[281]<=2560'd317753928310713586540298462664295929299889208391024408555736939218561786004688350639338032633197773579088244755610302098701786443849174148961725784110667209816716310082271999654957951291618028835850553883881281945489965153134911362793105091560098096585570933053488678905742460211877363664200921839936662449056414479612522335570650244605896409881376619519704251701637747599877015012010653918531827489460329719059094566710859879384070221752965437194010537774639525451328462781394785862521023684554514929210866229068041954890539580685776240107831884727121461998238280586761465913532107640023868510748285574274412231685823938048737738506330585770436244823700569518588081474943538075466763073390081475988291307621926083554650328098870878084306002697017373620777302517774360875;
B[282]<=2560'd346640168219941423439422628391713984263886703685131535420443822611832605293037333574037244518787172703775968942732286651639363198996520056094789732631319330240838777887360463577840927552306084478136068263117900069369054983563132136956737393934329106134026571688066644906031380335181623018587968642600533409945063710476427440871124385707217012377501075567700001674975824023294806620316769763374931925913939898111832312189827625966718240063741537905418750462320996426506588565801821599782695274859803299925202479424087227951494752831457677702004270028094034319995835677308599377152937671078686950196256527157081787937237864013624703552937319638923724680287671928776348631462499712500464842366294963062226971376517690816888673834349004819565948713418750840367049745461834499;
B[283]<=2560'd346640168219941423440982461496531257694782913037625399236413697344452265115959338427353673822990720667709456007610797439275785516251183123645926678225799734802090037117328540162575567999985994372592813821206334863640163545790481358472597148663889714342565014457780067275451999339793385267121747458811582603295044260782181902415610072144762570657968365571780525325371920205391114688339355854183464382774139458752720667987704886010151594880972095853417055978717421171840798207933968909058328585340225752424783033958217829955301581159019745085788702299214308135291925634520081350589080965249423159753203710218961853293558970649706675185664760586643848738128852348622239625686007798795845351828997686766735321610103824074697369307187195090153892031344163369114513382953993568;
B[284]<=2560'd346640168219941423440988578395762609705371605950116401753755397320906330115331328812468852386497868685624766778922666786709881353568246333605622878032792873659343429094883184064956013034323219323755819050201102844867563707125677432883157647597667742964348484450226273075338668700261586353095426271219128986149406158602143599030554098052790764813931780368753178803596221189551130616536499591693990183518732567007962233470986668899580553109853273854755830141732373906956832042161917561388007397070944211277769507639723699826875282710183835788746902162017531213276422055838519602482695190468681112507180757064229433149017720913792438233894689142236943709788602881604920477548709989357791542016399599173856094942447415064997504468497554059086003157489412683246773099425903623;
B[285]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197362591554881626737867273962924929099675963525137915904091778949339104316394217713016843603161012374287360889466219408083750848241898797769930648045743045688749525373783608158308119784151720703111636031376670383939478583652322970557734487404089330385032090814126635783115460588062314504985543649541832471850787751101818687191248752137759357245262119242621515800739553994723763745103453538351256988045755637990575285824607511439477695053408861658072710610089665782839379731294171936184197313158421152689964330077542462004594933484066689598894281021960037161728;
B[286]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197019365148533380923415399582536168996432636888872647018924890449265517180842278172079195175177564219023604688307968133883547182986598235390410962638849613276383369464554996690600726690625958888063621426488205360857307952727879295589043663636094335509557576978151328542804877480804550043287128126456463886364415909023073166305848453548668900837022857861510841706481633672438188901520231856076096795305886257304483700498980040395647403812559147564816865900422282628884677909332841620615173837260693822715099451849768151191986993463027117038308062628083869484883;
B[287]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197019365148533380923396865922779648780827158177900795221967848453454095044652718310837480068906341835080797981119534969397998097201822062436691818130815719659428946912125200058318188757318161271213497263277666818431513922056198384100998589627928675559298921429490833833759859091091051251378766873333807556879764034746324119223566778838556125330665271742425432059204353359740318031927021163245927668891323102168336762730048359012805140679763234696372874268439444158818622254779211647364262039251705589127138790164461383717334120704462470224538983381369794081331;
B[288]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197341145121396147756073074618384712962353541362160115379758921011107620259795752909733521878946468545593690074329803821600848644772588571801200460873054173121945272103438669735448550600063702905837710934898054218254626575664706038185238229638692723675359721813658874286310746074688566395670291757670390136084846292270415057288177384623039544356628270953596698030985450138460918215067271619280992308508283332513552427057875712527701897800954437199123569818050044029174134720165811193804399082423322595795507514201293442967115911505054663821496187703989896762195;
B[289]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197341145140575417786714599088588459881198745802674115218212809520185255283991666562891630378244191811411741567859792796487826428493357602975774110696588719541770283403971034353807790413525065197270707038601780639559522928281651864165047083526968260332548569147714273205664037512803235394055129903564287178607991381183247203955755344790264580523563587829939980397009125105844560961057896178527173737017601890941056727495665530046658263942385482003104244962821572437168296781581575772921736363793776659038763412294922391915056753446105094139528264159425735053890;
B[290]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567090432925311266873429198564184566096113238979985496340959643469194952133656835746548316138577005497995757447624029654308311456576051934771169379826663669214958456134421510898623358404159205096585273386580881643479678445821050156363553394595049845864962427699643404045756369353647048344760331500762640750764696974867641798887922823301646396518837505786188359727360267637473236231269425144112677475650330472705062792495713522731141693158638161778052446667317006607003796799194948026066385698883875399815766067624520126243241569723175041437100823052760626742620624981840818713891;
B[291]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719361317906850676857186335228829570195375771814607004827685064761220419558855611127487821085602613746027010565808752893009244212356400015098187109763188538122064581577551681723477911437147567632007399946644908171260143712932904086865109060750256954187389964669495484615346655876665070728800098965185522993397113894827930072338236235353101005280220356432262028282837607759869857393558032689049195665062376136702228990564420366385418878855914905129624062963932643900283869960324640033615991511364553062140433911668266562788207455870012469273645617613168373360154839089381743201;
B[292]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355655711332078306453572195590646943291720107179993066068724984637541280959265064180088169580435896105017360440926786073362041534912615781448683346753256480856693681614299552195914362667828769168502589819044592880369407939574046603673720852225995410400087173038068091334293110258998506772447658063812953951482907861254841026745130712090255280097099269561971040529673781860699776711770747820339146312390095103883599887263345545596249258848963859255882948085046190661897272141970501529732208812963913353872487086947399099769424727190003754996787563425912929704816280863136336;
B[293]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988033723812451869009156094733522140718190100808646514905608457038366627437579074121054161720255725945152036117306675986884068016537369799582071908641823013201065431465822537161864492778441632426042511114336149725287116921658572547479176607075403372981756554799675872465308436121353182783497684392828491159133464155090449407436781484079974408751881368376933452404756439532623068281376398274312218228645143655777014419888014808480585474863871632472053983025309489201045201841507930735300784585636028045445723305539480368582042644124394833211744;
B[294]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988033723811342844742784020489969899972921540445613474233240690772195962718896772977547046863523033584789382928892767766850314628785929674404824344692635015135388053920364090043372953508031962942816478692681817232488391462858236316093160488243009646956388004164317028083265596224514403745006759953642476230649539774109110401360154605175670079745003529510390024660111326181405694828715331843304246953556836217601954457558701481908031807775139288973839231070076954169808451972976994233086393583915905330987382181445076540217655618851711720169620;
B[295]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567113522630407914624097528568898781818282409608550189385854914226322757036883144472999169736565565374177767311700895881826058055960241032737565718070602840518511249993430048883288844839401628995704996137111100247093717804718233705301091297772828572763196710172702223807710480668597771342115070222664303155947597686049990045383630627416672344578057258956178768399132881870867357832493131160636666325617778399339587073950719366133781685719814827886831011076685539247335550845226580094999253625183532842163693926507287183272171426947915689750088375673994486014372961287273117253667;
B[296]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988033723811342844676938225318322563983949762419353146375418041336479980914823331964498796548988979695926205626186669190805361543770292055247912831334056263807916268903556286990403116539378021661026464664009037191133942514672152337519459981276439366477255760944102021711328593899538394494688879996985840973108105023157249274400680990752629129135406146194466736650374459305348691251333539133824365787067414565893370582197011984981960840092054784787244686465907604014855246959090931463279634185814240356352333344738461102165609590011684071834640;
B[297]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361560783658706004732103664600641902542363614354181395244446888154755421268355708871753778087647534500447196635385152543943035721006511517283719605503739652108695175426456644964600192817048457967132518885274252790795059133437497404314402144815968255137856776960644583898048330473462768708341178880132399706986127033702672026717383626829536338836730706681906828056711754067859792134772375719104831641593604527677338648424059723702534308676709374591345222354276153144228513180428613578634103679665966716600404504119831680819700580213870619223729593097227321127126893659670989200661760;
B[298]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988032565457608061109689092121611278952783333352473830933268703877854987356195931216772786368020973601662204468982178485966163616183979992319212899039155925833747184486191129662370762517315788495734495413869557281528970448298193524963297280141848922494511046853993819237012027091717187763381776133755902794296058154620576389927442176484306688650685329487365172965461599922277689867759264837684299890746672735226613137922952041454279315886419437134296518293426067735129401650991652067058662147872596444867510887932290943267169333678927932688720;
B[299]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361472119191134877369619651720082072433661069698730235089954246520197486904000888303912417684165433164939353047149554433814553218754744984168673558277585283658366058778479369824793097472888332731472498722030014843811773032285889152482778224747501862128377284143164753762102419962396509620922735359843059256863829530129003807696518372266492201905732425800551317227598747286244718275662569052835658093432627271170267666524052995797656137074628056069543277033179598341376199038918974621865930559742851191644909924419812137541568310578926706107394255951904747761296545865782473961718306;
B[300]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361471748210099014912036036603426930469372213584700595561729178296067989915979080709075952327491666053434314810378149440013610511648122733910035992161340201941985899453457009173919721915735540252066399711494932561126142789474638477854623892319304822078569855136602618896228721631340144792659520190588165540119635389958662017085643689623762598112441871940883288245529036757506501907548011656460587503326307349929911813209373791173597276108298757602273733522362329300510952158097014037008769942295789883759166206031767110784886821633631361545302678783865084581152832364396967673283873;
B[301]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122815751525225115196377771817401757367386462545557131520677961447685129326677368151404776737059354397667643404877592809114649074442525575662981111239553066246250667941330975492914250537080996991535703616572387840285703802376212346012914613614871649680147836618826303580533098789011768007865678018960087464709126163338629517337402105292457125661347685383970824961738856426907963052918389158077549250887826069631673437388002077992143102017026415460631640531025746767244374721140549838208072983249781327026641768185848005457776935065685418940179073798400;
B[302]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361560783658706004732103664516866771136115692876234950417220619484370766225027487859616341239196425107187235702540821783357248581152717226859686311092110525413330905466511127920764159586261121626658642267230488709245235769380713499800405692267002702624978601424893633491566048866366946632190767071902917533615222837409809014404031244738303137786889182164041928233566223157298924763596218499336322892198803931583956625910957610352571773929706381150873364744087426744276789308405299256463760729518138411942769218244801587630204408060972203892236380767852932963066947678973560565795680;
B[303]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361560783658706004732103664516866771136044244596062906033682082908235903977857626100058876769565067129089828776698737264805814103992565373953941406450368175156327099048422447861590507062070007094951789836402892901584933122724462002760073283123522461521082138350714332404817085686391090032895411750075728280729315343797166470717099819676995435337186377414803993606541870382109135525092997983299438821011816694689345685553718008582662630045507702317602302293455912535560669663963950188088557173207995071106210038776706453322280845856794167114858295096250550409360056836327586137275204;
B[304]<=2560'd346640168219941423440988578396104423301476545977474942047666673634590095409136184463660586387126194780246636445516679603967610207560672873785916196666363008166769277468239815958546324920157064463275809525456367551085255673218288991056542706930780358153998691145864962239433537024176590794849114601394414961273582518788590237812900424314098644045747216037911053795972470637489915993458715780659665630785427358729580861737549040016196529181562310921552268696969699109413161167436128314880793760352994910246707195645703683596781662600625463578807210441384367489617548974468450550442831253184846810568135322109935191202192455973168279487299908313444567416785681821096634127638719451873323647619915869679719377414140818878546460044048181075329917483535130146821221300943950610;
B[305]<=2560'd346640168219941423440988578396104423301476233885454447611804272409397093574543782048959773067898893985244428267329366620751873840002172752499030843396787774798990026498646748665872362609697108394310587915809637182933929957618467092833318931116999413025187535756542447361583603182505421850593618100447626069436848537699991238859553453831410777508602466224608986322508470091390438126348238345385454579123149626474140860377789584109506605560713862235206204321695876113495570544903790791668233674975232706640862444146310011791439300757361247731279911049936261890847625214414467133763594149182408613276852780566012572806772566744882426227183614488692786453661177173973285397070344533017113730068274113416568398449667460472563848779849779093252784573659508191823754930306756786;
B[306]<=2560'd346640168219941423440988578396104423301476233885435917859629898776014542718662163974169951624181541902443423122670810929418712654957331650611398627065077062109327828315163968085058295367362701852356089860355057936862836421467850794459404923637988904120142502179043904925562410103945598319055838918758832398484075849311363765447621933487090547458033587801087019561886842998657534468881291716551304032785450875424149455326032636318754532593244841867509788394047640801814037676885238700905014253004490561843540767312913261196403048715014390758612535070888179909687563317568074997505683259729600054116549454076079042161881904177564144635418742264181085577238797739929362888863756746530018196927307834257500477520716457309882706192850308354758797682640146319985894696085915009;
B[307]<=2560'd346640168219941423440988578396104423301396649205842767723611819493854373822104010099445408180586885318458673093912730785476923093888963435168478451464348059109250797993301760824542428419595475719635686892365812945570017049961590265590113907814250719162107828945168729983219896928275918865678453227043657955167915547766764008851622427610672695766838077293918661834882596097545269939075241638473624495834837327353782998189253733416445362776014840040409657280523120832101861294012136795788102552296927645442299989202470473220308011547427936921082815015417259376541485657631717544431264029585063961338938012248319030149533980867092568572025203086483922197027632716756050283571843052944623886907587211775828858597193390174764954094570158513252629581885068038837731820733417813;
B[308]<=2560'd346640168219521066937486828891007452419661995294553834554343263970979204877566674004431222817267624088614193523866229107771663641699394886204303022911086858950399054712054270089686697782401570888860626141158726520363299680170394762978744419816718018015001165756910607262824732429972149902450198250171800200014175124136079597461831284781144630295994464889957238368783941544453523730119382841824038158361924595730736008150092369387180990529346588532695512372743940126513769814368385484476568819446594881925453656551491373048405033971786398038037997909650582708964284268563605654954235633954412824979880320429115776126638843442952534865062259994922665147855130375855545648564344791459991383354597568599291195092333588936944019885105690579152263627351293967984240166440338582;
B[309]<=2560'd346640168219521066937486828891007452418388640421083120239808296147893560470781439972598720736711895770266461054962436559098567128784388792957115218916868022914584338409332822952081567126488360933246101423450628970136321734326417988318303924012248881206349120721810242987680869224453238912744365321040200173257657219119724292562757546930784219863923073256901427597502804326738259990325304481012616531941412011285328414314945647997709497822282622642225351572402245977239553920265804666312994735933515254255226025815063241848740171809139791627720176815900253831562519585030031663187902627786264022839372931490296015568546813453032069037144739634440164924197116078659885798235476829678300766501674613732633074355049957095153283083700975344959111715589913177854266913977282582;
B[310]<=2560'd317753487534946304820906198356137509167880937792738419593881201049396137117862720919147420191031579819409021540807078298533830516174747661319350035741409823384720883255311605077732380988068437898163912476905733304362515587890645904925545223720790208117626145173187623913257168279933671294615311818488909499210010628059676860892876562935188343120114350507574542375921393833294115763255887512631391548840967592061515132680664244251878024378059526057127979086134092900220300458009127724495933017554948327459848559708036638209322549717168723799846284202733384793972992338026841891089028540998026089451479590274826368750761483326274079006919876176619199968688913526013572140337049006550727648883355720123273484335652539079434955602469271767161666939988813481459189495696527372;
B[311]<=2560'd317753487534946304820906198356137509167880937792738496499590909143089375243973557712914858414797008282643303056300045936901180062108771660033239134295520925397067246320131267745424130705747144599464653005281406660103303061045290446519820935260452357789498917292113822318721080400050271306597000641473773371163937411352194984604356667400243160120382429751157688449000563948601019205122257552488917679900184739614387216320151486782036256450958072279758167237786282164835457085714945120569891996443424862045189357233463786242213928123178938561524193897057293130924222723343745317016627432715997557978914459928547613061948937138241886078200471695577042861232179904104655219973099623832156619450996476547942577577030662221669056628038625048884059189664621453489213157420826627;
B[312]<=2560'd317753487534946304820906196863095721359691411162319286742949858890394108415278665140259409260106879799984137078447975278439948296524640158416172979440692254031328790661889818655007572683860927852732375037564532471543210805175835612471763013879223981972852844224093731834187908419199124840675928042190371093873093955829231759013865622220231390316553063246586072572632076109782875322950556360640175304206736804738280649748461258378292685769326486379794835388458186562256841334116822001424405107961019924785649011228442693928859575484544730607603120409537597555371535865130116860820266473150794798353785340275557927665112191698261147642067436238357436872083243642464398095078085938959850548104331890483011730484033441664584836481294942064620606714242349358945444857336173568;
B[313]<=2560'd317753487534946304820906196863095721359691411162319281936343002134539352237345174649307257866305351539473040538043324838102283940237970873673350236521254975182907198340719861905024505141583602191998927495188960745296500184896814224479192746182807573720570999867471351345819229151793616133602142352266560162741710522090871864461361893599945972495612391118775145150600010395578104227115147124579472082297329600022727007264975243275867219672370899508013852532960136623344368301784355534784749752485083610190169137750665217206882264331929146038706620361299772920517777869574430441028973422974499279743176224748427359718370426660230703108045230082564920563829105284004609622256231068040411935356495170723835665469070658470733821220975874714999193653004233958915747406194034816;
B[314]<=2560'd317753487534946304820906196863095721359691411162337811688586404473928929542049364674719962046925866062158345006912361807641648590285380535046300098290214365926248933854634450555042143128561353092978839462262967514988185461265498750412136506452484447112214135921674747613618810241039407254269078290079356060492190081029745766475895672509489061099490009755608968162364479604338848350450854769016463970423429195475607311625164058241276971137425773463121142629779542429871510756299682900166080740450785772396549146815276246630498436315854967833664395030073367782636732801220697269259626326081553557998490413133437110275707224057795117065128104156963238009614616466354160336556357598468899431551061706564337111764749713210116900346682734515825351248387607637901868895878273458;
B[315]<=2560'd317753487534946304820906196863095721359691411162319281936343002134554353030447196958756435477478828486417709489131245412842725395571445905669536450740998830845736507297197974926460774460928955251915402986280433702067083623286281857393283127465235485095425444191669856949079435817375733724230390758181737212437707425345895827536777267516136526689573209512901528558898563274774638833951658753781327015979237195649101754637897823033244784146827017595628758774540169649159292335450769911375954819272772565484031576809597547646997359305222515924789216583270394897640268937320141245155046284646104783484542554551072454524778964494221601556185132399464351944863347002218041354305113417749262251600112517024135292271693814632790984354746038446572392031309828083541734907922360161;
B[316]<=2560'd317753487534946304820906196863095721359691411162319359143570385691210437903831214442527082243226087252498428349983738811388816586924090578385145421950890884966004658377752863935981211471875025795196975970614364721968920466944714308844910251445802152123788797315528107047314002956132053142252846998952384352254595868999514823982215432998528034886796556398493057563935606114992810880478978986721056386920585268134442673600755084459524516371885240598266175748821240348588256393691803201048456646508230365008829234858411733580549702744322512491481422783441624726380463432665906122722253602585196646162220338994134187928818026318785430261533059529388663747569241525029138040719490393222294425777153941781211982198054657176257243836465378591911063212214068660119689021334029120;
B[317]<=2560'd346753005094586844653826697597391563598151235904907097363227980012941001124239606847938592268058878585857298796588960848610858188262093228490339484436098246439993522127358126573679451880958743945236707966628198317736393925715119433229087070690455613259520652125038012279235135046519542372751722698394883380935759048457509059258936530600204160388863753251521673012673035543347755619200069027790754867524427095642595881731575449198279609805323406555085842961747819686733575940879581236162129204546000106314606061181132407296386832039677308617446461854833135049224521873186429364532436798849807396335268766101386354142019638613092042423102397705834342871677256695787541784686847663460432509073133545950645320756967017491735412967158404386144245824332613406530428735353520131;
B[318]<=2560'd231093417931475595679102140442529344206006919365358596121294925400655587452840865083241317940322326643560833456576617428573562604815717013082492163434828768933257771512959445468244907764672998020647676366064855139036956061209739604127717276590098190872806053396042847365389542237537014132301271253675135907570995359627716883754346863108231834853893087650665672643048073514670476473218115450728627211397923809324511902873912530364138328534989805052991437794499170327543490783452689064711873596384016786069482858035837052764690456642728814753295582311589579063668653120855720238416095535743693112657851658939952865129897836411342967866165926524163588927378295696781029848993968938264082842617840761895250253170361098707596782358432303792701318048335949542774656188308205654;
B[319]<=2560'd259867287669442144511845552963585485560224362507544774272171196301984889656281358443266020446113497104946470155168342713810890102580836042027392181678883752798239196244989427099856354622506742720630149461627251811174181763413536364312057294706728530473344857952822686207977227976742682745185750752370103068627543993351278004238705767307367112014278329689949902565759825164472980466475446707523990584859027697715545148617954537456357365883623261557780814922193240270928055176932746976885752211491439276768536697567324855579550205610353666070333754718544885245443215474514537665961354933871925121228916415756813398496787171403460265799014880994583896716431548379883848409705362721607757381661917802188636239736412742001918974871258472713376593439418801258727437192520610384;
B[320]<=2560'd346640166498161082471717000794529672579508242939218004648311389288871180857044501804912631419446898317683142923536394151754308368700594813111993903628412523313298937902475599875639539400037587553728189659831804345794205813256671187704070980709845529374464181289282214844282313168508345851166126124449666918887809110938630931405865326718106316713081553555226872013642030241590359134486128736610088889755999675371800901366124169582526307232320216864439000934652196394459599436164080264816582759124433673427924522057408388292074967572893962292733507391388616930360267162528931578432167715713536184161924383371362030800325784290232097629697130675907374833473728643560722868932542966880927391591891018988367711670475739340368612014281047820778029429160379192554515271019733089;
B[321]<=2560'd316060906873505235576900002012374009654430029806836164883902325789641940985008568936362585226680291753146872962659636110852745830064426494560500201557492681022745045154315160785093182122340253665297814780498118716342831275220917123028994443684648727648013241632433607816491306545058813873955303001371719493524387239996243188426609986533047580977422264228971841332203427495894102902690901417039223209369178959623979959565663701148852856905648029554108233503159644719963444088012215932159724698459327359918179601534322497576069628594841179853790855927457462793739536367279855691393845301540576007967702761172173433240203613442483894395099924469696756024437412882578832276748823326753811714765341561983751008288231307474615719104083696467727955852686269682513806805342712584;
B[322]<=2560'd317753487534946202194800592138713702222860203769311019687932674225898274078150484777729149509836634348723979210629667441997355725378176949974953394673786798620188803274780146425670198966079184939429622090877987097928098654682177166796675779968343636688225185417417679737038879733532477427084830566429105681811199386440000306637485434141472092235197150054350452323880977991935128985880944152604401767722419764498252102098517347109985558518166989303087189791917424550564042704434891158923052275812690285012824759395986059632126390624197766270893545670627387223915077487756093525614558710573311041310009338831952220740670441431925926296381276246635087045930130344914996311809580193313251475412709730100724377445742612913969499498112883168162111603630806737202952365322313737;
B[323]<=2560'd317753487534946304820906196863095721359691411162299521692808698211844142165704747327457866260690525845810512854482285598332150893651466575461643165168172885286936290018955742748673360289773612238662816795482986251570056681338626225112436041683696748586560996323398173213980754654131109469608322263194036421471714857992264883696199827736077584647230694943935602065082677920414269004224011506288520373136358211018373051566981685740102726013533998078133903967200845683957712467523460760274895362811617300800482784686039508470279269298607503083335351305728667756925090581870290040554969397116458318812889261403833184964849126772799017647821679259113615400538754894219984063576437592157644365606336008712669414183973265117876186446013741874234745248986592897276820096355009024;
B[324]<=2560'd317753487534946304820906196863095721359606520837421234616955818919699407821542277576063890415250723739267907519043404134341220388916003493072607520587931836604232604177612489074669217564535600554636319881252071484653095007028167871902083870222809484691467307977868176561134659228640019569619750494415553674664427354701901757438189369495563301037831879437070554808386395170878399913291132339651349404153406958721516768505442505403114255194832200593686136949343709852599331368687082682835048920764731512081786809471123209327446216437040282757044412512599277710718263986035704258077598509334796523677323722737955957494944471257784321917338108529286638409433032290944981820850836365228025334584260737032230318635751072422169796877493419815936519839361963449839869614638040354;
B[325]<=2560'd317753487534946304819340246765367383011010734416601004832727433169148998644722141255619196684211293433400999317532303199999766015281105126695530202733684075604115973730634790684988330577008530827521005762088171090838800041863350391726772437668961367661179723107836496469381390502396553409723935971996408197474005114412782897669721324891968886899801130785323508315943329596306950583767950411954719353217819911428214703289767205738633659555041695742506199557723362650573131204367405898751719957145069622968527146211586051184908412924522510745702019323828125881311750515017693837336308901320933907636166818089362515812601031407589794891845102932586661521980216518751927380206215904172313921016471389310749843881248442845718095645789788374556521166570136986076397933609421251;
B[326]<=2560'd317753487534946304820906196770099635644715503680958773701458687331100384401745602052369610171522703377693847481147548436363462179474006518011806371627714621130231804135740790535951467124870270722179543340259139781983623606815201358724096997680135722110395925179107302603812335473348090824301464679160714904018122806219084184394485341915287490049031400994358928505045094433581712438733620094603853987436240301877771714530526859688315749652949641890493580554656236636513258626921757602522692543284974864587717523993535531781104199262621905011434025885646081254092578822037767957184834389121040445504707660432684527689567188388550389024994303275434959421903445599305151923154217787890208509749489203910345987660969135760053652600777615369548080874967302829355271617498843044;
B[327]<=2560'd346640168213215821585127764456826877489414210721824209849586109835455313546501680703169052663209646119895333878137546346647805130801090475564189204803553430591592770859444654007306586213979687320490848680657460830051961619505754115776634389734804572056413714584981072644570540096402927243219089231375709581330985531285024095629726941650346124815461439308016201634835203295236228335999987742160408286635219706831373254442746404763337087919048592636696238581748503195464988928799870322422455601539012408003692190037668616756043208441296550463861958725893004081296028396150006920022106381606193361149505399911636334636142738456530639149309998517601228763258806680894748368684095808679751501729342892752839245907391145452562297632952389415109202359956706419712781976850177108;
B[328]<=2560'd231086420723781065643201911444655533564470654863477574985537838353957045725937738658815310599045626852227729000917899369618059868742479373791775602494602042549365542783211048644963533242978644570001898606588875098410875919024959967876170108530263189830985331062482995470278099260064878453689358331020383903370718493350084909021430433360782889284327605992687442152758372753164985907766558214216717151736738239377564326244172719722795245731407247186217024528052245010418215613686013774220768494468823165246551929606780416759157697285795025531993053385468394198428751548421432149195825437196989457406198233141188495868498889967772329010402968689815094527663799861982587024677517758661834606785164574481966609348952991557979146462090932278689759734196489440984693910712390976;
B[329]<=2560'd288753527585369407195769726124550542439999628249837264713404757724042527558586706768271305316842535069601800923827830416680784834497829935771821498716589242418749937517994671403256840367607801817666072335039899222612685502614376622259733996024803498871005444980781016893382399007732680595998303526918734340398862378337657355294608028786069605754784878000065825838688187583780231826917819133792872176149976490813075819631801953464574298462537503633542404212466917452539642780070099739929840249503509620229742596917118676798445895951380023858024245724596780562475915550111835209735783443793531985601698439941046518619089603478077626900350635510654402463832926344451534092960369246236660752507851890122306905407633280080761837284178593611145203193946774499134517004481070144;
B[330]<=2560'd290679275083259650281787114505612290569079038576859906521698813939167426988689902381115682157174849164641686544129393642409252505831402999812323476107178095174356122171327338987297624107374689130460143520532470060292729398485002904308385374948057648354832199930145654005082662896407661949336112879995697324829711196087299696578036371095397789367998718526161235233636342052956600819473080793123411461500724917050292567957791222865861992292536503240327724027824081962632793393419746881111905316450656715525190935835543805143658383279102634537342898150572585538373760624913728138688566223528519978775296599018911771069379178593321256163949736848961321276085379968133797340411773074922794773282301320896982013556600597870488488164223709451870384718677038523219045811080421655;
B[331]<=2560'd204125461810830363726467229145894952856291385198917209030715662464308586860361016220423983644386079737760982832182884909367068519391258345758515773239287004638903498382513387070655136805792909986483480584047668137786569324431281254677473187128846801129585781064321840686623334238687451964253646245654002265388099908430659705981110332494215593869230522306436173031853358777886860999313545491784475581434391495480523531495759163700555373121047737555108731877922983745457192493349792671704247672055009652889831518162440118341704061761172716244183070608131867491965149265273823812128440286080211305995428465954437625351013242433359043711946445385335657879516522080749484654106553674196279977219909919407926058919896818272980607899888049773481181169691106252811139356918710594;
B[332]<=2560'd258174710451561757228305814672544198989774941598061420117678239462066502414607223486599620771967923930413876905895402524554887156195295200326142642401596048847949608112538986346481743393889050781301588506241138393747020705603305134340800792523040053959644601255270111541157082677092446628386074039595328771320738954870438928716115877395761678493696043980644613473604071597469062933351462180261651878361541728731437204470043610894402118980988020430991327147830422078917148579206807938175472698064960586593802032020859443331964286768630876179310305149996772648881318590005706429155240444957656519342323773171022201873251437176346845991085872542928589920948592116783428077502155855119929614292115911206579389936150766650782780228327728411413260511180719224737608827121186596;
B[333]<=2560'd231093445473657249464126085919728956506363447855719606176333774641554059281114916530009899827836766136798505119197077930797165863243874384568634479812999564012073947603803268357140926305631703427008953523111049889578600862721304953738722077059467403261324465282835658903743632398906498163549640938361575997140841938363654292388287211523022730255751517309139185679543290740200883595038780077087071037193357396731867893299324685231370554156966950663458292771740226981877539945576587708124402100343823487458642302642242029728309907380876077662282152065372209933053324835337495368030928896948508800293913933293553306592182809782980485838945751333751587208232297061183807701350833344534182066375780488988790859732895406533165464100555137682534310723207484940002228222931661671;
B[334]<=2560'd231206282354606370198558490021580844954873209302937098685159385930698115721620017818407014904027675990207051251359470369028149957125090745648965183314068125917614895248559831148161557151802170792522951555414181014093840975291480260955720343222586739693990438463636586295002152525651743314816019547801712992793531194880980550102150600068105323640593539811218472379283904992479149836931458661326488448931736041778292620382657004672656164425286999112045027151643116854701894575539477340334439674354347141137900413472049134866698809486790366011412996570313949132144728597437789932640529113382263959358735150489901901665105661010802350663526074165571009305494317274034463843023224037894299453368824347865329955755883624226824962672611201359421297373039930626178851329284846178;
B[335]<=2560'd287061389300832008156039550176997572852029856850443528706494468340284052229061628375803826150440325514823949974968303905408899783413429293201898188948312288894467045836633529166220819949818312212828509139507614842392237194046171396995178698476395546568556709118294546890667837257125305805491290435972112048409259574632429935451392186819478473106728857896016300933253609603401829309347727461793922430099412886284420765696448361488988005943913628635704078989717579712368108002662117687388541834420933159058379430220765506474030497618022134284438142130954570830433927495778215155929595646516035248162271961297045617398607573726483589745920533699372426100406164262950803928928392282403134614447555362181129074478848926910803164656537067649980449974655080584166420538231235876;
B[336]<=2560'd288860193491661523228792500288233408531859295598040101771935743480078500731298220010234134712626200507078291221330804695817930480722579336286960533229644454512855191480032166828956304796839829419011604325408541914203170265521258291323367681810620223558691029023745730650373487350414559021943493059827476161571920309448700915870550510853540648872187235140618514367124057832583857129939130966549710306875792895546578098514032882134844945170926315191497801394766141186308273344192830589191756863684379147096343700448855446940972154735286273019687022981395739763280257545197666118543730133475113027498376553772834001774407774390488252606407208755573763284495473576838891846092036804843341999319217363672838853839634009751968582252496915010221559411562965858346160659439625824;
B[337]<=2560'd317634035580204607383632505276021373275503309057204659250797128361278518186462414132590675455649182145726199538026822892249212744534931761680608654339046049709261824511863654422703208161488961350544137247339564207730506356811197106741052064552707392541901493556156544839607043972844148061559936533616144258588594861087647837197029912031324334845401049699076989156100002660409044391606535327652779092729960885322784818559918182458283302065323163056002839884945840247607927657021850939085176825119805408357291141838925130746239408040905403327271388764024865137065085235236212840057925089060471664481192506875967007429269490726526143339085430432069527654121592579284516429307829101373666151643720501609302020355936989071701743446795812998879497347520923530605462974994284672;
B[338]<=2560'd288866805134896447062259978217194850437037170880399510225429190514792428114854935947356246721093008799799833095612591381874646592090798252193144500047157790935849499689422859223152270068269136090562870353368970587090771624026693510063785457073460011217352943045801603372826628291657414760765382079400076758860469470652764109859435552151614011045053810321657131542851142232190368253035793461926294171265774882545331945089807825921469401830089926833329371760532223595152214326888080483491193253868312523045677770804151871118755637823122800232671893994352026781734686413743317216105761155462913912120817932499145653985095115339290249652213791074456693196467020524650507809200798015727578871152159593459540303030051152003779091621728413995035505677665749065392127110040743976;
B[339]<=2560'd317640648830935543586196610443773827370044712068348897522578383429216518829957987281322762483651304511733308987153121919749484895319256993278167665771530552181301343280042580046288563755402596797176816768799570270469452193965128572232202209952652828661090371912911607659836118660744433279339756614095290232638637567085859003819893832984191232215692903248042072052653338817204328729604098111556747644054345669174461173021662173597214162158240768931641768971144168274623721211516004896254896867957993778410238490434302077701394630117543114718989420406937581173219896187792278088993100420314557997346689589061501590445920884381188512226837460708566923986684317522339550629038733458999149361207255420539481510363958149893092992781863524568165690012014414950561594765405848152;
B[340]<=2560'd261785104747941177727001333646884974969923880932807337941654690738262645471122767058599901613201724551190872382731961116902463832984852375982106262227414666840055875434983360387251336292944897479049304489045470833300213005277947949453528311336753698562934894996699562699258250639920129634183944070514468762419798544094929999253542008794207299873767287589777813414204289273064806216804422802731921925988895999670808968542248532107505306515395644331537513441781560005887371787779027313230206891067660423569515507384079596458668117570660102039656060157505327811800428786023158258423510317457997100283464679784655344210225097714136223690074377391617273225056529829180751502254629726757328409041394207307954608620734603451126964468795642380802183568411998489660672396795148292;
B[341]<=2560'd344715300444194144340699792701463869963154267545303241411011084673362581617198450098066682680972075793618550630987563915526478280530192325497881754868641494767650551626551087078302041039351657002486549200492006833407022872748225258345802851551215710135117007908927662639135331804571893480910812126999951191867815831769544603064361628669492352649023888222967747146145973905504301197837531104203808864306589231284988242356423665024772314709790226984752621377503021150281206875751200116101057493079912148788783243250159102123073503224672449023738589989588620984708388971970382570773620535380903526272462927185652394704420503788657600318105422148494177162552177905193574287826191262304210873771102040093558471070094652150364434172512605082055002713804393023422338491920045859;
B[342]<=2560'd262010311908211026393804604341950848078332782968288416747299161141317293073905725124888787232878492153259138163461128341225893138176843058426540945104599255505873370259980078377080291197970329318109525361555664732497390166549828126107227722044731058419857290795050876469691095495711057594358888528108469834746828114408450341223123719066686913503386687861252812652670022287008328622293277111745669251196799955891891153202041721808946547400857020497931504481491871018768693131022778464804273203710243012899528561863324911564203340333895844629637686242249476534074555953827293313040729161449482358413315555720962063455266271914616959285213692528002727457967221554055989543296349047015092088423394535848403647164754032814752003153867242337235146208595179177345138686012004912;
B[343]<=2560'd29037009017182740703509297361366423011974600620441062791458802183455453104411743774036747849093284890588194310662106983594389900256866341018657900354111067030663935050575985476005216050372265787185083999252814416578862309231665642044643813379656902865863345710903082328682421360084544128029840873177738272779183934878894816959033485161805186180365711002322858934557078780039125068289514674063176860361521039750503710328895601250846505144705566906345172785743915392707131959395847708680000943012523331264357533508318691329264158322321320573512282072962067407935169683679964295859008498284760631975480434529342293632163672242051141590044644103474237721739701614703099509910031059574867458027128228554393498007690607599577960195554132684591810151980108211451422273360131939;
B[344]<=2560'd27088437478056201010721536992932335213657572890714425110168654032825378907264473943406682712105372744828226782796188145634359152910325854397702900976563563876605755766162027110574900914363577861488486758589580574810127729574545699347261096629629309234162763080627327042842205779163877013163329745475566875449854958354979151462175923437129349535233523050403989720178344469025987149533657418025651228029397209839606352146280952384315059582896785907113965418532120831870140374810025682129851334655679220972108786087459938490515887645160680306364354192578621293370280114717570101433854989442180215058949395357351612781660173654354661803381696084741547932453115219279958990615915305442066419717199005645964733722764662186049431667080014519335765934183735536326798523640463426;
B[345]<=2560'd1798813627411595857540039797543963750891463348939783533457219736036182630540355015840595650331306945483720911439864962863106640480321244616639435086515846700590839536541859954846389050764629859152296556623525398944595476243802367914413500545874307582238038052161386702418800330608937872282414321122834551662590074276730599921610822501271194715693026031500483211195732095660184155245551320957868852598062931061535703897051355614279663082400547890611754656720082471104665319446724428853422743429398082374350279872113807113040690763355234238172348667070454659205061594997884706418831346780319104826183394243942106821267372404044709747291745970115767219530588435340158656374821751739390147268792777572975492715688673000263525876962592457809583842324513840487179923092426757;
B[346]<=2560'd27081322523427676400002663267795189050822784415616359460662730894948581425511486235990469867444091979972767774034683308101990508387897131353524198244900696324054908194347487406569479698551860104715752205181960874031007449018161021759247926613800014089903839682468791107891802640625382391724727367149837708680601259022490647447495421737819858945964038715981603139223396796146392007421679819872414882933934818143463441215721339941530440623986188981733802901573108941330642699445186182247152428375342544412620788320225380779795129900807971585306860996877595852930948106430215238012824129165052983794450280706416023289522935166544799848014629374713727814346520357839562687488338494424744288779127468833960944321670887600819837335915588927982891828016455010531552229019747696;
B[347]<=2560'd112432989393351520276984298050539606857820153986027338401474401490387473680250754027015207966420261568216670099183547550011897066373421700333611268936288209825414799987545386524372232904281930485778654873969504237543806584032398889378165292902427063927662134196460413048847923533187753399668277811787526634118988145192361496726259073425116004071607174492480362663889574767003831863817434786892590903906286270931523809743662672465312894230316804473899991997850009470535020231875348438353333006682910639504103917265290684065039454853522486268301966046959040855483372347134312413435184655081327924260166341264123411694858792899032986040559027164343657876442003474055786631696232256429117629670258201342151880054135160870522259200943020667656618690495228974977455290845760;
B[348]<=2560'd422670592882260642076838129933010681320207337220622153050654309385940456044017979282218045469475024078931608680478753016444271354050306823822254809443448722591010014918721930263380470756803919686096189712779248674913592938658357959970200135407606010454384659557038197847064094915222766036363818680227281850189933261804458847529885874058819739274452069496178285588017982515919729993274435334096766217267149106295497863540565223689088890936501667320962520421961326503336673831378691613237024103221385318522414611111950803375720304011885812018874368781463882293819811622502915582398850358201041172460866519883947489607347917504983689375812453354594446953003512542832958478801435274257713792480375938354664911962722441163971214787371086705279926016373058508117861466421;
B[349]<=2560'd1693032292495350832233695645547157125036511595982662141616850039170127957571877366586842718353752883724914786459458356797773179156721991369789070834053782145800887973365139181634235949228409055656712847538151349065529547248492871734182721043909326463832486757775356020466884637379560169163426747362382124534411039744053907208186221884255776987638185066454460216364176416694804293231953772128661793640298221284269097611961055662945359124593806854948077034182601906253997128850072372248234005553333635449250424674320317751453158796576103091743445218183027188153010455250486312664166780685280071707766804553309062243286380983923818750591101903136184597125445878236299465073129099661988430242565225820664029283827592552681516212559275391259491427463191344858758464959176710;
B[350]<=2560'd3171203279955923418714505557678250280104221256252711347872709313901617127792131723679072039620664942536233874947983486645921330704839116216901702148264369794568099001711484794225974222933705518833390138470176896476643902383617210439666113979922069044807913371460964443122453608576696146074282777200617469295758758533461808718022446005126127115528204590430601394181718463131723255149790268642860590057204707564548866022067943940635593385152506135716378673298687589904801361689437499798850673394830812419946714932513012288894200340985313638506355150446688490795810372952953869245188657478806413948979953082757277874330268011561060251822282829600056617090790747592481093132598019109432401166728666952160903518077502916015061698993899363224982362130597104399969072222724;
B[351]<=2560'd12773995960922336413698189767639283010365339662022546979462191390926870083701462263754303266016630061615045193180019509962751254360081593285415300495100926087602710753113694473853814262018107574514168882005852640590513899083081644360262044080963223924208488245279315477840794682104604758289254854001755346611415528058467719833190283321571444022361367793021221488676340201143872800026292269483411609845949958185309232745010881984726436652859662934436165456446218358834759593363777501272179907709405353456276335327775691382280470599774955761848078104439515225783218518237517151510580951382573249629983349642466140062083453912892294425619884049977399837269273392301467630870622314552450296650318197077016879724235660219096386324134196040492529781874248097520841120645190;
B[352]<=2560'd4020457981730102801956177112418806336012340394412192933511336889402879446521610640533832448412683166151689821654099731161729649686428187730115517884952415503790638285524171210313611114419326239819597849075979471538008889796452313780836641025527019204048127871541090368739562482876907887613861476957290809575375058315886444122488670201622460227721003778288106140301233191434445100336516149733459637478748786738930664144724720720666975201480828317813958643169132511015066069054026475681658852478649178122599156363201885375626696305418288759585627270059408518155310544593019127146764440869858579544236537662896658644045434490354498847668822276669602099548605499173695572105231643258898264256309167464641708025955265549383158036144389153310789510551104505610524023595827;
B[353]<=2560'd4433584377995874312324054983020067281194460802350845586497927891694663756055454985838459886323984529542359178928101557758817759532272678324778375331830256147108693809520075286110466657069569709220164613814037543507662016125037334903322341854772574058772629894394047423001328937158686551691473896784855994321092338813610872346743908275968716812045463248139421686208443804095859304412620093329008160775405103381341875578649076324134665506490748984931294139350338444140752499520403837238417313225161911861717621850062523831689485072114787517528784322379271099590080540379210970029234719852128198877846416611046233712649143683788964173619416035702327706062127902624191648898884798045440978014967383875881410313675634897007337116682974968283374995523308841651319304556800;
B[354]<=2560'd11071054291864590120385783856394281804407857551243123318953159957539993916012669229378491089168258617905922410601591202282999327379986620486810421950743230048073138617562007056859321604911465042979228858245039182069801884950271281212418665491725005079081058612001277610026473846590149951838506200873299438027334345732428544787753747795034581736895073294314327587382407095571085535593432152977079965984383861086133941353984039397720946885804017560960540322231586789378777502447609228175399651496191035177546259043322917504780885767185786771185531926101730693126437257257025977356347296159952025214514992247051468602778706549101133370232159732083582437014691692626048015336817125897790082207053337777254370549670374648904586803292690575005914433277596755892449403101205;
B[355]<=2560'd11071155177431819616665738749868841346168094944602547359664078199167782391661229543186391760905238687324277668471331266952708527176986686977699598477069187119694603426650159779705329743749244425808499721885932977086953081193707160510925179413028990578470070369186877118417822723285894024334517863909712633286499109923772485881646272786215129659929788615080221924659504433986137353183181914784503971176310004107242517969571356700115459871575758822173274889643779814149854436770978902281513267707507370300206360127535300580489412555992240319423692352578612514051589433427831194631155052913572154573656833564117849701359388594033851540464685415568344970673572050571030940988213101063248595196496512983390974596390223301465873658467838004100184727495542540306599887520820;
B[356]<=2560'd11045328472419530722711103601402340070018919999523941448117835433636110000074561052525481086455315268450011203741952650469816874709257075152167692602786114213560037891085543715655574433925880683254214794591226607905007768706736699934909433867021667383091307323376389396141080706711083905397701004356157174628316946495490825537451960051202305036307813524681087212812673057271378480301881330550487588213342209917543798477218218524479396882594469561767392715264184592417096030804112379566791314503457683542350749964339754964940843745993865062265391326965444736383328206015050959418766029591353746429974612639831945661618304786381489016603097947578785981620726777291870006617453794911802313716993936312526141074042252039008824891095404253135196054968242218094804153141008;
B[357]<=2560'd123882203144010400490393439838201321644092535469098744338895630453175621773170970191991788521382359888686382879012334447200744801738777513762612482137680110493835967447039130081818801607191970110926153314140699393491649259743730764865712994129187339494402211547506081866925723363085166809277479866862538967001209225173147315036205645441546492207183955411634889426336131586537722639306291283216154586182907042913575309357448611038130277821721128692031567913493418987267694174429906410553251183973252702239904139990355491134509107644524298132767565187321427041997617123528002246739671353018632865697292903388923101873254187453951813129410517037296373972377837533641138865931739692407138205175242376327602976136790706977372378108441300412192841914987745631797366783750912;
B[358]<=2560'd1816461149530437117425149070977861590030730833980996585509258444762524297583600639042449601316448533430350327324683268349570667152611238374630844197722742817127391020268420417131181593943435767911348417399764004500990118064863652207624756175523539393670366953080405385867943484833438089396890160040235756259108807283446596162077469808441364572307084034453894295778109565244976246097740376654094999654339767358980347894310453523779219185091468908066792457153747843858904838871344413541927964948999755780997932086508172811802767901514438160088478939893159613836359300486167658824295471292424163865741133967356021412081267171524447219629246015096262214401952962216000872361588783293917460902955424547232638202360000593983493394049509542933202856509443545833830437539086339;
B[359]<=2560'd18096018994755728754842244975679952869652557254462855193746350400788123074095218946256357261679239666239662244301092122585881018068648348662919541950674252845427889275435507750234548109145267954417960378313003648104684841790423406105985492307211406951887055036692322258566543046734356911362412427298986617861571578591628567598954085413151906383161769059824152301511594503216066037641798697312925802927992304642284408256667198233935674774157210822639868519261466562714860768664606748675713456423305726950769307265140925640526893326696585004866973806614490473898778216984044605401608945943906898160497788985883003900262316713724289765358939628903380815300224902655726564485523598448150186046229715632986175940035189976033020754832012211481737956763819513326406482329873;
B[360]<=2560'd1809412072784440068320620277432767142439581028751092946201239860120350799358355838450649964466134308494852021332426248697956393677319496576852872212080907179070028848197181890574871566017684291930637565870029420110525768813206360618107716430743394801986291369884518556116514748478024039382499329611575671276514025641250993531028470103436754631272996269267257242532346704760442666563370939721035910152483599916894703378689385474372357018275673308806580444358307446926516989759644900450864562764636200516510945476179768825646728870004046771782291211944862436280516500857694649631916802421241762528741561442196633676337165474511238319005548106208026657084377070287937266950502529635454143196568820976108972884068254035883014558135925315173882458712412348880013329300459793;
B[361]<=2560'd1817287597422576927782569829179471050927950145642858448252387142657262748298202798379083471321887702916372467174235142072529279702574482524016102577264393622842295215878818272154867213005765693821464936756333333721931404422406627329148556900877307668493475057799088060237748923570919369304629885110794805433673621297327098276675412992088460270684867556952393344848420429843445827319013107988045473028973298111436181568606394489530970217214004280197653182387680157461435086693778414341365735949651567649521123680630290229356505276649193794397977650989103321872068042318871450221640507764869108045716576179183252948448014529911256266423743529587204690327239992464127437703523128910959246247608539651015266417626939051407691913646244058621043515407517294001575083626209282;
B[362]<=2560'd27106330757801270861088830763127790607653100441577286721026171886590549507980852630005529280886856821934666456772351884877132182822954409001465425467993280335333102627459438755682241815483264622612463923504326947690527257924013894884493928988487746368157401742669781948808299449758566099590242263600536139968773456212530940932983284732288137737385779693554046968721433677542948953071391383384663754817135085109232246755168221096135400008069272075754713651677500459518691459716348735300502600797734922767988073206711063029985809119095835704262140807383795121282683931420204263534396663123663372242829711175086145993836765775986982296607121135539254999090320093555729687965569415245771634400035331288057190988352002554463838180209588249197455390699044426302393122700660737;
B[363]<=2560'd130881051225700908712188262866135890810792362013229825911195701757236774809292184756008242329989573825503565485293848138387915407913699934215115417632152912055611692935283905076060201906590080348269050040927212881534828724409289337630486688956913720793194646508204423116633229608560144450723413496323416381687551412164137666331745825938545106101190690592361912340389814382902528356496951233812491375772502576734372427469561111170008926380768107398473605020928271611583425425871888951749614270907041752325457851814222512202706554714136401317135411320702945844664876969528717729434928499771008869215809317756825903962945230475075247532120336640803546939873150161204110004409274468327039335896852065882228839001526984630121287015127830824416384775999525524233699240972288;
B[364]<=2560'd28792272545320026746382198515766502915433039936344902507211613091652400455657531789513366693535354506032524205323283159574869206262930096040507018647763164769534235179330848260815472968390303567923953429394190281413214498139698141094894308452049429039975195961062506565117505003592788670431696577314409296709684148045320542864800945894854003561338957206561587307937341669772770005548832713598188564846007388542392970414486812241314256038583108171227061714463534008871197062998557379376653033366125015678146726405942511872540084000026375251994397055402731907272629712039950875194617242244775308072325482932216221472440263619181660878796071279216358540910140290633333460559073005454996021419865824354756790982949060646375555939153464748403296918479085036584969577995182336;
B[365]<=2560'd129647645122353628001074517791869509475019654956688160375070478223654553008002954435445261871782571457969240656712631001314712384218292770473461913538802615100485767042987093381711740519590076167156912247740640885402001889866315298716687190733738478557284091817010643851176786706912841723496658218649578234268345710403441078771406382767172042677289574371056157302973419294463598573135915414043168573181887447309459884634793417731521496941032185455751005281464873679485446989661304155574339768326297914889633595313723429091918138471315110113950557486031288838552920676601791352295337121889673855524910987548854114702940327294529800829077695979753375727406321343934349762242767922077248737016963997748039877709438319429651388445517686917263077433406888943276580798468369;
B[366]<=2560'd1718931977810135088461774374876941676209916755673252929050365147937477156379687190403965149653879144234604808171606747998793380201939131400334354686624524918133083019714049647389508838193077412228076878843544823967016105351387563335276573253486360903696406267549948546379425197314998103710094694652002156370538594730770111385383797269756570299735697872883727832585291437748562608377810054578713456896883444581766767754900896275656876453596326527892578257153199222677106780835391791377538782312432250500816173324748667231404356522930084624405993346580985063566233173968840578478989718733154500753451076208375307233117893657740879934351891628424273546207913025729460436116682783133665483270048076492345053820126528155750593767914157528676151495584827252649666586181894177;
B[367]<=2560'd142177733409606286757219600723675117326535341923480581148682329943790189959872763837317603212496110872620495650337443366806603094768356767284241331515781416877623388174869151653705734443434993331449790567741273110435560290770711608066926335875984246119932532444921618339545546021460517113840462520070266781034182811245664174317712967067213444710542645499242679098245787380114761701690473920528639049472887507133207444815528965396986227110643457272285291916518259013660063837396690872663958865373539014284503827181930890568721964580769626190007613353630283988300101512492012324696848747804930712502195967791490301426086975894171607336433929083385567790766513916380339744936933221762012205655713507587526267692259223098763135371906630152820509989708679311901204201603073;
B[368]<=2560'd22798329097307687844484148277083475097279638052977494428445782389816007969530437702872797396954533102930893867313991092572065930080319388632814580451811861707791741537260331568033461954842944303149745345459808761534052728247742306030664214272774353786571865521296027287647528043944141101232012760368743820530226112005698370620797753389850865961346324327773086819061704798433721824646671559303422877408843059464811392712362858283817591304687828817231813994763719270342241957955496217206145291832763486099598975278022685493187505130163752702750351280605946585967022796084682345964590144288935361271491080094518576247147897274706087855504229505734354828762290278329667838813023499793965699051895655076635441810764903962950684635087934033240065;
B[369]<=2560'd5890709092508123048289110339222766559550543700560683939941330397185633572074130577215319223490990070284501679229699358483378652582826826139183040611788762265947144416390960763241273522834419812211339211993960867547564008108313397411649540529014512029109332532896242810563572767140973300192708927487556324625172067605818685062195575431232612374139335768552863172442441555282981438752642002762630682804102522542387361305253466916864836278051339851575935971817529364023285970628559035253860483641331471095316525998905488745996767240929284721257977081531279039067160819750315387013098889401410883383664904242548726570585256573497737969148585350721419791431326357364984531330187429854930452037431334077953389611400960688384508389024231076352;
B[370]<=2560'd349164516133983252332716805237657968280226581174685237491423208106564036308121799225175458650704874688110095419230177221915826305604644221372583374561721239881477704182445124633958742493235892471474695537525280026510850525753713311169790166670097141490876362053313930949160205347584118201938957762857889424016118636440749072679866800182880087388567715518791714680168418303602245680743724302606994478722262833736293136168710571889499584225032070784912205648526341067986662502716298522945530554126053743256110481549555477458989481604967586078811716166651876421857835870677154245514801417754533736505736620696753731769745440100422246278537556024334589759691409872143236314288089884769562484292450501324417535053053704703162708067954458624;
B[371]<=2560'd21363351290246281412849408225998775653228730359772848071930886796248188470873268932259902118683218844093723896269369050804291032338011177030197820782139993534594100621147679541445957241416991326384742383056041081852460129032070893250071684612235804249164974169579496938770154013360549727521236025754961800948958166602723302308685136438084561475634896367246132930658178128374671695382295297870567668310506762499900944578520108588946672800239589505258516632467767151486707775165771039914189883174228542928329568026629123791204797581470915777235198188185806046890735725020961747351479320843063008331186570384030811894360952376311331837023083777059142929267798132941228298519025177954011503534164550939342009653034684390759672960772863005040896;
B[372]<=2560'd5217104701221436823653762554649857160319371686969910157514097568112800247566979068484759022756197576361087429572312945322949539945801113141205348185989587935386924286176884850346377002948900212381850799103812881394500926076241940345752047037820378103361771419885941470916081207849027373094989976386305192261591815108723664020223575490620224083673185159115528551178347914819985710179792674059663279802922867679326074985861825788083516767271074503273149268041557690694265754098890222320058713275922151942158218702832585085786114974152799004394862196671935858594149084613104563556336469886191799041034509648387489760136452945459145195468759833120250970812702164555014752515273645830255990238295140975605498536624983833826529718691298287888;
B[373]<=2560'd5215666867478140185748632202797783309832312819341049771384778003391157008402020471307210826908266569327152989297666907505128321444063319992147303147262132768520806632800160005046890120993815654560903847966703050139478413688510873492389181069880917374799502035543168033294133019905712869733413026637195228250118804488613213520360285761120822879363984935979672638620050448210062888036857267682082311441998639245453523753649691483895499918644173885653616210021305834380948728985367263337302701778630237984979308796351952036623333235021943088960899685208546040716319908097441948759268519234286540792828646569049501985063695625413712753256952997853944013270224965099303543215512479912736673174926692641043357601289352094346114798873240207392;
B[374]<=2560'd81019570741491303426776730564147229239827060298609623781569942111566716534692170237068491836737989071501856680248912464539529105710923095637532933918524513523942683838763092898951291149824714061689506443177555734678999713860357107190806998556252518989169114194456717756508031518961122087469023554923738099495024399898270133233486639957909760870738718482829633238782592773092694702045350882985422548315906093456311567119658756240775745318596940393428107999374292669596374691719812870040553925718064356038005776664492094913647971116167882038812864994624174121060639272974563296989666462318673888114211135861359926548491413985529711794561805882644061294219518095265402412713033560009003293610036629710901341796702801268505063936;
B[375]<=2560'd5062487855714884506332720991185886570275076312780100261989150323358687338959518523069839940508969801177344478671375307291004508291999242737393205900325880039718736168158091425860454475973663651667314441465002525840957127860465112993079239851177346575438994494576969514509038558897968121492377765234455108769579535752810832125686844452898816238901807571082851950383568086340263688565171768193153246509216415439740865626473670747730340029316476375008440120888464953967340775598111656729349224560478061782806694635195726050562347223577052201873607602366417092889392398674593474781006641773353284753829240048973042475367595008276353792021404233570213646083218473503978417263138904654554823820285414643569198783120291716466234372;
B[376]<=2560'd316323439522980975204659822798492738906757922897432819670573669438458307480953532351468872289040481281295670085224185172708045100771491626666415705397327662138823034664791911723806430289248270895622390702355194114137996982920219126127874235016177874008652136518581382011907990510302839021949159053538836622277307693957185272526364154441186904722311862154454435601846205747852097482687498832689495367896867998764918242022816615512866353660342774599495394575984751164328059662272128201174695656133884359415646242250183159056792098922582311239289997193202882121669478480515793549646975752929064198568632868246369864070349784387213116816165067411461601225111755095507897938427363247073627505794286535117458003750448893440045586;
B[377]<=2560'd19765353071606805099374916873917320986471171578899062206951978624465963991582408994249437997104740028139847010909010185790161777443706181079942071352545442457139003190444616289368512614333565636437900300115936592108412537562122569732722647207336088151776296173998653436004248895347903211589275143087164919214654501454489280389320023895258147131620618513516608899995056528680558340579821501096308566984622639384320674101541714785542698083330693282133744265952960026490587330547636475272992808984722255673299417170199880620280539054928848492040531202445657763997679809941766997980722543165673118401773306407571296675843700740093640731995442146692577307249685550569393900678535200439871150471995655645822396150105912875430145;
B[378]<=2560'd105844015879078622111376856045945063345451107374587511611438975902983563222263827957806097164695604750945663384248480056877132044974957035036089732708637540012113608920109938384109077757173961495711503300296938952067037633319735239635166781710657932451937711437653283088681603176188103625691546421871011459646723462728477298399667038595166842490737079160652034882062930989132140240516218250850422269932158895565688851506164088105813336512862033668581118131460035981383146536550116410054427758365487720140553284123703279170720921462180698231693889231657690992514729671460136891998579534988981364988899096169347279999375162832471137886490887003596072088993003249595234867540143335053396423614080111273572599201796096;
B[379]<=2560'd17754795570684222452498024990272947324141124153796922576859474535435122392255915035528967307060306472071892230065778170370578339052677350288760718683880222150213095150136748653939201146138714876337963361103885992749967534299144299127706827716129375691823350764664123861124836561379060997354333807108509787202967218192940498099847897890792432168294301790994886154529442324522796035911715104717433955687729894457650513383161120397049353292858520413379226979994687564258426368981171430110786988621296173210169557818738301991957249016816123437397029844419160882735416472303857451929007169877911014150024207192789016868914438583102394548767373638804665579766167024175345367512123831848368519131429334187035865463712120848;
B[380]<=2560'd73955390214271253734061289446511865964532218298750074907774039146365771723684205471169834114236433902603978870207386296176398789732847964688657295778066290045333910310919408022195088436384052915033127055076891773068703393858020111612119473669806984034840190110474978332949068531665778860578702666298498993530273366699846323603774655737742285295365182370028020994849189038599351177291399077997561376299361201236144775507863128956428258925604384429409216795173086227551129817336661630282774347755717489918619171636174641235392506363961987747874129089393658947062950201142307061576835529556335477372541058542294130453634684814719278720109762680073365788655094591172072798238662779136011479894937889925198442369384464;
B[381]<=2560'd4601989183336459639191606828456500973356309606278919314330968720502572470283661452377726396844708938076955960271268551595577904430293676959563964988433933847538755513684083481253287759841973675919247546886908291088830501694375357918525428342224861152599290329782869004163787235193518124173694343989756444263251268057764892780478528053435486307640692056428822412093502866881417980560349244988777415304768697544545138625701316748086759969737637102824565924015841588250084526488870903925421196910632512285343955476876605821227458717002601683448497872956796178980669813632216948332867213433044953768133779806436190621010147101930449268140333867074500838080816605427203686373718573945138730833038147380263420246888464;
B[382]<=2560'd4684518926687037760893605525714161606683514176923445398933393274826038122851970510340010013581430937508507883468637915810023115369454851433828237597564250463466379976497800482464043042101734342243408502280323693005027784550068872450505211173567831303932690748538772327049607500640746491250124989378453437467379353756993055402908437960581061007961660583561715802500332615157292424699887373684686521621849947452165868329356438223988657562764083837976643089456828895086701529834889727109772837465542711817379027428703658842975450929083158846477636457847132574132388871482071185487083711768948566737844577498663003311618399052872187745893831413229422510366221277170314503463617189925889446413072307936809717776;
B[383]<=2560'd292586242493234440242830380876841030547809808077622697708637582556583072146590597945611532975283400041108177429977095126998728999565389767404042222847052110325365093255369869424844908579044523908771049274598342170516630019463250154385236794077129319016186636579236403077501053562750728290788662801885182983276635457064177472493466595551806442508717904932644805534807664046120468955645571847483656259670831794021479331091458783620489641075587089608943779943941282292140709632401403901894564855282871652504525057855946643323060563995788066031355667211351990280826648947272296765918199717974790816144982887231288052317190110836042611341085323205567525230134016728675091035973409400642384571130250832620032001;
B[384]<=2560'd1143175509063028536869080292967834050283664652080862936223730434803826870833508300456941962073486356555052187026995835528855068994726773698149484890526544628749329107581280909538812232068295153167302017846357354119991036310133824199533202090512275956968828850950607203691050885643042447443847188034940608478033813389499253955876285906590930146434727003340326780953074286134030103669334709208581041756372667414808216068539604710444406878449446844682719480284391543703652802430465471472999849202650173495870807140645353806162852457796878574622933392376022827193139714718836920978704410092713894191001470332164155665379722349290058817757911308945965566488114425806035586853328273647384306622820950000795648;
B[385]<=2560'd8667230658298935556192638798708448511943263604210819187330477369260760532348937766206224186006640140833876014214901481308900053080695753099917391030966742153367711783099800033981237996389563382104195877250917567467034207210220603071638548233607475369219066015322323483736066267888684264074447948358179881887803668103520834816897964702335289736978577726715373446824546110193951620752914967819071565034828154314028049411504019353753937261516921154432671244853815142299706310384719949720861767856676080377467862577390964766669756256673540422558920912664377002406957460959944728823442651750068781313697271801798986542575631754657395621132224878361223859961098963289887523437483804123547859274499352428544;
B[386]<=2560'd4464571615034770476949257265312503491626110656165841124871128744989709921326976613944669759980438889955375512929167879760733078687151994775266462133915639472887241148185029577537893034259182827585771240816447644050868515353562669390635613467865995462146119295362185950530358838441668678495112685565556559156648941854686107707103236752837299723159559270161876400044860791229626939586025620234590337036160500019733957332673133827413788819481551538266818011289347636037922616388498142196661208877848614727745647461210167190817377725896434254557091796381227905217130143712984902908209498854749112779260736988597902832553247914939192585040651814410047785127734151327491579952151045438647277202046481072128;
B[387]<=2560'd66983139811775772252020953777725520700786021588172022601229788635689862813858951699853563349959919415142057076415408292622955784799109081780928379478146321092764617848102720058793161587632852003088093746520319627825557200206277498506807787998121807983592713443224115154898972645118004556285431157113536434890661677515607129989126037764271073945830732631328776339619506540202902732091801433153693539127277499990034781677629190206968109722938280433272285695567271405017138222753553304078940397845264860399961284455204275216983700437136651542706791498356457207743695300132473473421777341282999214786474124439210647075393166648348480176277178512425303912464605229042146682990134939089545069314964346372096;
B[388]<=2560'd4185480290431868619852565438141202338852557845807287640694888630284142372944430861367900714620895216892601280275388693804303117237402597612036234956499401772787300360761047523810053131627143204101642443841226830411195139790239185205081153954077286860673279708974282312849235655842827205596259717669834237103261026074754654324112439000018138823862573442064867338901315298803757294889455311470981337925005525027069677608468120248129447168512414858873003951144366137070183607314300355501049452950825198791171365095779982194587335005835909737754372538173059444500146993679456444252631197926511366662322401526337652810978780661095765061526356742603320601124583222537065530881622591592488995867235650109440;
B[389]<=2560'd400785353137346596115460704607271546206609682149521948596158173019652256594043233178578984993081364812410356808261979344404873644309089338860218009089417078845798060469010737568774471240242478796077073288516564240049832913009059454510407082864233949107379027995444929807408344244016296052724002596580858389098504250882295234296492856111455818640147273935613434336485551354951710547472331644252805602121543030963669849198835884727818984829629794465582855181119467976764364315387709393352131550221101972850947339531273529202617175236322225951738117212092587224838803994305669124858219873057481951111354463824107815445695361439577559930809237932350794780348404871641023901286469442859949427098991287128562789113491209134709248113367285222228642205108535296;
B[390]<=2560'd12828159211716870479923636824733980678479828995339404417731211781191424518744625796297475967213981712660103585548098936051371552519418034317541039390210278932988063982807511421324657392458809495237932069409154566273430880055935654610401189129115146262906545732866109704089452842660069107372396435804980850078290234087639544956494707655354018432603461661257705437992101452233488268251011824274528979226917287670775198083683171634516540230235022517636298776266748182977213490086554381123213524519194485909094234901710782827722609993447387660525078642831304836460014443614916772159841685155937164476143994403227102554068368447431031767987336596688000596423996506131012504749483885448741613418240029823392497636891981450622720471652904717066125274245291311104;
B[391]<=2560'd12804767449820017847632614557476467791618325434020036711819688484759767437986396786403927946668525922011724960598120010456467940010854220231722321324046634909250798932551937394450685325065668372220725430429611570502556962551173181610488891557163838989532133795882500723534204305720609247282753843930623425359705756211212649523724534301359610913423026437270108374098609467214368393484407352615951268920989067290798249023322334025050094817464505441027451481809386637164943989438640485477623301241926181470652929495566273286145479644741523150740443172562704861243497734694416008041044746774907144858967493029403326996555072138093078564028283252727800626869038724927821090780994555670249788407684590886403416012372963458598381459801101304581174613130474422272;
B[392]<=2560'd109016741454249125990573393814407413037758882684390258038289791454389619750857931050241916266475541557084291851859773360179737269859573391039682769652008640485928735845457460282913905602382112759419822298464255920896662242799450448791815488694588066149924710758290645006272419387578632301412597165638430030285322376022678144829510026640867929129195589031882200608426779247359770913026609881609493308872644045502351841177555540344990262795248360273378972471690094884654798458088849442713662181970020511061626885544835371101867371866298960153178219182170601311975579263444995882894947663009149794365009250680908905974041595830303938292468465524416187158561966675513459984132909629807854367727964714789519968173528200296667421861065165389074096834862664122368;
B[393]<=2560'd103026982330438231806869805262035003116429331390727072872701442756889378589839635819046393120234651255542518143985760046272043000704083457876640687446634768835373616546717461225824654295930382183514279190496072639324225533399125760821184765599001910632307307932791279084597949328049030108626430196851708595394434937175131862352277689637560649357991554866181625459045605166739685531631956562860967817498572497230724903445199681020808458544652359692544133164351256040696410712693109624351791380766301055012589946759763502212612609474160518523276815181766985793532466457983879990657590471222154671529404658449727707843901881884058177670763319208137707076887402816522614357893967088188742754567987167843950979970310397749345775055405581632787819619825932566528;
B[394]<=2560'd6437614734768629700104587567754299210943668019526696299063176055410439651889489047873120005539771651531508369871141645599659224934227839442441154423622968476742734891638264551956397627658047737604210919229572085839356288143291127801185592766583496481589766008751628592875940567242952136767816752502440887880463760509065400968334199021959911397751860235178521288721123901775859926308798321002616226637112983963096459618511926631064660881325364430799581352669768061851335865647459533257514294364285781452846980764582498474083820495432322271594243305230647298332278420629820360694105685283002079697777759968558957622687537251676874429331512891168036709429620109053447377102909251285619741370947156924985082976675320050682191918509386231425845360295334117376;
B[395]<=2560'd23489251465925075230210151185774156554233534484953667316032739986389538193089559149557302552408464722169434480372331282021158185487400436747296586100101689568121091109491216164216046348025254807780332018189755195551081845884846116801386263995284721936099365983312015155384769343691200307020775126092794482177169621527480637485807626099030631073982746959445031837302271108348226641193498410557343758420820839223344249747409683751704502216755923856507628507367907613982379465498618958998325499586378881972340891224682712355961634381718494744644859862290339645747506308275728813211117816575198465692821668189904239464455547260107978430638060352503505315717013220729232741179160383188654656677066546700295667172905194964872885410638778314684851072679280640;
B[396]<=2560'd226950964506300163895327879686879413190268394939194869290553088321072998024929926822283356119754441469267322452740612190720632134237430549970636273531643066667380809714903418634582426262221903966236339768006128768171758922939281836363588542549517792350840357740283219280861541991083171292370311493280956898732405025369993455657848264336907953114661394045363237640186161976053607412361749420903390452588749212685760782457184966907620956799835947674635786579054619985963633572536760350500779964307799625416525450663981610445893442859891567776818212201374657821981749238232348416373677038628011213563064869721112610472799298627250498941059014541602792799554206717116716269377788313600;
B[397]<=2560'd1493041787808189526630419137355951764459199019333429443015935368916255410388342450639531113568373300383417760424307677376374729827081739851909033428853748093224650108279417337941948161432077501504965771326173407160039342449617121192820468052574135487067864363277843503088622357034128883374368177612857557980844234000598752432345514273094489479368350909283754862601454597522727331993775323252315931362475536575839804588519600600044717145558339151144226569816912804471866008611511890807850613335270428343241224131229560470723801762966761574194293710090193003453150169560152801892219652128605765838968530342428826641709929241025506317734903438404818946356036832050983216272339237484529383168179371696575864793467707748749661543209462845040297508864;
B[398]<=2560'd96211974006015123228890870695476079128313546304191348489864588473169337045924697513162309585187823279534156372635601753396951302501769325485138405466641157905672344268797937701775770966987445869504049802192998170055407555536084785417222561564452955480300920592086943248369475817265582333404926398594044410758365914447427400129133912422800904695115137929704727251057607084509002452351362697943301872122893627803292689159997178362819530527080665345249748404428174577696793635198997034959773244751857882703260613181373088995220773678312365247952887676742097299595459036717791794002944036401499015784891148694071313562122408866700818360345940919850740686511888933946055346907858436973475313255039690336385246053771623560871014360311206193768500887201792393216;
B[399]<=2560'd413227281832625178624377940173273591162540363609555784489470831439111381486194876550285338970405736458241855100929749914339507991469281123866255135790414725314116992933493461327318008249176977833691632202369417749102511739199807104687284737448853043909222502590174483278526356759190423843193117454915424270670508742210943504760094337534403671474647328496831420286741485889518529691520555448820079449783785577452925064713791428694456406491778611403899960225825872726972709863869381424874106330782757421325405100439649123114653157779599091092224481382601794963512797563988745246272064415222338923837229267677198597476998978928152463648876511997627373554003411789552860535942826967226625013413075074269829980138370014007444723022904936760433744351670537725392973725696;
B[400]<=2560'd3302627480576900045277944190604976378912910739056775796140643191161137136822816672068975550738343136495291137686282827595474639540795864766607713169999696291636489922363218576064347822565616145566051491435515871058351037410995774910444469806162944074559232763676152985227776630273245227772854649504214651873979915117460815403881342331877048793181732138798885048016705052406437076679439365008816251898557559840287987029374029838950530068998124222079851935265836930656105702942152782964918357375762068822692659282783448733940341625662352147852548888965944775853233337662798168216196585408081340426970722619743594916103074868938535649809155062779862640100326092962992750592;
B[401]<=2560'd860029666044216403279718246047628749594245417734645536424901238578750269875845643737530959674976204741520790673464017687272150225838105516786882402733494310290790381432961839546986537180766809565027488932459829415359056563678469777129075410539602058170849268681149146785530256713049157749344253363564471057948548832682451682725031230755873526152988537918431275580433100936397101397302356183076958291050990862378696908281480947416808744678162377717649924765252621190534655630280640270968324188954923863070954196318832791063304127515956646918467680280215008674126180181364484177087047783769134822520378088972349659344028831538001327319196907653692026535365640087142400;
B[402]<=2560'd53960134473244257663923381946554151675476574431959456740643607384227106989175954832193960162971939150945410540726669142390153105750859694199051305599095912646592092097676592012509785312388552521554318299530906491588030809844953404048593239318209218367788463601464010901864547783898051894545343578870425706955576669698604697631420682104774695764026114434601423466176612317325801850466837444930138611840622729758310249207101035759736350752442970176890729481194649459148131789789764650517804752114319839838962965168334372854629759079433892116772945019168314062976628739080306006800857318432789212814133867374184165598146040082033553001095005440082564273220036287528960;
B[403]<=2560'd50590851170528442469924034036686409671508515735438646481693593018546606398027116718407786623964665902646582612514200169992083457384006918308989623250258589866548495416493092354212367200801155237181460392478548075097822129010185388539021426762398811703376882401932052123980874514307997820839381242222920252349365897538211324649181242969452329581180399793965249944496068246553561384233820653711990483597514375719825826081923396083195191626163166099390653586551092260871091710975168485243430305239794153067038678677162172524895438195413918232076798437791794636846495022780621969804488323643735475689450779351489315726460742447874040617903293296193912439872225527463936;
B[404]<=2560'd197668546878914856118256231353719449244528063708079927970389590305161422454533507139299562021142570032584759073704613052319872352105391271242604804990500728927436872250942926301011496169872362454520294017154772907776480576701034960026898014224320304115225273334957843502137936366316106250721558773044632320522137994770635908293100454508719896253620365964132534002283037030671419646263117525525404810331138440475103393401006700484980253199069521363180279111381436249370939599886305467775043955174616846694958195148009235956674611250963535033391270183485490813974418728554816983513351188433693156275770329263070142571123275668990606157104974148819059448174449000448;
B[405]<=2560'd196800527309160435749293526195914967554374265772324650573058265241665542873582889750711481794933230412591804575787324660603951587772009256225413651943183324312637240889057620129441773488250087530437187649232905081968452630759867560126487448369892761858977526654263024456072561594162958839979662570780546645432824221085394413732056885834157173377919008879891696671855468676519175928728864182910452141827762108609402030216211550216526092192857027717267169654061365913685864829708109646466776804142523708013033118264204481148641435796143039225423227900545852067277746100622059042360458732927433541858800647253562841157053471742650310150159698271070486346630376194048;
B[406]<=2560'd48048515274689558292910177415122923251760005619308829380968291066398851843661479026729405079452228030408532883044228869901226415825360226770973426889342776015004953567658143322581585420305119308606117269216833425183650797968412063231937950422867273824558263102563967396579208549735704630862480331486624049512360037801411534371777743201701288767014915897587730782490150733599980758667586177103249378343201636644327290806243459911054234869942507726740010973036533766006124173071901469340564244760652525762082955399762496545050269699556035979597761446927952030754531354537741328704403227420871395771142523341401172058735482746649294715762023147904959243670781952;
B[407]<=2560'd12512204569718033164482190001764712677756554887152306112512514553358956937386524414177560280328254781529791162326606409904199297026974557072571981275791762822321763705606288719233957055782477650455080803853467832177957652342829647679330121529726111158827218983002351973171042146984360782024877658161325460992343634789264550700284471626528748477217051879386510486406094927399255994771133011912152778708645699286656563985407550799232872227699617960151133620476464496137605510234208524605025795977300190159429785906873223178579081416466243766821583561555159154293203335350385729864768881579653765037920938304206240032951255156854273194218076418358856394997760;
B[408]<=2560'd48875842456855914879678186001164436263438736108671269931148860691762681969721710669953301219014043963504843315050004953866237823828074759259856734546030362361914698818197524612547112150505506938461838465496275426926065408156527119915142101710166547076667215999652779968060363692490133271062071523635558529618303160168703682417276130321837833238730366218822945633575719316715433904741634816053369359534767356755951865113281328260749862374765978251798140688786347228449734372057881406858445693901835689400552651808398500901667181522490793956659410901044663820054484010567446262596387798968425806753661658856345462974166061081619805755641767088833362395136;
B[409]<=2560'd2875751652122056253157370280308016895892202502076527998661658131443732181873918529594339791406834083416059888434147712635875902087383653994687333846877422543652497661902955532809112220435016845821110238420572703780220439929009325705216414750983706710900015207586914646711008138334965891059183308175993566084571477944888626491734947594984528486056252420521248990195843054983051751668873006401149247819367260381361739074342301473547578416783611071479819088447722761442335917907689191123237532075424066344131058715626137309131807964352535516665598457120401099918620689829779968020178768597037225612385552264367066485598601743655575957944374205629379641344;
B[410]<=2560'd11233425558539875176110524770427302100015223594209097958299156258110816118504581897163781683377931261674551931418970510301587541314586336041889335224029644060927216598018764079489635377123473886903438743821451716519739996474923537725959735189686214379475795118697322572878996199725205068441524347197615136847697580421384277796918807240012800578262188913040140002550617834596236424014591039426872912944459276017776231349647499955143990804791703567044459496172395029492242778648452998048621136068422765724280162965883158875893575644993312835262462674984466196804197169555913566227989307374825428519254115884878694819826567655337928590851348275319013376;
B[411]<=2560'd46451651406788871696489030128204993265697670177788861770099039518169007939483465303075847695734625214702597750635218758318066420448602843740834155395149161689812715396734844288847015642421363467089424106414142843624564762728961484161021100749917828122373533376802337308886833796096320582889569888655133622525863725685267528789384152245451971997045732895926066181836794104314532661286497290627851297532054796445503513601118797644630102802637458468608326781800480332268882191919805923864575324636066162561468675344208519314983128786753224538006390287347322687932838853163623147480916435565689400437251666775651828469465464742483758968249206374924288;
B[412]<=2560'd2731867143358834214578654664710124436298605868899388973234972499016861885255040292844793548744451914499448434952247173461417107440271175663936192070686193263347192054571985999776086987399586751491425554719472245276705567602514513808443315877980585099230469859886202265352747831273630421356443763856385597620020675993793492072033246130615561707299635762725145442297629737491896522398108839875731411247004878958791064002735742988969106444628316162203136653183901412407229985682315394469378961619391676605167131076903993072047183110045581383955425064229861204526017067436971790405481132003768333746193070354859716112089827893673767557590740000309248;
B[413]<=2560'd669726491216085512492842139083118432240842883003764896381641615480673947073414366031216543004122187495305346465719420789055915452857600546764196291873048643670698122868470076620425955098667199970402680163179439588416421701699267132454105457003014488186729950936152341435510372419047281536482969001132165220808248713740041467669873031676249016969151080555023680937467822389067943234483873052152747398455784595266988268027649134820907013400905611645010944545149470721959576825682588820216429060428244817654574255494323238099616971737968173946308255722186418445507817653163725689762391228791163314482771416093418444857759282748422301816165761024;
B[414]<=2560'd666796965012748854176328823707991594324221729484568795484506752720125048853068664831304057437273246307537316001948723512177259983237511493728796835384432948223268598886531958056167132301544323776876649679439341593440220330231048060060318582175216792092318455426555120983955013961476238525664118180056799754095774103802247658174989731743590073797111713489424651496813383698007129369204718765831462411008397639563984954625493576319524930339756218380100015184925860234189608896462065463136772694948291307227683048610304310479585022741523565955951827451572918743496163984383930308629686080162437279752675633227580583893123111905064684992044466176;
B[415]<=2560'd2605311529851223425871517378978753962864355180491149373094425968276612862714315293200298648922858863048285647453857871005851057571128272085322372422899244953230369387350786824277530348990462438909475726412316402021238527900483752435684638579525058874884719878205116846339398405825950003883446169852089562597052973682004392773651546120822760120318263865109850915883603566497886982880587789640521842436365717925958971159939631356001706002895770035272158196177322624539197808166919943422279872925854528379910365075898965028001302575372949415586990975794991482656363240779098929616111714216727981141709293823939901777980427028160788962476032000;
B[416]<=2560'd40084359876398503263920403629739058798637770770969660754133210542568859628435807219442772863937765334867915590768758106080573246227559272207544580414660195401720530060030823015297688969968975929218833659972581672122269177685490148414631377849354410764056518147758485580277845913680537457778868139742279674780502323883248137220039236081664216592958811167609175656241092684172430602030111111642002080470946052358520038666325958502390274705963388853872716290644146853122461705412170374015697446534167542869423944984408320659177911988324644376369847441730975057919046187747494678498965634849816791555777384495325373682687311308231184220160;
B[417]<=2560'd20699409315623259706481519202690246122145990772328995031465978655603878777784521239660230481207288135501520802250333331212556943647571162886678321460829358628575448171240004921137020148938553436124610847669609820326911581860372255159483268905386687491405464894728371594831047632212175093447874380601380422915245713141897850011730083692285179717482958745407533151139284839544530133427438800688053936001743086034570445631638999737481797531576820074892603038296143814657434244146765735537413808639528489145474208506825710039824839752663798865202276032231540824859320900863321666065306691009236569723656980386548688868288546518744432640;
B[418]<=2560'd9783704367607217155965650421168079295256024994337022434900955900297462975621699987735723326232031290514423903199134080171537176923859627549590959028128368163682282194606434296468541434880447607378259610025486136855697459809501670415493916711225558490545129113358064903154830578810168108594383007102539159624001209046683013359573641316815605628579831529631836737949019446562260499790088191837853694812603246186028488871234513606259453881352444754517494847328643397225978432205408374542936032603518933844847252104489447577711566828813665033686768342938438096105505818407806126525955632871096987541579052922727112610779702899561725952;
B[419]<=2560'd155248102161804532265799015352372003944753073282127399922613121118285941587328041082010141816604569914898148320257745456510002216022014862691825271081621371542558628617307196958778920057651109299051193602811075102290285106277434211038082090812023131971112559580820782156518766412035008997399771307797913459175829451465868618532013756886987103740346090748090558232918725877502297347386319614033860015982285208293739754657531995406478590083646382071044547190645423450408791631729063336375478191536942736419717458257215154646272710692716098833918453256314814412329954580691474467430161117068031646389871653163720883129309858877916839936;
B[420]<=2560'd149285362750795478616626233088618596115151891446191283922148936167838125378017172010543053037639133657370510290049247410295688405786182594570658753455450633015367922031772071494892081492488605663495058698267672434335678533090669864936587102615420225864863784511666470094926900077116369370497085687869582921257903351593621151642753459487690506647902755154243256732488151499321549480885443757762022363121056281430398741646908837589713189152279239763284781393922709851321660899991947859495994800682114760867401398280576111903582154232265805827436190259964453667109880955330239865971336658984305106909021133870527786397426190909440;
B[421]<=2560'd619441373819961736995062977770230570646509008597609665958377757846483370892313422117359782783531445499446504607341623852809284987131822708692549844871204279301752928217869266433474478485749903316687491003300073216188548664722230161398475954202339036436275779526481419595115200323666274917592498137252425904445542869322084819489019452345156564551241007176353020191374973390167814432034797011357431766399424694293269238720726095712815210825914511697212194344405470274850079907956021305270325932386642022487514841637646591487533954550112469144096636663975288697025127878556191583867047165651513666479456797898627063470102675456;
B[422]<=2560'd38706293626204174917915319523918868819543385905532313764439825136524365713873181338689214009830514492196503106619248213222871764701764222469081812914197872132340410115937559456155849313496343203011407125467782593582241812100212191088791451857699063857025319841848752285137259245785162421894920802188158410581975558296975639948653442027958686229274373514043832367910871283726488171634935898774877987196621407479708526605462842047623184179400868694886414752323452333082162673147291350895090492643268312324462684088891878250414085446792348647946106893756449724529954684477288273978118579256729515181744344733014978448794320896;
B[423]<=2560'd578477138529316728128364394270364147576179648657484124336509229182885963021267760282042011573884135503305267517950476023321678659033464936497185279565103083730285599167920435348006752304653869042478045162098543473662126940082306217180262823295218270126979724171484750926310774509310822212307127316004741868338705071277581774054963705365915582935614226234260147587299764526338324336199062507180527797525068286515420652825069656611897939040979269368676043546124358131156699619291798294144023866238226775782137728218927977084014103240666601467939976567986698912293506434022004057607557388925154300926979124159702825623577690112;
B[424]<=2560'd2259124905050219418599973124010168814431155237605020185632529857477020875723843613741518559465888645980231469587426657031364874100287191067086398053926451168012507731304912618292953569349728138720029440030364294863266522506834489350340245599520260525694538265674089137250866839098830988192400458629777466265388552264603572671407885070783380778070022155060929010481602801392153095443567715613558709843634080327266987457798853633597142040840365082264702728593168157243098328921637676160368722339034400393704572230209676165873405775283465194547541421448453626447577746262465264168895103539188078512803900663524819986703974401;
B[425]<=2560'd2298100263170018917009698555547045711334245033480007977141604099244277528882340229441160715826877080073437184162890913590925572232380849076690031762093579334169572403586269242180832392873207426691766964484129758625917259564997567576982543200307664002657492806571223558998240191997629079879378407315616687496456665244562330260837357542926952045638214025551382896696205190349071325414980900875794656058384807751036509893541280686940115834911680671240600813083223011974527813062348738145814862130479731691105747377258014674570853924201810685304412849339161988961700238801209001688599871200971661166422454551846664011776;
B[426]<=2560'd596116262247883622922233253103634506847506108023856972063112939644088604094397050081285724602178568123637344767639645262161224040361271286972474551165624341470620904812785892568540323691744619907411751618953705060352598024769791559231289866869060469039608086590951094007959795585553383272386891910314453406656654042890746539481664669851549991214093319725955258885556256549197794791125445178516278111284782900215014170510788857100341620079619088235739466112710009270179083673189299751152424806540143722640799620850904962813241993167050038608742820749577696300878597125425204580401337822711093271232160903469203456;
B[427]<=2560'd37121856896787398990369676030576741177812261630039655216356809475175009905790052686797351242246386096245223273086919601558792207886313248310731789625828406944128834458555110123868373803648265443128309347708563191292380329555626536812389537859647910939969030276716733565174628875319940035841892577033987117150422716277619306886244945842228931122122110892838111309752983057943048661038570775376614664682938041692888949752968244521128530152565925974273865819800121773238251337819299363954004818001400321535302964965163120000056705270637774978876587622402607732838876271592880304800238138420724069929831980752437248;
B[428]<=2560'd33004044833135452603370796523296335235966974307234532782697001159823087955912928021969362388076372057136101180267476602002403263332600785616246341001239023202686378009199558579748858411377957562894552560322331432732214353113852653169416710006598266727676742186239048144334337314752906555176984517595659457804152933101116273962775580862742724574708789730981187375396147458415076742681407975248267632753379645203562851521855540520444410955459200408376516299490284661960094260705703291619828574351743061558846135933837924559041127506024499268982002412876378666722864938870093327869516087280561768422518984120729600;
B[429]<=2560'd8061424140310454880900279918290852478258089644720012523176392927296596459535969526984469798231610876626501388243750636663092309017978953358817054163388314512031495479526267346586847016185898541303384668721379290258296901406399087409099314824378023337850964647676398941620583743076749395976036015858435535278770253658470799459865988591786783674967492363067944131571195972822248159478569518661039825940264422927401474105625312467370005008177939045511811446010437663087539245427904262110130901105823026128386749575786130328747199344158769708251703385498162449389827407858181810025835006115675952541402660864000;
B[430]<=2560'd34470947149796480785652005224947285203139703410397759192756712110399638624550160117957566465458884852444725257212270130085004333816232366614237973633625371677516166593972984613955656656660470346771424902269017164954269956475694774728099878205616650151060060425475206591950784809018225935347534470658858269531518265909154840277134026697173309411287044400282734066698021780117068407023330388874160773654466746949593373412709495030151264641622143426551191641628698524636099211582659123658040885448200552791286042125663070166782936307607629825338754503724244936241022682849011256367386100048701748478862744649811802193920;
B[431]<=2560'd551543044290772466999209368707138932527517800189565224279318798526624693754272031503137089454128477479452381310523261903948613766944074276712931988887296310453252522204466459764320006592923099602167319412514199237269277173194692037822697403135621201042440539236598018378690789424022147181068763628849287540693278432312743690270194482674915576885807270821466461440325843580047334889278217775526417550442031768028754858899468705237118847040572760867663783654964520586304500383536992946921229230514235635443814917951068702060661236508673492739234084133471770516247714690877808805329935899173041893796624792482698349248512;
B[432]<=2560'd7656438804794914812417123055421329900673201123420705266701169535676447238388288843555000082405213490121234688485318348365235935767032169425937498517331510705110974510303179889477640182740650318338114739571604364879466049676591703530842446624143420200913165492523331144498976175277927455668872568830307780722580819946824801705593267133870144820755541918661212530394862701856990178340843007756582546416545068833666823972398565005796457989822271820902061024525253729687418927203841733656345175734286917906729775369402334595843655499345300272616160911876692198669168411545145961111473802484706787415031808;
B[433]<=2560'd2000610589549994062289857177190539379137075629005540124183040054452758291095599674164031242406241988930185514111832430317539098219622546527700194149018802847157241882927580211789120109775015627369998748635164193879020382796399075399342689107218627833478110011822949621789394861890948072703190152450839517710154289363380640289553157202754345801107212450301900891765580368545178206252800015191802201642771505331086309012469104322498253058852931417255255665174859668320174147410869828882709026420995289819054589806884821735633731016537984762507291066912297345730188329213264555099713833477785008472064;
B[434]<=2560'd124125716511805493136071219538922243603246833024209656653711539214556179707501950463126304854110668275028613101778598411994161898974202255625634976615579248996578555305558068202398637435573549608566365464516716763695983079260019732484739389076307960493473464310954587955014920922980494030943533185717976845674442539697887684281736660169875917051152392625874327439201164817441701305017872255213365820076095146830687906011951596863454941869247227944935919229003571437845071519255139643090769548948774295202815764409964721043436785602897306952641596492115992422427539745082375673374868254988336889856;
B[435]<=2560'd116795794913119249769295683404946229079500625545310828963074870141971129648805333384512800486013709580249923637156529434431655198725644762616348902854169962538078656085032176836762880817135108147697117484643775789076309115710713502794294533134410631518945731488535053383210129219577284546605425667784736987253195346604910184837386124840758173694446680769995244596933355903554580979870226607527850804675660163360353020394165560653512947430867676675369405614242104158662626641105792164117705791514796915265638177837845067784814398885857290503210565996619591381880277131199540809696103913176092901376;
B[436]<=2560'd456233573971928566894565770248657330766841029366032781227932261803367994460965766773100602726503777947816650918247809546481000727148185052077483190870906352733033270697889462198752925925274236879060108340436951694076494243477145648012995554473434662343200673116297747638271054363616094655681385602970210766438397693996623014417177006786064314369573100232873869847475341607926597851387436457791723479989055904174597169468983819950031402531679543376965257925552223923875871988212876414272841978235399215334726144087267596045502365320535016133061606581144547723492608084974515903969331542770057216;
B[437]<=2560'd7398363015128399884669230311707644889471426425959388266254937342252123075631701528437094807517826366948308128339437000883759789899211841930440438231253765851412776712653197652494893932942423491741146767846077049699145655357286444137853446719753484754791729688294189596342045770523227186207559653695475017135451293270574937514875190133034886944462603932836993144189919951922247108431873944142069841066501538034984786035995392525942720476588560113390696905655176936659943445876355160944643285470635710748219347506628981580244109391445038325836011085281751679490126005694191149879488407404544;
B[438]<=2560'd27306917425803680745399532359653921199618136512962453048781426322097956826706650143635562554371720260976191303055737574515523116112738092892063787213120499983812147569979792676166449863130487661240141831113732327570120775922117716322429264883783157860806691729226497567571789310986101540331166881222980879392533145437189548782891523723235277666681460239804205427634903428525004992015708452733247185446785758582841060762649890668606544329233587501199496435308495382282277740012767963625485783719619443643050379599792460652730850898092801924184359378932353550085681613683249248533601058816;
B[439]<=2560'd106252919470556801233693270090743885491106286213760166912249898509334833706519328435180739996815985436180647373630375695243099296585828671047959304419570206735711721509154483144612947441146617690328182169085481085733723888652537645084600864258159145050930868173662976823266661382756196319021479411263947043329548565611621217337527317471560447414132328685861512731503024915310241701642810618072250913171402345890813947156045715443599843143808416458301330964347794108295665542610768691198871686685115259772289717278864935289710467725163385863494128266386209937291316163403206720237862912;
B[440]<=2560'd415050466676178289241786203694770249443489680948470733538432241950974692702771187923898441695630065314322883802024446257977645580352091709997410288851237297270948410129995018986738617316887617094715594365738842089099212057299003503487870301020815803903959868113645360008785878076346132786148982038559661931238392688733090128675373631276565910207778750372936694906339062760014733291410037619845972731952567875432242552597520222412758964832260373294534116014756713287302407515054675288894231185812467183566641576319124999607760380955944403504280444418332832983817360196300874266443776;
B[441]<=2560'd1621660236201928286499986123289647117862803171289590075386996852052515707607208425049582276581473263455705058004193654448948445777490957636525795524848407505815634063486603689256823900211496589694621202639732778413905899758637521396393287123533319522386560853123547546244455114706854877998326429840478867923840826000710483497586824156636563537204870064687263188229516219230879752931192220645528344570737351546506680204126875943543757950811678272346160039371974933862943437526651603103672217925588483878629925463247613624668491373980794128825925879084932302855072087600336939778048;
B[442]<=2560'd6333161107380288473492103209174136892863661301320424407503063628314557176037370729992778533454328352456802155704634097002232418063569548708112971742529888058696341092063188840900522330230432205825829734681240392399553765647316224291629374429255003048847801372995527879938458532468848548495583362887223285927606778145040219281919891617130342039153308023743407079329522914747303745039701010816751836885950104407296726428949352141326116482792259273978875850873060327594703539174756957186449052323966996684553604212176725356308095569037482084510700797767677774769809897722262585344;
B[443]<=2560'd6331422155892634360270098696092531291624822516333409922957531893942554854193272668733530297885565687904361978176569105217588662933137079232545654121052541368827162643035588880502539965382611233014811592443423135420728627425174721869839048561484412570454604186050075123871843584739993999121933862028093089705188784765644848171540399310167248771169368621714409828985332864919404110150891144950748228329757611548177024800340894845123041814356015958552750084880008540483438167319172099628375216288626464936817438377495342488894161295425311756895275127534660112817481630634458742784;
B[444]<=2560'd24732092643836218448717087237330820698612448024611148978727351061888391795310737713264261674541452721441795223620180090737628818038488129154467242974767881787398462458611609813492453290037348506985266329783479457740754391247143499183942310402496800748286979059026634263474524932005726188427793409229298619478585909330718311842512055476133522779355704264020655995329339655631306853539173044960658806144242209069734853354631283165392074810013558042108643229827617041933517348040560504485958113448884053033990126011510079522730974533731821589980856746361688241680530245196709888;
B[445]<=2560'd1468387807174999947067579053373722106580037753082625660613209150308299146532598150241317050632728977857331014375712641692422247265108141919184077429336956643159925585461025981624458293407677494802717067916004496654163993857384594419987024567674639242476974659020215779808769791463920206522650072037032223993148019705135546751693878562606601142520143576818819416427392293875615456069473329671393508732189000641488273329337307307809197968209726899860785444109800787127468578230095773641635793917242799858081112356826468917067859165146983345418711560751193587704047599616;
B[446]<=2560'd23580580668163234444085240092114506121523886107087525370647800699088975667353240394644562877576083080072362574232783859278518281624477307947869067184948646658974350967398005717979017860952558257061436948078768756626575061815844613099666769907949351305011558053801938647150132698676940533306302106457815266993674642653756090209241233200680856351522362717877697611768732350760236118907846555518272802315893081852123250476735458002864624853697212879099224638019649380189598574187299325014496840470124053964278025095937177893777989248470730128753530665291514989976458625024;
B[447]<=2560'd3404095678729953194445350767193377554772305394818209054158020109413036728030560691502229786231297301535950377300173248329349969560205906740852972831895066909191364981765034092045342735629559938563706579704572727059856586284143796793105409073499553203249706946188296189931228400920953535027642761494899206531188696232621501263587240926961883113713698654099745525294552165978990334427428559611454945374894648443070790799357379404972643861498985295176412028662719109948146151584451227077446466929688576;
B[448]<=2560'd3807419956475406532101045332951036701115542510027811749401465741396419878278743424312594864555870532270478706741486738797532105562499869537920430169867333492273987444511347229364259073288848194772354962190648448961297061838118391471401398145754456971236783406892430868326692318314206608480638958344965696193849656437400299376246544503021164816668012901929452341717901456609229070962659151972712412892656104914010709133793102856475779060656245831294628328610292409191986070635878893370335037751959975100416;
B[449]<=2560'd59100688741659719942749924877821584257333112056241163058458134513405102104647708504128654285546301593760068299084883448909334507017779280843015304270484241080770738343242865448300470126931394107251255798027734587858343388430904599613310586901756627471015808601338149185728800401562984381063362948057101938739346846105795561961637740139653546698862894573795507836801898330166087274512904428559819835463152554352476990038174648152383642149452724393070765640199721884110470775262607929327105085212470822884710422784507905;
B[450]<=2560'd14624524117821039677256367059490237319380646047238685368429784868001898463734153916609127700720873974620968313781895460242019273484123220666544525182638352547645911917807790950852696540890431042227791811266011771308783321459996528727155847700582626139225911078894065080433737255735623958035961742512892666799910941397544174153307877964153500040976408304711230254158054236260598499459600342356098751373102165319391647794245622621261816659529995471925595656247388047584440297082998449253760992574302161542840320;
B[451]<=2560'd4061368421194579437567560047135901422245973094860309456605505289793787599938680848989772930756819129881745804402733733548275651011092921060682120970775010799278814185060937471618982609375822600155012280900289660989469042435887832921251214561447476002831616718480205464066979771585534773627829693594953869332332827272984100695140031900153444560066979434917108920795738828817888851570947046212734579305746803061266890529934181023982305648738335580930421020335642206763752581658849682824222417325308539293397654257610820358649151488;
B[452]<=2560'd1057906232813924660752511189917733576172294503334185907086002986498703309903388070524052322245836536623245074796683122289277605204639909378357101952875300638603507724113775151827066001204387811545698257702941082617838962772838454952614930157451542272055961726872097402512361236226778175421054036684034674513503864115367581159673401926642923108665496603471149218399641087982770952492577723861547209967656781808912951719044431779308896067144016260677295884887400710458173758702278952940963194603373321576475704479928343804772352;
B[453]<=2560'd1104979952541304111038417197626446667439481177524809333230226897933955412163091797319302720083606345723098653183809860562426440960484927352720908489154591371191389959546072146176141926755944013262811476603769634866967391012110919115636972356430096383498059038082002427626857348450747582111620067718746727855597514704902895491029647163740771382691435021510876628931276819715703769900200315672082619199579802705433212058168335807393699611718276159355098390398025226230957287668157811653907952261476296242993300155149143836636695494656;
B[454]<=2560'd1044345983218480729687467758841778890240210388523603063683842197285741710099658298764122361896617494697725043230039835209422400830703812647788374169336294672128499297077143998941615557497807527359197558140373450546931144322185828967856910428084644653255381590771214964434763912722157508253952627616524972764452131805368750334525767570889418089644796759482878001134197114025044575586545760720166000406834482038799895764925777101426166950456521249747723174051452037170828058655500913354745556929815389426169105316207628471432533508096;
B[455]<=2560'd4889444834773350727970927856762950601011131213187756318634190728266983301734138803771683460002539823248871384633975998702720666702478471474105338089394870892685408660212694579398091726744248091971355984703640533654868208760184991223689170397270216258015645848229634855786810979591243181562821525189083457261879748078871167006603285425005873445531916708584391296217863403636656696793555488242356201413074744000081738902709437617592918161230225244698599847142732199478330098633082929258887504534645090450537036540037327138009907200;
B[456]<=2560'd35532923950314040371555233996418615656447617690238539146959371986022792206109678041799221488951283430456014754938233744266582558224172189085871013865500498498907118697460000900058252692829444547957332045328413014521689407863938805410341629192057365368890109778500554930922573071833010205103659946557526948495399908050295616591672457345343194686373971226445887948692820862572106913373574766175859371754302257453488041975891127972226578275030048629901981605157469425742802479364165313833308347102684519865090746045046167182925002621073876938294923133313976514303154556757746635214254300607971499956245637792070314612036186258014208;
B[457]<=2560'd1109565847988063696224845352873564437740752949623496227822692462621524836530211924974680966850216832901387650706957187701203820925171788058092251780530796624470752817589989881936317610481588862676394708303399422503522318497657108201084876503178834828805578537026517985474938764700679041583905587826546584682597745752887150225596825513900477440098656218721715220892267818164293746879907536540899048765619276698530745588548062733509608845613737963337180876586042234868184295600062093015125216275422220120441803315535975666566108807168;
B[458]<=2560'd38255062034877977026177430990952923613463943870659685930130103617759745372704032637476828005426439748524180888007875670453460111263669772904047693340057990799911178895050649262958455479373057822731656893750054002814924384903448855704194997568350050711274871141433994239689221031535170578713176258982274891573520673222003857689470752895932409276548616629710070452621658004581266482973299470515147869125965756226250871673055537281763692155014625099670024432417610399870120614243227040710826780834865676706434971272315409133601221363108458624092249421819204699789868906261771233920753425771776116408478934540379578112755630080;
B[459]<=2560'd614463660781673250365106002283749036033562724732187758088802563991857915060418525501427928489607968127247041478034983017801875056637059141227020814410111718555376336039338625383955145785546643676061364710015250263963015517660536203750500590968760496993925096546935910023338942818120138815266426659363604710196922427545518423796913807718336761512931906249292989460242350588492623574668622276433296197008201090576260983664813654083012670134329079053956198230934015717357071358059129231494258554238557059446286151542652460397520855969501069045367543729151931635389916643997041541591308446807135517679546695197406209605407604736;
B[460]<=2560'd148053840968278043675487748069868570782390191710724277435355876923779975663270771449753700894474177607122735488698616935222721316013452292064184104000889859413355673947174235269136521262670216087466243416738024214100067543868455358191767404861728447576018011618731925805533967487139417475244082497617857419578754590678608912003601167815325173892806523453324120503217984429315693356854396039233162184912500630622436647338574973662195963182960787541565858118838077309008938215564333838893421793410219139290279326789326388147153851208948337638126456898563803892796618413863559635487743778122378669738080554813352574271970319794176;
B[461]<=2560'd2386751587479084783067464634008171421557021195198603656518735358348016781620299735265953848423155179115930140943553938029843353983896682011585063655478525689476423859381859986783100282986498650302541491599250216431075579978194643848945277448271732191865926683992113565907319798475682690855187501758080354557531470186657701798246266882321123730267626851738414780411399363808846173636030456830317770962036011972607822281554934321019574132491628750391091499564170714304553281534768647905457340047945071920238054796970194680691945193289046668323005409793140152529508522619216522976997527427907807475821246135507426446450822918176768;
B[462]<=2560'd841936398104496881132935423046398685275229286403152049668558544893480021002839700525751375760954307627690336016570167637935520443357097454760057775738365821362531695111620736969727580222167890992337650367841149785000257700401558718768638321087751579745211836606976156540240304042183724047315666420426346042272482305208206916051046352846961470636560775488233712129185511565280127884789555138922970705712429087764966292033633692527030562308693310396781891278151004613163733591436242275648175722480511222991108041518415440496295339373653992343383742321268687886510943598888867079028560808341299318507156033944441832125589585438099093136605883298747470262141072517954020573184;
B[463]<=2560'd13523808992651798873823001222073777849446997989673553648465361596418168648438443223972667443404837465696653277170851089602721564966060818140334219443420943866342761897007010230017343731758589194245170669653458336153060977852566989109733791960081203283592390946380085140344545505626855605692995921425108969459352165435380870953884680522073568298418129457742833441912762925655686701129431145235603557781689823695499904846336912640629522599499491004354023907804515667285270618582265438657093948946128932963820817085113147419809796352349701426757322730878378128811411127930255790289351487050427443545430220163663973305755490671584000884544455650344097042959442179211581049602048;
B[464]<=2560'd7024863791154628036614424982945651049763186181362448336321004134464893485265312901412722365035235431798031615811684711166928422262068303475427845913996289055747463839839763374802428806662759225603692159881466484408296272069972636160539748598865460264094868967658891938600935134267741205214574679953056650144811996488874117696231001540311874042979938110987074772540215927135837373848636625350978078665190630145922194517968147960592464941663814181012622029607607370107599820841022308200461047519514544136948322813783635697056827265200677977162729957791734304476898468139427219643945451417397952163451356003752352450848583109574216658618373933870246246191145956825905424337923952191140450542809089512895489579420570671019691183886312340939853709411679973316086918545408;
B[465]<=2560'd7052405550912491353564068444622593558974638321640420593141894269817937695146099565384251062843788570519763978071177184905966148535842517951974185830066757542975873687009736140551750691888288385583111588533466816822931317584104815885209162129237317033070034751130692397316548665206175000804461703802094724860344821364539039246928477631941250605837974623839005781065413476266905477108984799839673781931296060037581322501288905583719753037175567242582537013619633016479520536606991800636864422905687146055964197044863912185206983048366815767656635800773378615840248999703184050338115373718342068121149429645664077468361487232626134379149014285543553951305265387761941790164292354145382614399233848738523198672185141690082929723285971847829918499698587695004801314062336;
B[466]<=2560'd27187490095373768866656252185663885462697105390340268912996236962323234001038299727695846890211354490043333180694043575367443350060536738963733150744583665147575346138489242405936064100247751883775497821036550072476488978227200617378412976145921740567841545903233687191819378417830746024889115842654259628683404488146723535026046661541778508843951584050270970769722529334302864611572300219076535673967088548661933749223216728484001597044670249193913798202681438924434285075728994342264310453319595029459246108350861030156154466013250026291360684501769974995208455532414896304017738223878992358633230309792884328332982752020502965821121529870068170778443020655379695072577828594099938641324610974990732570382405813065757848328412310068091160503710782045791154756384718848;
B[467]<=2560'd7050690496378207249635476162499193882185989810623667608830920116958959703795668509513248516316424635066484533185987051535200839069190870695619994922358613682071546803686754358269511898208498322092726301762234018127227814790622167572236963536291519752787108517213395430180398728798839785780924251377604896610048507888087253277622448104864336095342007120228425969390251828351959926736603256965729503137042421963837992924533443984598596843290722921035068197457230561749161169712173852702766612679022845777729339559966318098721788569010553642688732563745731754843633648484657610195339273370959891725688644889555922220208350537424017443328545612239830573003141247809620115977329005362334196320940946930848634704488185820880145234179012251487252793790043146705070660255744;
B[468]<=2560'd440668157658840634450211847747990773821109300669372193680922265138140020140244865432216943577845542486945899494021708852587240088859272437405628164067283448869288708408975913116312350051188857027343552831224010791632560137814969296412753058123788799251130083105610884822683681508146383431220533319570235276883325073051182168414387460650984788432305854497631747737546624871270224784717923030146598054235538922810741882453841177310366379856064386193892312601676707746536882459923771671605361287219765188714629281609885345934816175696657264519226785870421647162851102966246380876720087582230774720829849367188012580782650315909186964920451817998662221963810822068453587923594934887283379135961066849301343684780241009441685207807532107011140629850072819374080386924544;
B[469]<=2560'd27548065201605893895275016815092551355112543856190167465953844165510375375878170321613918423549900033987297920672303720220921201794285902519344623633300539384264430972961464159189071837886648950623241760550376929974906153466365731872478631595619555247640107945779452176064077480072978801672040924236514097665814488927523671246415426883826648747041756072458507300282048875999321152751198841303018840778344083793124103082102430181942785511315947168269147356951854139705824551574651356442385739277332175743122565756988338508736286912537029638101606964379140904361848599259383873369903186609985138885718528812191942118862424846303701662526702108842257649038179630965040530188512622852650080995390463443886768284023973115139114217520280855668471192154284602168149278720;
B[470]<=2560'd440674461371165429876417531827802870094204256056465902008988901576839948051625062916171308598357151131834561631425752138458998300447891998828306386711709837082390808332393757126442794358774087479746001769500924178699249103353353120853294897536328911656387259522350083931975546234857047499897657292501126177267673486426761462761118766778859965651448407646129236259626531468167173929812958875979920207888100280316599367946812027471599455255873684628394540957662853128528057958037421432423167893804693230831384983584793323197930196665415316493036154199573320854711464607809332851714536916073793597586431079384128328553855198768769555525100973689551487271427348641048352978308000367299430063366895475610692349447719928991403898396083669602268625512876274539792166813696;
B[471]<=2560'd119916828657152135302748932403537743094615025381481930190780897109716353445238682461886686670964511771452348588116668130454187457281287622651502244632898176473099153751968170724180608088886884341520357788056368446898079320770721328504222252077603438257535936157762251684667658452490218082221911227420628428715524209848894844167355920738590300754923803823111431753681817824835736700785413060969301200615569179166807728534655811439475274927087902754980597339007188730095152644878582290014810859646067086502435116150520158030991829363811780294200957115447590438126306385595795149947654003934311776472515608548111546981701851013271208501720235329152879238114429199070803164593615368156444733704793088671791773567512405566323918070149338485399777860960392124788269620658176;
B[472]<=2560'd88578709692552567531994696877192844054783052223455324498549479127214563286009424607940604117219077294303806868877179257242025774254921612342775361998477803604934668523495876239864228164155676319053239799642017254835178982868005502295653941910871130039433974748574143175824383915630838866810152863242525864919192769423851206424498347912575363747125217396478749593138049753389930535618921817668354888967455150844649477852076423553096715743663061601833591804378142618926822988504600105318895208252162615634407099108777587584893917860955301732507642843160740886588738056556931576950838723090587786873599402404789212572061352476379298334711582318176099806303965350486988750431716613533265675130772676106587226677422412888562401276461119536892281723410825078158580544713064448;
B[473]<=2560'd202206737131696770253142860902643793962996942683750308583543319105254822981769702796268132946164238561087553522805316340958825283631763597435511151233359262663685450790138848506647769041587359452525927237058779648360844933594178165703809320448761231703259068714294169004606818550737965761180982510858596647656383340138625035959223261867382604507874807755823789074471540987207680373979829012224512225902640058981537410775544103218081344899009381729670883907217959568407586961627305194911173978175341389038936248771403946953296031334995557653575205291581689267553931804966992606436581531179863671422038051960805935390963919451087546529427121223425468223797094577729502777413704344342888371660252641103935303854732201159988102589579843132690122636785388146795456412904325392;
B[474]<=2560'd232786022690669003021107984954579653930663622802977608384395393438615289176570733506188295287719308549319251778892840119731671444374508670960542346657462880154579154457978640469876003713956369742293505997749852937926872321464855434205473585624782701821443786720067963786963623725361082710698251781816161520823788636310170903613105078541808292253307704238760656168469119930201099778509313670064641045612945005215060517960461596327180215686957622636885036506338147718557854497833261611656256323499173709890918266717383405302772326832851496893981221937806119056421767421904432925912201737688999913463864295387896356704649211732527526052637041642464284398375951306662069751614103011401185277633900286437510746552526793725161447974729420492084813074149827206056071082215997456;
B[475]<=2560'd259973512799914427868665841100064132955334130775296493738914518023112812036433164574316971296901491207608048917976790437254888955224378051613530011747443135025592646598399904913140515501124647107622816329927764490598997601339419138457525635134713323993363947409904089635072616431711563410859117428022952210656178721170609844322238983663937379648165146621512299578964638337208456219270919822931396243756965092485982197320070622012260474364818436675356488635069000513423599651827550420084822821000073333768689736573722525490037267827321993493817423855761996828153618133516622186786394880451514941082818267674850190318922075825774559841232567060427556690436773386507158204384627229466190124278186511150958058092906941919307866616777268449715175453622981018559298392273522961;
B[476]<=2560'd231093884533947889734268991835940435075553562158201233934515684860112863254567669911303305066538767612318902486728687531771043269248765420273525232768286931932256555141189464070353690048276431956135437039422430724429259435047019316965980459275041208251021934067896300133130461931195309862095772950794469124469881628483727728540756152256734804488647494684827817445742134262936475137620869380966679818746391231754785125710406370127824087146114432573115220563348372565174092441489288025965350959192639410044585399751410447713481898966877995397127758115025532700116862477948999992457689009020599501270155252650498394932127156525785810363206527090098692237262091709762772991062942144034432852187572740159087913351560844197253056360959925613500715282156064110877959867545489681;
B[477]<=2560'd117359633464110863205513229926789107402920834876925534334911703923947725433265753532011627462031738292062282952227387643707255948475088731701125800781502889405058420219577532524591169327931991610378478837514425337148132676125251509619950406678706204720306305836312521727696176237638076305550712746421130739934899698614819567650971835505443631771922303883608500274612609037019788818727604382247930814278793614714258211292457296442060918175744094306540580471359706602881382092888064364140962206758094249003625685175962254912162122198950376442843465999898639658817004315799236457465852490000317608367922578789547766291714728237441766842547511403126732629334578760409430019844187637553132031016827052312262662786808943086719385323961226059260889337459106966323680400229086002;
B[478]<=2560'd59586273815900966936186018454575680998241954810537439500449433791868865150274677070150577161144317953513698192472312697946478636708197582740474791298848463707831170586386354806562753527784078763600188858257100775747868904232324626970174569807056419698048801761929937686367231667966839572106398627472788375977314910633239671855791561364656868058760032770353089456553444302823681608353570928808686833372522508777465406276360708615842022440851038725746780203934082230027624674589390777734913279295347956438083142744845515046209292482170181438930905271312335102561275123860641438435970319754031712514917732260690935700291949532862080776916649022927516175064778773093860509456987840759693155067697878577870829524946827188641799009421640654127107420316557293648987760186512981;
B[479]<=2560'd117457926466941821840695740754478637940381819086616500533253102861783707937945987063075407701911892458358792299337024361180259347567819763486701878339667537998096568433418217801374333376001499265036608773365763503872723311172504419501892160311377024027441335248436036103762354449690479052312958637047508217043285479524839896375587619630840327597390946738625575855649315588894540230281944863667297703176429842430230161071736515795047800701276971144671019435601074832706089769670016715834216060193195919051756729653997824106423604272832595842665602904872289009715659758599444404926798643117141059632815942861510042057939511581276281766225174759649183582900716026477436334352452640256054858584053549888708413941194635412601473430260106468279963408643069657303771459850744338;
end

//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)   pixel_data <= 12'd0;
    else begin
        pixel_data <= {R[pixel_y][pixel_x*4:pixel_x*4+3],G[pixel_y][pixel_x*4:pixel_x*4+3],B[pixel_y][pixel_x*4:pixel_x*4+3]};
    end
    
end  
endmodule


// The whole VGA 
module VGA_out_color(
    input sys_clk,
    input sys_rst_n,
    input [1:0] choise,
    //VGA
    output vga_hs,
    output vga_vs,
    output [11:0] vga_rgb);

//Wire define
wire vga_clk_w;
wire [11:0] pixel_data;
wire [9:0] pixel_x;
wire [9:0] pixel_y;

//****************************Main Code**************************
// 这样的话每个VGA输出都有个时钟分频
//优化的时候可以将时钟分频拿出来
clockDiv clkdiv1(
     .sys_clk(sys_clk),         
     .sys_rst_n(sys_rst_n),
     .clk_25M(vga_clk_w));

vga_driver_color VGAdriver1(
    .vga_clk(vga_clk_w),   
    .sys_rst_n(sys_rst_n),
  
    .vga_hs(vga_hs),      // 行同步
    .vga_vs(vga_vs),      // 场同步
    .vga_rgb(vga_rgb),      //4+4+4
    
    .pixel_data(pixel_data),    //像素点RGB data
    .pixel_x(pixel_x),       //像素点横坐标
    .pixel_y(pixel_y)        //像素点纵坐标
);
 
vga_display_color vgadisplay1(
    .vga_clk(vga_clk_w),
    .sys_rst_n(sys_rst_n),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .choise(choise),
    .pixel_data(pixel_data));

=======
`timescale 1ns / 1ps


// VGA Driver
module vga_driver_color(
    input vga_clk,      // VGA驱动时钟
    input sys_rst_n,    // 复位信号
    //VGA
    output vga_hs,      // 行同步
    output vga_vs,      // 场同步
    output [11:0] vga_rgb, //4+4+4
    
    input [11:0] pixel_data,    //像素点RGB data
    output [9:0] pixel_x,       //像素点横坐标
    output [9:0] pixel_y        //像素点纵坐标
);

// some parameters for sure in the reference Table 
parameter H_SYNC = 10'd96;
parameter H_BACK = 10'd48;
parameter H_DISP = 10'd640;
parameter H_FRONT = 10'd16;
parameter H_TOTAL = 10'd800;

parameter V_SYNC = 10'd2;
parameter V_BACK = 10'd33;
parameter V_DISP = 10'd480;
parameter V_FRONT = 10'd10;
parameter V_TOTAL = 10'd525;

// counters for H and V
reg [9:0] cnt_h;
reg [9:0] cnt_v;

wire vga_en; // 使能控制rgb数据输出
wire data_req;

//*******************************Main Code************************************
//VGA 行场同步信号
assign vga_hs = (cnt_h <= H_SYNC - 1'b1) ? 1'b0 : 1'b1;
assign vga_vs = (cnt_v <= V_SYNC - 1'b1) ? 1'b0 : 1'b1;

// 使能使RGB输出 // 范围内输出
assign vga_en = (((cnt_h >= H_SYNC + H_BACK) && (cnt_h < H_SYNC + H_BACK +H_DISP))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;

//在范围内RGB赋值
assign vga_rgb = vga_en ? pixel_data : 12'b0;

// 请求像素点颜色数据输入
assign data_req = (((cnt_h >= H_SYNC + H_BACK -1'b1) && (cnt_h < H_SYNC + H_BACK +H_DISP -1'b1))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;
// 像素点坐标
assign pixel_x = data_req ? (cnt_h - (H_SYNC + H_BACK -1'b1)) : 10'd0;
assign pixel_y = data_req ? (cnt_v - (V_SYNC + V_BACK -1'b1)) : 10'd0;

// H counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_h <= 10'd0;
    else begin
        if(cnt_h < H_TOTAL - 1'b1)  cnt_h <= cnt_h + 1'b1;
        else cnt_h <= 10'd0;
    end
end
// V counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_v <= 10'd0;
    else if(cnt_h == H_TOTAL - 1'b1) begin
        if(cnt_v < V_TOTAL - 1'b1)  cnt_v <= cnt_v + 1'b1;
        else cnt_v <= 10'd0;
    end
end
endmodule 


module vga_display_color(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input [1:0] choise,
    output reg [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;

// some frequently-used colors define
localparam WHITE = 12'b1111_1111_1111;
localparam BLACK = 12'b0000_0000_0000;
localparam RED = 12'b1111_0000_0000;
localparam GREEN = 12'b0000_1111_0000;
localparam BLUE = 12'b0000_00000_1111;

reg [0:2559] R [479:0];
reg [0:2559] G [479:0];
reg [0:2559] B [479:0];

always @(posedge vga_clk) begin
R[0]<=2560'd57773361369990237240164763066017403883580237145113726174237184464633430536881379704668765882949592769943095726393019195080462436110363548445401715084698459841028804720554902658797917499672002546284335684299428851956696145193687051064533984917986117588265178082279972299963448370517262940711401196393493785948946391031390212656556196078529908776626520098456552924873713331570781743344007272375654812391946626983038622980391777307398228455721912090214557028816033489281662535282256277936157945663097328812396618759730569418434161833682606279052447384793699421351145666432457118783159884422467460781508768303013775325807625349073694943406561017475943324878474682604333835662100419831213315705742077550981914250740031789378960689210356679965010245019266395543649263974228514;
R[1]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216088429764176574501715678693841121967005747024074171202276246624088493021737110524699468503125261701810236879024817040830069340769061379279873840948439722211629580351034406346611401581758567459769282064012343433941323293442646943430773547195416564914482697354782658914282337598440339692087669623842130433660382000798614631721697639771750262520310434245839077123876327820676950438156811783014032158960479487655080012756721387039865005655949661088204289626259320903591019200966799666230500896552365794627077346660489231099739086310161685650431601195469583812466059903344102030012484897204042957444661445739434209243740219843250908962234992368789134055372950217250;
R[2]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713664168093303524910524452971021490350172490437450354317788664934684426241290213337230996453027222904174072909745368027041822195712787735534177734524762104051879940128748202768596837656022460235736229405418116829153124227614529894034675531120700559133009090840853794077967124796479662784386085477138356734953639084599901164502212000999199846592724083100949017437838690984147965532103752764267723902025581347968441414756199250378304553269598740910085392756620186487139974671238414387642749608856059769244395355471496258406201497544120169880374351761307784896490999979584268371927157158174870201941787391115795171051840526176990938310207469184241502619672376242281259554;
R[3]<=2560'd30692098227807313533837530378821745813072426625859374633279472014017725084571737912433901425251006783517886740174884802759395351739350849896827899861749878862779748577022881944868651600722661676566575011048452230221223228844741781002165358656764311248043797008065665858311197977789489852738981996677925463363453940761485231938941581650736137272199444992429990747765471568206604260816335895789745552689506320230048975817128513437214414776577473685708320464001876218499491098968630421386375051054742019730145178180257970951194389867072233349762934500677328186609196933530102595878836502922044829061080386537378917832637661044580598062213217988030162663890992245289257188925808648386371026818194078477172116958315263694159359436283603367320975536096054597340533817602089506;
R[4]<=2560'd30692098227807313533837530378821745813152011305451294277942221797086083963356503086880359007406440266948310936451834750739615634148023284954389064762283809336935828302565986918637568481961293298878944554309717815161532424378801406979614257263258798831516965528472238966316825136661402276463515125837102873914220503442617255076920930442584298492242984955486846082067547086784124487679610934875542805536768030560710315650163080083461474184200593123880912778369792713999373398053029104786826781095602620284752208541092792176921609261161114292920884755459921480922980927002138087533411607297392310147211593559239205847617391138605626605928180818276444493830926783147991457738316715814963357266900926984976635612346160073896314496476167480011607541185787931013158618452337186;
R[5]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478987703174675699725083475815399968900807590842845489558260995171488520159947707181790279877926310771254769280586542744827918100057703622466556989012755670758340944933631687589444024697178887451180323965527020605167072868767723894035475864108315467691297843489672465763936698519735085163285856945144331545828622621777740111855337044153921297390757054460163872846432058011989492667139067022033017353005124665027437016174598347659906551917911560368158440784344930682542765505644831421369201536609652847972933745355670831166946410418786978254126395062603036834161847977811626873970108985727738539551587450510526002491181247768256560180969668604819134280760369087320496029771419378792931874;
R[6]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661228337411958397705942183078003852262345519021338547303876438626762374586278906266824968170714550572011111305369817014004157502333022222607221998803717511837111783557950693373286481509525038020478427842498146332318119171025486380203349924186038585457182968459033775049674037702434105617821638910627835641685827602148171788449442362428890673440353893563812044794362130233262138235007927854794113972556379034947381089143541543805462535957630439727825340610556401528040532275390090830587842418637833881285476050649429224126877366278382281162988194683867341786438576625680766379289859282365444275588431927226466832105114736677033880745576727320351568919027414277956130;
R[7]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661227616718640421333015426271627208581362591230083995801291952254796521672200830716457480355152468402572808827371221927929572757393964327899000909086975306328409277648164047024307714445545726697245131823913066439449876077387349488603925008172744089187704093106423790873414702623815711455863643304688464036543229931113422718259615122764882864979858234361285355909374605204681309062399152433320483141046017484670371885637837570269843827337473987875512296330493698309207467782443639509492324690524985884373850041758092182843604416140145733961997958277958773189341270714818600787555705801468788889920955964564172251657635190035917785655805118394890747196693227436646946;
R[8]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516479804513887292444896417371762181161000709713768085153373143030196806614527170808845080655822930521734703617094073296796865624609980420913154456523598113580409695633353262931999136865180691564256507186550180304715173916042630109830757232897751070177884065717851106558278445780183648676823415547724570008698754571357211806859109698424524692351651367547387800704839390803636878102474107209364163087812580379650339215798907736690761696259600484244999417137391231866947225687083452469729851008573714391118704579974940816577136067046700934830983617597654623159020452385950089813909939350777243145338270055953855353172229571096182291491554342109087294073640886854261114098134671229727805678114;
R[9]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516479804513887292444896417371762181163685458001673307052009043586791471421229999582145415440846807209742169854505089433349763973193160174993690785591753820243093829099554795717491278318997651658106869117839056449644986885454270737246423721194871969778106910540325695144915095665951793550566480752875693022406731307098456823636855505930734402512387565602136962719148921181747382410581673058060694213752620539997364907859384069633938709796926570609461141918080885098258138206452652718514573131239079954553768598280380553422279833153474939490268775554038894838486824230852434102975586602593692199796148893462965752114802632518037446214703997677023006105555046774465938746066927213394364867106;
R[10]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770577146841253006716859050671651194216427324151852519691032985088607556505151543216944595795796979507321307972496371515043736824526805521145902840578101662905565657470123075981047119535954824270350569510972958522006594592222195373586524650066147204783218845089299672610460152208032041871122995529937091173067542373540673959967865756150032833391312788244701752289126137237638430800910743368506691210016277400415940304687529495463097575203297658615017949538388928247493943257052513890208321150256066847624732058430599422385503308274431138014274193886272307171673208271690921344539156057306499691298763787755824024714903894453408818784455871254467523827946217188991864018641519215515812201898530;
R[11]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770577146841253006716859050671651242074967803215427862052218139313921459498489560711432190865931790826813053658749787612410757884306883841178783355085511103376449297413748602098600411371519896577503220114810835088571494690897939653762930109632858014598857622557149784458348534935596538082151858552199925907223007751013012981232062603836861534584740159494518015086093586279610426092064029854509524665974274754758656922506475143339887801310058934563030724831914680347189571212567168207120819070090014898934447950187115967003881234269910936618066013263902880470495055655726960496384256125746307520984938133514767885993152796504772239334252063845824004526655018718621351876771242234487150362108450;
R[12]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770577146844656387931809647169194031097842564863688708668282928215194353203274973249964507359616765307549012600366109823313748675153935594579397233076546247526379596538838003404866853941540927543791411120123524808649632201748086011755784882819343511078009050146836430117020445385192449178734307384452633554383340237951677272739100538625402455777060963823640647463073417310081771555590587377451329641713390103791308009783742779070333077069458785379145697910107378052184344616623554202065766936622649727707703150278031651793553886997997672440171139457678770859268868472922342328548896565508129339296319190084827224737920422202416459396626145062901560977657367719256641665552020970233124586922530;
R[13]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460436004455500951133535289977962086482813396623742845387405627396667627003888389847663839254612124751246866695494814846981868481839718103862091948852888606926691384013541689660301117565871615654878948164851830808092541324006725202275170220713405020212330671269703161745525937500469247311008172458273578169433120538402635389024425591338120000138715847955772368627691804238130967992038202739210609685841959804981690817054523159044664121652644044215815940327583419251959509941577781087052215558617912831229603838868339930848565842369950274061978184713725617839794651710865306928161851241961154578863894436302034546224437698091167810031881631285408211131541908407896000822989320668976031407429445100066;
R[14]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460439761126785901079117762509515395512153994510474385781356158826256150431744019643121246522469170410910627958098096812201302437120632600791487210392633164134602897344129868363444960065932787245547945334676577570590262895484015118414978887810483373385213284787914905134344366798113499369369693190735999125908436080316067719474820596628910659937389028824068100756319597500781586365356840820399189967539269821050050769394965562515812600162604518743692809269804807738144443041516172845690189395686383179417198160593659498625064028092001169722132214537890043497402675179831982526826730462897848617750745139825135338137370029748087669192794888966875647539543589213119514758348256687828882569215093121570;
R[15]<=2560'd57773774597272069865343387443957577157171419115330751726028671677111126571881120180076725499374404477624141084618576618988030561947118405339958765121562973059445710653955943953211226048191052124449808868339360095192249762676527520569677744213363790990162129253519361892866462809135601927043196658611136009619674116096322052327748488824140232475572928196407914842093951897404685369893814664667825221211016523699444492249710401582879724456311794026059032845368918437794556567726287496242011783715291691427174666100556735107936946864320723887784987310607180173296643042917919733827940469031872400732466204883710281366993742979328998463584949517348025201300038563553787909474198250214033598292147213024894888214018348547848691931031742993876569773166584526005545580833677858;
R[16]<=2560'd57773361470875804093833019566451488029810786959545174181716649553466660748833806846972465752516924522999249499874769953927742992076926484267667269471714596692472904002995130036422065131958356176079700514940058214216446728287604318129842854162236295841569953770603035943831572650067133483090163059169929234435271583524343118399160877208007233855965807616970759880682253600515360444611985278515424027616781969039011346954994249708163359862180560651569728049427401239565906715211967880191437940073362885434949951952773504927124322674959759113817614447998967517975541079655512684016067965977845366843036928104618889221032177165512605885870779147713545713597779217845684787190500292725937475449713921996811347103256897184569036317885085838824176500855424621159851289047343650;
R[17]<=2560'd57773361470875804093833019566109674433775464096976142774271424736635792587648861165766805244872608383672477961986805567690923346316645683479232565245606614909389537636457227536738052372524964957608537348177332123493937917282757528339935225431899093034495498560421107396587460745175077183417201728689551322645898607490413446198925652343968175150787639707364078961049466034735249016343639346282227403752287081025271628692030483033795325387793733932908505562006775552856639552758811248536801175876579055938824502275674635125668738374113882171615325879277508011817871972576953256611874614160316403033380995203926213531526204462163939872628959872772830129405947845172299906385375671964859558635406933816238879513613790243207710119154800825233971682898364502157228529720369698;
R[18]<=2560'd57773361369990237240164763066017403884853611448456386255867676658629671397973046024396669717504161779406207433729881804632830388313982112693717344690234112952941704705490473167642925897211836657356168768383279665773847924181611295628614152549340470985191458181115937155024939639275459054007112529367370630635550795826391349507536951238852005848112609170450200589531548069513773231551949686680256985184540808808675484340654693335310425185700011362497442488260733650780454295487466917809308488386891788862786710633625638210361143245910833584062733809301443081269173907082378449633299252001601164058226799463248232030278372762326658420503666360035434943332370449850043493079148391725980814098981652768716440863558012319479466877925739699053421983004807204435176967060464162;
R[19]<=2560'd59571728114694891677698238079748136556057732165180109097654362621880363465268737487360071908961733131164504939192006519823980234891618468029637517931610246730999394990191015120853075450684283843740434658679518057653530228806846836558952237115222639352060483755624671920051920477941884392700064774772255352155450249419754165628463633608862375751395375611644648179659999779039325722497569628997648221886473257622174964710047760446494064604419562100120119276738798257878639216781704934790801796897608292386967630475473192575720453409603653375592246468097255808774559887711900680111132881020770595623469842189686112151659816639268966762871319380123136302717123961260580995683697796195638483651311451102858930104152141504234595323277749127820328946656571294513889609137660450;
R[20]<=2560'd59571753941400006216771902103370816045601972028715787622899576152871784209580395884329639732451681690721204826241716275175276250307392354816321749849389963033638190747429773512875017746615015998028068028973099971845587919751251637660724245741474581988878169270579084774328333318471646743172606864845169022726530830940804808894476511773295499433129154661786035652938976446796270403752673192709301151171653331211659146286483348704835874677797659661436896973964627512297735572123933752333716997198612023827309549802726240861311139322249659007172962260623117036869938192887566273514916699477005804863368367411138578252362682697176909822849972138790004963833524897901326993848610302012006459197142577399356703267532261928150088212478912069378498583626128760472653992678269474;
R[21]<=2560'd57773387196695351780706505306281763924849086410639552313078743576200123017318038823444762673309893740702224549084415660829651178305720719879453644204068600437603116522976601359088293716169880283844329931389804165030773303512590463094051021114826609191183966786829887669850421303369613317080545649717477252735635427662987752532993244140406124893933609911112789673912076938952629598182435710733446588859774301267485833166052078658337297832532490630063200297076878284418742688818655008220831313186393135708429478948905494594174771769722516875272934865527103440169958934313280197494052930541998492868385971945112146561623600840632331772963449252070457666304477218990909911036801708391516619165531233857366789266779092989235653367305753228407773578530318045873449076946772514;
R[22]<=2560'd84855037739454993571676354812050085287620902975521785313648051914687671805555741680075379630184645753606064501268542625670688398569170826904819160369167033581690368634141524232846007690201067183835210862156533647333092486565685604348315718141873669855847825215196623125840228899250310809978044100481125232733424617155914057548455742114858709247379782104309649923967170154452137245294154399769130932711423197697044379939513608507370033880134493682561741162699764779822767829358514893790560310186314284651543783811841425208319755084398727483063751820118055457075008353219109122796308694250193435939324840645802251828763838103325594559365970977718459750683785967146476490662920872517491006987095230907818159640744049733519748277950897712257543576497006446736256324696416802;
R[23]<=2560'd84861649375964315574534703276604848906599343724610112110207857906947313895283423044253936180758442554400416019252901221443715454146489678242932970178078625063688789813374140501473168536885747187172449956087535917152426626059934542303685565884628235870424999475060697094511227702764069292123761917808363076897232550698739546972055242379422498728026497984325439997061605980135048705175467175388344528034510091427070149444538732741170395334615657171930010458608884619431744777237056401943825027465547296924129238512125094104360319462851844596100627443207692591363773757975638976643957015807339679234902817388390619986385563428699513292088636997384125836205330879424183176014210926836172100418551659552887770620749017964850644822342104861299940093626832065245436954634494498;
R[24]<=2560'd57773800423977286631199288167698527425283551472069132515992267034625772758056592628731792675974686172113055831683685587774018553159458732493094908281600846620034756432176949005122154059497817673958975918720683860322946254953703997935441407175043329138400457506631271083418840576970037424985967255116393613351892478351682228223285393639873422626412127685581945262287199940436041096935925477859887686102365272739176599785921608585519187781364394304951755167512585694166330563402125335118914360719196681938222226622886784686685398574786188453559404132217012229120318156560941479976776659956047868907528884816397743774923355449185663341893307650004712280096539471137225344042955237756424188018740342974628325423784776236655561866706258783679791095404379028049162181577679394;
R[25]<=2560'd86660014513199332527338525956260624693852715527042283708600032213176010953371552011717489775079219120796266846697707884762927750683352752182511547733394917588183677217844803845682068743843616621303916913975141258559610146501285186272014604299418773168730938210191341330988390895648904522360187009963925445061218318876709719320931449359948747999285685461742413446120894580288098663719170092192512836768230165079025728312889661182968313546483816946188244649267047924962930276129476569706430741900991413788656825941306582278735878946625565725643594724730068437497830119381134260595467865487712671162357134162070605251203382088183327784201576019656910643433882922222014790354693698915843055834084067178326181765277591804611848613557768124263464470971822435674288525162979874;
R[26]<=2560'd86660040339904447089907176126339298658372385550005500412844907312321895809690773594729787991810126860132749379633350250610523899379677833044574233793795125174668865424858048496836108325384418940790253154761309240566234132550675206618642041830308171867430389161944971336735593916210132022131503530537889276640071219741698132106585619083033078011939152519957903070068979415213717612557968256672928519252437178561013139846494255541335085634657490650874728186597025938793318471802674701438713479970922766770069316053977301031567503364609443192865008274147269627258508942448598478158278572359056728706631591557240080030986537164228163400683759323271928779255009644467443410983305858645561780584692941748688759453146918036906572334709173412634328070033088993272005854515831602;
R[27]<=2560'd86547644233906525683987586255959996178780177997147997872238240032073269924095194978006632401899283121123159986973669782514802806617610392338429356188969010571405452728691543893886078557031259378784701744497890552644424698074255220202923599241055182339369292742282041704193838968282107348722417470510026363729128538109701390388070213211521405608743445275431893536783715770969424151178325263197093878177645772979283183799834511316411771335680431246572852585309424200902827184539073956062131391100994881389148516651124884593556520806061092836269099951461061547986220524484233583170111118780297363967311441660837166650709627727135236239650196250340110051823069280071009638244155378367711833864098072735636665017152485211566547812428152915839720452697845936937640251913020210;
R[28]<=2560'd84854652053934553616298397146624536070538405817058795791924372022941743820520470230941590271712037180602919722013743340454328164096577216058187903529732050798498586634277863102569602142576291516451026515288934382451154787808809327755103774427980792576872258156047822403159640862882035327291064441941101412182420772980914398086519994979424008127860473672084879593065895871789924935146406586154777994941426366353735256351612948067531739489928591117718907137891727967351293934361974090100438830448416227896771334931776106721073589421338727550823563227038486511103420906199040018121767714967660437023136383361959210309570147128873153967453498893275832288057580110472253007465240434725688514733755877197293623892297599257557389657279158212075623668066763231393243529114427938;
R[29]<=2560'd86547203465285291722482633879994214875815498975382692729280487970860287460701414385200255970318623556746334272869381669311096238224468381210547890770423106354435688581003206258407953893488933786378791751915781472531612365244017597544249648277442070230123583307952948019214605531007597840715936387558279604095131424961528662324132312998631503135389959116820519422192572640471630263442010329949258207701526306317463390685335565874054041007597969956740717950506839656760509799215976725775922632727885979057554479034001955848623026512638874018429794958727338960576419281895324545614036925602851291897515804428447176454222114615066182882099044737877142010984915940204950536035299599612153072355618412392530042050399408658175791155816902537636026998207822435892485463037129506;
R[30]<=2560'd86660040339930616723341394790270152571184390368878512106172621765721761786334940882317348557350115981369538283328281307380971933914934572412019315683515460323602683126835711739208266027009483980063056403761789137044299932557788435826725385959496673747324612807970047750311784421496086925726238433309531533625184308966626480117925629871939538614258984676207805307644116444641756444329058617013468027523616568601192605257497789952848450230756953643323492745599653218312302393190581004587989248981335753017744959379788285806784946726533178761221137690711679957573770373013219357439161499594901346473285352103974364907452831783993862459954507223018131790959681413478751892490149539995229508689724957635794938511251978717343928600180224075707355994505089151502967251521450786;
R[31]<=2560'd86660042054983714243434959341365726246495501958022391305058741483538812193193512051140921299861090788630797271441700407132062652736259783848185445206712890924420752261136589925011526371798819243587942597496120514131354469309368529728818924387321812522608260999913810195140623009015812785977759473158622388249885673805556821446548211834368271576699838533418920514493519830693722143502965448998635824699131719201738384309681366426356354838822652438158917655932935060919757430635569367099944752511663786231191592030186867506931887112961013482100795520886875360160209863299745370046711447841909152093770400346771215625321707800411605177606495687822059067536051707443892351518632099274447971843916585869092640814524572477509810661777545549210451381612593390039786637906621218;
R[32]<=2560'd86660042054985349471078990978866873383091253928810700187133553067155743843200631518745500737262686373512211606600663811041295368135079097879957475673853053530199190497913877777104499248986550134855620124242746994467879621536033113987131746722757912166507160203623231330756025300266536996397491376234064128643431893500187293052189737704638924212782143797859339400465394492457790930067517994976831619134652290051505460921375358806983168229107537861536530742276403770391883848554804535534693160013240732440632153859148089486517665037450505671347659432791099686377303995985548588682448883339361870345335605661918560385387843864809000146831847049702609616071925845801506719456126904210381434281977166952342923476996665132398827404022965848883340509063816712299970021253395234;
R[33]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190657397828370163498723164913685864674604617611832076045901993997060241425768530503295962087441676672526096593656057675529032768822325345317787245001546690868033476231727400250427677543031936970352614325898729171163338123081017573164312718840866067197200331696042156170747968491170799849874707365393818741831059505494822523773896582561035147031496004120688104659795679187778441920133657501682062924203244353197531261743320598589302545276603401799649678068001091681851430885058924638923118150984079006652750602731440828566189645072263058271840641485688748303943623249718046003044544140568077720876050658336538857831623516903268377480886996635707503599997644554141416005752978621187735647620856754978;
R[34]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190657397828369292234014971812035646943822631590102383456438229367811963837047098782979556255159641393552570655490129934526296865439669799244866722657119836841084276889479123542952554282470385022152274795495621957013480389299800462920665170810699985243856780458223868360843374778163127160565177397070711106698505592927449940797414710756915765368760968703584625403297349013717095289817551422575089049273787086692426910765102735892019283623395926173089909278744886942519602601434478719990081749655260981101645184836029094194050228683761617612029284741559524076190765264426240417536067503343686247937430731350027266912223302643804182428842464628197365534632658852519579838334407258754467459055035298611;
R[35]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655778510202194070040161637417840900771471126594280959895654037703205549443451705331734426120302890038027626411650512251466303380351849959568248800570872694192159108235665223117982692034753284865807005281431807393147686334592744165370486019114791506275256411762253343999288511676827592420567772128568766785968295406151420415790795729285100265489881441019662675831910331779263387009743619300066762956453000221421940406872330379884283866249880684697352142141649249313444657200737042199370064025123557634707548023007465950754730725955012173166315959801014856087170437732410772188639969214737505676321789356282994820385685133205978391940304285333464365761427757983256176804850455244240309057696563;
R[36]<=2560'd86660042054985355860247144599026105825370384862450713255366273309420535690531809473154932743249057817960235194511538639483657108702584117594483549706751669993070060604135443235778016595193572530866041647824603335615946624991648011946306688776333337586893825044884325836406083916308991286584354641722301564662847016434433334374352514722325555239091441758688041587303661435674280792999912751013003971620549902391436174574767265090172318172955380343109096374320803588016649193108722850005635171263569617912065571393519190174976399184967855484254137357704749615382996489953129488088395423301599118179602198627141036077497085833835722511209144738720831045174562152776435381936900858090572942256301072510553897862018364809863945259366808264623663376585822018502469380100797235;
R[37]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653889656877323188571555612547409708236825627004531490970559363074718354930358376364126985645716118612110964145874307956049559112198443894452957986659319575107696609302942473597942669599872016311265148867229023005173142254772751930569000003825840204532248012810675726609370890294128222379096465142468906017735078404235596041513610336176403120317186255558238468077373612703401185314589231420607657466201681264232437405144331537838648832357875437908038388363570647727130423233122483543469278939969751277342360697257895316307984859161079954388547057487937484074020261551183868504359662321516224398030541164744774538941282045048615640224802838567082354516877311311343561195861857178935981929449861939;
R[38]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531206999195592058631515169666085870834112215180850712390801272940727870457721771369136713814219035557895172422339617333997389407243558208709928066636020987871570716482981243002303478933367314551356367101769105652767502163755149642053652315807525023245392905916975246841618000391795168654740183356848483491110660055349977867276867265485211830769984595523755878866113883992969540578929834217104591833860336645959151897799803041712681738528943294636731407835904570705479361248817178876443015977666559901284481937915382242958028520070787908597641591323338589686182499710885422517499770322137144442249643539449574790018369186665038480849875047590012558038448088104105999938940218063493060079969658482144051;
R[39]<=2560'd86660042054985355860247144599026105825449969542042632900029023092504966583652700713258564343580945446434503036217230676100177214570808110423548599902692897236229713371170339198121667546392903080238522631668676183078894976247648345234481740751658215289813668522080149862384027219361491548816237799294768246870093499258909754380271744639050254643749180999996873876795430651270530153152125106786698856905484544072267301506091070179026141025424573837248111327709615233682349410074304490502489993043075809560734034023659792066176487668779371481291609180005771713020838670742115618772734180585023102026930464068158579812052234981384414556401660094492808766172282087665252745720022154211553524721713288312055839787382764257214440802956844999141290532693954263320443993017496371;
R[40]<=2560'd86660042054985355860247145999094595491657999583195198385710377805869607512396466731678987761437164972739107030858391033238520402439539630334889622473537769223704632270839317187942177018404210977727094424850787920253479721927428136085572251020596373980629949971442245146379685705449409672537304522564597712924107208958314208419091156163789979313585724578363181082249707468828388402274707269788218623638066568898142327029629448327660211516401922854060996102493235449118519130297447045948581186117849278097339921048144617437041912330332475395504008331440676802824937174923867845712331137281204425048898848456099691225611922418826310914538946403218352038094748234235621365429995829856841135583715497922842648762513492360395868381273425084582397999893444004480391874140648243;
R[41]<=2560'd86660042054985355860247144599026105825370384862450713255366273379364933412339842983667055047579406082263711460100440995334376837721761848840631372329508764203044248349919802125093496978063216703683188686996590615444302333877479206426108392116004896307220607487467785168437029651672268191249678499342200570378707334526834768521380778250803137546874274698295843841074750359029668018132410204531675088437274707169953899582139330462851165060769364792714018188986665353698532431930660166289366972965911796335904748989053243367277052308974685592458146172124511779449724931157260177656609321916834440369489465644343841424174051710438391100523786656589450857221135900635791397372221889590987958326028960106638809298239411399053972428134495899663596034637604737731530175510950707;
R[42]<=2560'd86660042054985355860247144599026105825370384862450713255366273313808258124961949203538259139998459702056690386339957481819378899749425672159066314793457451577240781638063008135621124236601545533106135810918564561510481750284939662457173114619262226107534778546517588708549864344255077008336752270680402330667102514093759456736893536255318470465215786095801727285610237541274840831226346291160890977179416461971452103978732218562674825598002331744350861507771502234248922500679685876761707952789841735843590356453424711021690306577722269957306366667617521910324448240289929818976416294594792544912317039349286350001951742033091445988279211328987374403734985852959453466087757380391244541222510046771399578014182344042589037074529554947025534796527809710348910537888445235;
R[43]<=2560'd86660042054985355860247144599026105825370384862470473498900560383790969233441429082679984810915182786798554000589142097913456665368701439641228964520369299944441966372142316836296012441426454755047847902133710679288449747723865415630375009040572882694667339045376782776900775377336546142151578099265244474344423257483945124601322886754020219466213606640849796661959172891400980485054038055082569629271221272748396409731256653140007087843266726902800804163647533299589847174360138852882496309338560180578725218191789624918481747782649190529603761616806285352943683587575505893915895564067541362571991386245377393385684093230353337641840168283962559436056695275959262571679457013796970412981947011218633499309393101149130729914652462691915708444771501502375625706475565875;
R[44]<=2560'd86660042054985355860247144599026105825370384862470478022761271364532961295257704729221021131612876770568028465369627106275238964448085990526283000209666828557148346999043649916562142048044789654538224907986114647718881169296998646297860381251367123775011475464341201410632095235216534223447957421663158619323567892975855817761605800733923137795239453552729717742211564987090535939419737951382539239862305893331275251186747432609265153679532732664258623524602518288937567862975673841714290405361197961318294155092667997432251158662727655910938819925580958746769581351758008426699217326433714124105112264325629694703848473695649774549596203759666456702441016969602176716288397897292071638156591009685350146744363269211632687510518315374964705984813915055130378960215683891;
R[45]<=2560'd86660042054985355860247144599026105825370384862450713274211128025582489645378578319359534944713072904378179078903205061258955086550259735056424359365807955694828947394988227746318288296013831340056171385161032690446591086833733016052598612922586478096519079627263377138180034100981624266389374193185674290954278371436418280041886491533662734669332332843602156578019197760209213695048587015404418379889032054199514946501514280483504547551688657794996230414894643074193333402105889151886121777962929599874127795621299076530964881475722283225284633189595220600366941235274718933372591375418800286316537973432950665001100806337831008952117972188780043702087134290044747031669105036035860861870819030368366053525311671557114886335727124301323014007162950885173638800361075507;
R[46]<=2560'd86660042054985355860247144599026105825370384867490805865641025949292390543496542608523677042732505848431334203470616109546754390498819825304410010157883509087011339056074816876439722622183531849093964254660698277164375661648826159886665179276365371593709108878499840102591708420057386504341744840850245188437196951956872157149438257289537378380712632380707195147273599421874549154142470815487018034175937668226408235301960324270534547946968069076394385630547675872100999215476757991762832086186350851553094119266118993156366870451846785516175551707000139511575659382588108648804839694878211496723776144920421227951543153507797380487212783117439520767903005458152049019287194550619050955583143923030579993844353335724763722253481270980688773063561467073665335192823477043;
R[47]<=2560'd86660042054985355860247144599026105825370384943408430996629323382492495282544801194201851668714806843852744017366940954206200390443704160354779651618464754910635216163852899837414858143995145742208850515986112831337224936263793528561737911572920611443483107843901638810984096480072664422267815555037890594797856123363715088247129490780720765788864730026535740616607630693950827787237217014825359952846254007398458708863063677847574531545788037542670095583546841426566795013229422231390425547814050846531832256637360966494161967215896236077316683277200747917986919914283282408846602797433286434172155988982326018770133863073202957289477562819910090832348621666833300117729944133716148863683519822875662727759964116161129879766580796007493815022778056171230519273022763827;
R[48]<=2560'd86660042054985355860247144599027524485315178286342881503313359107810210882286758420859735697677702715371224890610223535319203454168840169112673762386350707273111350432092416304987347201827089904471491364658274077861817454089395882524183094291436050836282680183711760696597995966985593914721487986095937378218087337733653572617363580878920207084070009259039877067514778625774367786200657459040548434018303378217066407130043588814946903441909503802525058005524626821660779172415231756529639535750313109758197850846896479395580784424784713625376513136954627422151127676269690724852166141113423351662884680657114737890860980501209577442373198134926068421224862036953346833978796160049354664362283794907694010061503455531824797591035990127798363773683552556536385966336848691;
R[49]<=2560'd86660042054985355860247144599027524506962230641077776001648326611426741685203825183219895866240491356579364002356310457530253206754002034201795084953760802861847321973770594245467025372329167061525642166234772030790923171770597914075954245251283042568345438630306915012870076946752784034073795315032882164432373955049482305821989331497146609125064748101258209444389814720368290319437971840993039842318424156272479663736966056321906409465694773634595308531499880158292938803971613789213477994804496055463425468192591475648377098696470188963804053865660514586640093550548203411518030347482601235432633149441912027233402039771011016136615960318880495174580731092324094465408519040656680315091298000873121178135433015039256990662494407219162694537064275278374643008760132403;
R[50]<=2560'd86660042054985355860247144599026105847101997153654925205710892427117570098319315596922880966436658556203602568488338170605979333380608179451700721505915991930054063847787019275281673606709554753470797273430339037216304662475378842362780203642370176966883101149800876162682929584475535753010433387703693358721346321035763267034940356925387000284263852583348623457456026286321765281183052856146302354936692736184072173933610663857115382750266188826627324985550079944329002456042464968755635736407285281646715129608085335038708070275193893804650032321334641530685827152357605974854374646979487930198873827595953867897952437942068739996765475422648470884018171574772717425157514903854447332351540395119680025262722675448350930966917020537781433578795032738975825158611350323;
R[51]<=2560'd86660042054985355860247144604495123384860933153382920155216575593502789486967465264227853012545893953269379804173428824746731646092879389397345441214307147369601249388898420866646979295832034206543994916270041296030163502357390706978124357888729507742824898009660153076811353570442906386252642132363704161150990411839345736769691335259632661407369119069733095904493859186660373639578276272661163412799110609197763778548570988250243956641048463053518528351283031585666048644938172751595020307631735558838704044023863121331103493391343487128623761335493384284380236015442734635786430243668498849295435071838711638336800105877490922097339489918282868315729922358719226896978518719485605035331404210504104529273789977424105193141238498647336174109196122448174399984416011059;
R[52]<=2560'd86660042054986991463805219899333553356456294087975538600474899124939883873852140346898673950175484734079463223189413310560910822457714413521657952037128645427440649915636808286721332995644758388077729815813113589675846957328274038199215589030792138397033995072804616843467602630128790390802193732825610428263833916415447683995523705308066239206226999073244731865848394332097612273973313519668736175493304099779801208710704096063921661834108172807280758731072338396611544248795578697631218887496928827811482497101076342881260008470924937979355467653601834332803826008580338515874911443543031784814507444436728334860296965371920481832422506841410554375371111575557131789861513575463441223075141977388832547188933489794763776361427705968815552073106618400083705955089593139;
R[53]<=2560'd86660042054986991463805219893864535818617753983843458711239995000166463410691050226424640965390937583620509999166887975386495656051557951067473704689088700790425229100032446501941656230427710592509771301369924363378125024648905597026395882523611836979513978352029282219226912677707927958154458689806896236220049042154549908614898478393267381741628623672631667399262893511034890040314930328049640529410515007244328798690970184573107682285322088446856844648762309041650930132398087020475850387101119967344844681436563728623247868885576716287782633429805590421808804993549269743024809139209312231417397414810890443137748042645626721579992907423733366837283923276772470335799340962712143880758818951006041834086288958174774794024735270057469042290345621081466780966655832883;
R[54]<=2560'd86660042054985355860247144599026111387384492907707816508030576582809955086093770473639743009215524073147139389162198128531331119567814373080521468347892160076526446537214356146979136778415577692839761748384987107825904465224524085871578225816709697912033426558106741762816332083837644462597280168705880488600075718067639077817912973437930030548867433537337033799966744512189604075349853968188374392900595145268188272855616970093546179583569361216741486711476729841546911592578882293200115566397109995447951432096322613839536586831820687622558547122075673933926602077743939834559815783789862825371785120486070110491353156011248671307594540491744249915162375342339296018194387121746917033812099203655543845194742978772465202081374464788743159640659153893502093655746491187;
R[55]<=2560'd86660042061290703812090662096206953526977180103761846843533160057564913533641316529548496579156688830755124329601510661902801047760447210681665988247260777465487606824949932595372924642149443518627106578998788849605093181469876554280374573284784700299416528530079985264839193049590472130274831951577290772998277167072280606438764559573910660447587892763065222571527421308907956040737989018421734665043409995365839191289769661585241994752983683066727102788997129001486073355093758404534685433402527420169979543007055044889312203965162915823327398837670992921749413665310253174612373087666885865062057109561537193768845469546789032153782322884708444665494402461071138206028322096155904012922279269289564443437046260008441564542008038837432609017077848413277335270869644083;
R[56]<=2560'd86660042054985356259661909176670921900115671537150718549270095808602670518788928195169449956380894487600080751486788342617758245904200992557493550791932161484308035803435780493991116927045874698677603486310549199463769060127472676929857317176612893656063014768373840337324383339618783424429594887890233992884772378946005328782081878853296665804478423301641872293730868576259170384555757057537839257819690251970432187068951483597327585514916505539831366587965148552850577021937415947968680466418474225834801640513670757040475024349442711756535462211883383994090760076400791901077856248753668439177350641282271085223195398786206816599079760612456305843168192105475398161264527086678505806462632499217700732930082085318372277054637730683392438148624777202709706891502760755;
R[57]<=2560'd86660042054985355860252879279559778961087294531968257063724679241628012323114888132273903295990674863046123341897961833080183342937132613171031102060768080241827386971198245589566576123129483677216594685414317703711532600789893343737014630818446589617919513375000112390020437295901385048634061802198815177529635876109444704902548996381388321640935511219127909470443392651278349485780206812366966945686557360670887503147811313877634767086162804086027575158774564167259667568720575416103226998746804926358167376219354288828678060705500316287378994075039513296937605029108578423838500439226964685175153356965693134495516538805021541726489637879351885808211500055129422641272967894666858597989158210420909386179098055717663291544007946404210124201081239883368011905776169779;
R[58]<=2560'd86660042155872558317473476393956806370006731699731253985208197846010288411345225679579996108018080512303140477682782058501029414276750142769240773319352283307532336251034764920748548727983268531417850737167659011810345720266418825328787953469248244737426423747497510714248573991834117154992341832256583937645825481032132361139168968619215193172805289827615271606713750247327720680683147849334858061898232072953145071514886973513541726206369765042542031712209836605854604784077389073871556150287037640114001242313642722430433731938148171270876078792327541646904091733744988891997001743160383150450796248638961927430879221377780893503367409198723691454358956715284061884594079762731951380485463231996473959243293848677835950508036992344012393661873842403658677160101753651;
R[59]<=2560'd86660042055011525518644808357159509687291433515085964417039928896126589523036157030202254624748351347726032316177712983415544815224926344480181451280092230480513733731852473090894348689112160045452570364983360406450457174953985408887907607321656775588617371753084710375378877178011321580925218561517507530380449443033441978121556865986133151210082691428903715907926746646488983199534555706911776629436604729625426845641605609387902608117295416122796081883574681407109470063003396778576422726980178113391364287138922140614816627127566105128471889545984170149177091707221802971952211709231557873960703944370540445142069041198299026618222883561103774516458185755624837808775179378085704302382847864104624506194896261342230005710652863813058352810289416753129021733491389235;
R[60]<=2560'd86660042061709418700254420070364753889614508357520476624721847807459521337465306055389381869949376590007380915637880869426450037489117619135789536092530397393851945932863022784825021387527396467559900916438545666252329053036781639038463359581704323711559190413038180880636256561073128020105037350598327671619805554752651591679236676555929692944556941839183913375307598826956062552907148929684487485586095053206010103874629023429709003614237620274158062630924146955184024662835353185610528585105702830476895914802121256876289461022881976696866118527709748142146797670490009332908599397334193689830455001318338486271207303318949634446854851412072834764067280890678919137492267658627226670678203799482992627192653923657606018274089623855056897318758379734360346225072616243;
R[61]<=2560'd86660042061684788434908905394581954282049706344425075286964609985642652802841224492871943418896032920217549067834880581168342327028364026700841481509562565424444504679750194453926303611173663643870951586117099927157088254226142055044924940080892482010876829113501699527993612513785354736727224336428738218836522903515473845347614013102648912334529848578521941485655230499593292233105051707831003364176168518680666868929309106955468830138409697890405768926037839380741507899051255828496564543604864800534136155758708991589921175442987352028988051086685076336849536761795789670665990635151958961997599890768867165253672411716233320894599462567959509898835662237083481420850656800581906291520653850831730768528997330294445394728776131916381729126748890625332872406681989939;
R[62]<=2560'd86660043776739430959049564356418068482798466267026363645601927613655931042305459210632621960045613066769626593953648692947322220930649655467775417323791225067833944398209637963838618216928797479491032369568743993350634981293284067391937476790979468979978962684723201343643735098506263324123787609210878912941327632287396887860931845872967156706196488095078673188039453156455307014089082197659108601219198261739905764833834663395952373891932466972639002788457767609981403853284278662892499114008624106716597183104282282056465016295469538830356531480417950311075682933737402319863163268435928323948760288777599869566816077748920891144742944538657102139917151964715192950054777411601410011529147713326102333381581204182035410436375916063186697780663278715230165802041946931;
R[63]<=2560'd113741306912222916102515745629827062024192846773927718299790363274151204559617680307635052003802028957875899325639540199376878760337092314724543667534944988169781894723172922937953579341649351582081891973233548183540508808131879053295095116121399567394249309717907159171800997128998960298614170432743606107529604609252205846070857375295591077590224406238376339356905491272859010413650985127707959827791231728202206490056528592517276373696812171830955169620102624587275029547663361542814339649378827065888128641680066336429917062427401531388847564651748485690726477909204471635618757351730018378467634390693169402235337565915335390789898219718563461991448867360983494256492174345159061931083291053766698616648565237509751676533037825122619104559483733742666533982811927347;
R[64]<=2560'd86660042054985356259662291307887107396128118975143391241736401332616567217132706008379085197971092225091794459131020786618339251093417034592598131674106841641838066241666930693489942136868867164452742704985300188312826851427890339833782054782468361844056237456371254762593063893246375696235840959523580585718604936108734862445531279209409324722263224928230836226165077729707834824289407046228829047869907569866137238683554422711910436635649786615326669203664097441724607625170472070983221933721735247090656505859367163473587248713567777977045979324762921016886829477407717417150343450162779919193827212598676872341666921873070558490445669464604127110581560391151121248341915635229773655737033433064079576328307468212566400469204734422694491056853570533748968307201094451;
R[65]<=2560'd86660042054985355885302346157210501844775657980102160230944711620244891574782170445457337435667824447536769870527047746072772298950173304770324538343618175406629605672691825396395552723433292116446955230933563664624532058050881568273474823271552534066877326005776170913892097980344949350461930991226400763110996940568016431404869062280821105230887713921476840664890142767459646825802534072828715111848518660335137271485924097614897905361379214277415776222549491868944530959290096060098504770398312182178894899105877162560741510405556782520067034420383360672449845755753442945240732068536820397947655991897628360200889698728701112301663438875590596484126464095259526015836493616443250786031307126692549331786140629771966058388813926783172721464675855753649771304444965683;
R[66]<=2560'd86772439875643829910398925496118397644980468243653935060421426429664515755318921277076319127852733209416501908299711696988293155254046791612362417364905859213671160076037874792454705424030141217605867752265571596673279091388578242339904622948807226508094172374206979659828816627040065658386017964171778203595418699048120666526273722179861250085521321631827114139636645351247058508734844328660483161103400939613095104316402725829987722071490565232703220131471519471833742619738063736289713065860285790535071803837714794729670655540030570216515072212301518457315840292160111705453505079395323573524695057602471633360235863757830713292934803046751506336292998519798034545184646627532574055541187515475645427487733407338401255389523827162851798144718621981054449981156700979;
R[67]<=2560'd86660042054985458087035474402317333893402413326148309711117877882198346765958918604498883896507696349201493982411126336264983311120353329780628280970259522076585839190161340196052780052272702927357595588144135085971782012684663860040659695373083628936331308657386616372736207541477925778905961528594554356131418295754555260146073787186587749870047183836210510475546928155366597090915605920686847072020595420598586263036594295558097469765185278054424251982078462968110031641042136147707119349572170574474479463774153810344382224282566105999663074957271343742155430541308348270187540261280617727712473453207825173904415429569151288666051404525816947021551567824014165303694515042605634583345133962460045887232992844557403372643903270488555993541902552633377734498691789619;
R[68]<=2560'd115433884244441914755544033004845702060129319655254954636544497884684051583106755871158390810372215853380970608756650521416183995433525440994104438595399282130233703793830956420353798466302025463956049202229838454074693887659010366504078669613136436235580922066392902297560067525071717831955055077265766172131253511771424446119109971706160633869443482446653535600584880591978119114706555859493649384918317176053472624900862214219787646542041300985919338378828160265584788822067836393431602800347415109408073047927101757206828229614490020541130336169572949714558359200679620043118713202427579325246095819772539303511437382544593094250094260060501326831077326944427596161439949265494841922048010288207792184670630323691940858218424388644097573714993642159546973423173579571;
R[69]<=2560'd115539670428615600854643003180107845207537251807109916959732824582815566427271395598547917968864052544793495271479965553688657493680707915504256453562814814528764779213603146567188314902671688873704715581623206600089056958493805583199900777686826911379607969289809338350955768423324414095483759172663231294763466140149232149521791089033449641457999281042250281842277970596425390052440037577276963361436278081065153963360882902132244271911295828693377491363199281809848481364146097597738230057190829187580323238688326697363967124141235999340550032970368346837349714949532798935931468183337206968590851195012267052177956373537295113380167334668689875254952154508246410313055168774522490398770138110060514982450428959371808573796503773431888037003914383980739999172400460595;
R[70]<=2560'd88465018822450516566516897040131128408816384258197055583990176216686477470385370003621016644500249789371797109528084905006900751745624425949615908663946453703242100018982957413131577802895784847597087230268427118699766740439322277514110383844563647734773164824272915508756613062195675622890233367432279283083085419530208290818062108440640030640428759748922028594632356258200438266006749952874221193225130195536651237454981467612240613469685944781973896220742725287949990298840742252805568207174638651062710709059300610408109035384781074283799409500984450740885940460685907050138570707760196335510137696179632695217423968404565979044420463618092642358165838716817111870430613006512822765288749008145716514000045614592383629683616788115758990863978296358059321242357543731;
R[71]<=2560'd86772853103345916837346171046543093612277487282210449760258829378529702122627592600945798700767238234642510743069547913744827939432382791101947639379330579493455350259506643304783041685422067580176592658078529580032018458678904275980890868995643142066568373746826726119462364420381808853944874233467748169486267065731712377268598841991687238001512177199057803860643671163718955167490691469905673838665826197518929478764577362031340784773721992129964060395053934854466994102806527767249491025855903969578238283646303594712524274158477855760484397457622333609950670220171989684426139581368104585328069295151173431262105032957322796638986095926593965863552997601419274785774594943717503942632020494499642253310261930603069458225876940701839313309784900960154413890334372659;
R[72]<=2560'd88458847961286593167586226609893460958720097506648808405713204722629120778463442721518952812420090890841436943606901374959230399889008643794754441389226150310001042724382020728970456775761892270368502888426454685644638801973023570803934373397208636922408726576874726566937248758211374880677894757815368992894624330278529725462820831765634588183852126291221659255478065216234023077356417880213390529624413724351110640890119861223924788930276561942604988408308097775218561932252421346349514346903456813526499292278184437378221751362955756047027611972226306643760907229735414419198057581988809996000078088642149349059935853989695728427486294428278509551647620883268842474432046037065570917242873907852383847893016385740220518285339694132229022691702557433345525409731785523;
R[73]<=2560'd88458434626813845760385081100673656115354865026685256443379080191129654180354548134697886455307814339074762265986201557313193278218803681810795960809643589764979270411579528337144758374546580327395197240779562147395696332979946926514586812151806826595674169909467070013556457990123073721590723461810810556114495399775155241687686308197047117485552765944453710482975869719850518563021500195142752937966046517676976068176842234621519392573682186856185494619306685369618213145239320360397891284647266821866438343616703927611165614151772573755600399513650227868915560045888478287178976106837505837079812932979785064707687100102581692874605726911060332628134814480451521446600574048825448803418858975577637392074241755828835027989774450130973888309188175418921914057916363571;
R[74]<=2560'd115546307791337021810780710264363309586168621823507030534041888172833681207658152146166617857106097449903827982813714985901657893079269582988416713806073451484736686320212060248346391874255004003930999462437265457869584657266525687728344287593003326928159168579087645391908330198872592019616990057629039958439426446964578408561275762289250530717223718744823844775385604513924304526691008009485981638067985493527095413455493497821837007212068540488733082189801394910079994557208587339651915639641167655114128598657904071892110564564885259153206337917204218575636306632015687598601973939710220487803863248214178673164918084337336493658013995404596291125132701857954961043920002214057023974882173345751937889938689624805328144370959448542637918490664078508519772922559279923;
R[75]<=2560'd115546281964213288949324523725287038195812116436194190817975462262962644549633684176970772107285521921853065353401622324031650787026003469644394778121857159031569774892538120014661163723246837362208398052341150453546324960877193483280761124841687127378656528034096471565569174493655754187766946457586601008543110879275314694001147669314969676594712033102445336328052568794062091665789606618307509933059211516862228307088751444735584836066907845955699585503725335007111528534040691636316732917269007703572467720294644127583628097987883082356590946032776496273502373153133487064665797871116195662423460097268323936011287266556336251668015610467698033781458144388223088809393039768083475483537709257636565865898777422770538083273404865063148989794961586560187796737659974451;
R[76]<=2560'd115546695191496654577102573731276422593524994144741432958744638491782414474052740259893258282697512219741469268071001186629828487915473188561862396669655586644328922486121088919745184815226049629075064442977145140428397715499793282412145348221189325762355799621136702917927498877264818473900579177218367891041531346334006821636453025939521075987392287214770828027633543137147285822931547851468594658722011516174150089642091204563832960417873122410822211227604952912257390750204118638552246599322293501471574140859851010051459605426027009701203345490370181512266884265417980904864769129107467950891210615951861097221442703293319741740303486449079755244239345786998859315548587104382585857547479040827050629888791316924405404447321727653849374790617947307277971290640823091;
R[77]<=2560'd115440909108233069408532241032113690959029811735111577758859172800590682417351064641362718309402891722622434518926197892364270270351109678228120185681647338195171722347122818263978535131475036768299642782889482803709288365985545758514160173055456087517526748410919018361618552801494117802495118967413886682183090921937540812239499074019358920293060296805446624445396935781041559095324948441997386208570491463599045154986825113085645144717970545231351949789382564148863773845118920936562958808926925133392017094164704147007098170147580093353125805351623606281527705619942455700457079108439395871575030598096583958864254931006904656227193129151814939674435906390078867767231564172552243389848372749252810709366572539478083578200125297312527847478840487284135115113196892979;
R[78]<=2560'd115546722739561759969462250653374030936717674404759527230838407338386477947148468341457112550273291040780727707754204862061197411877253444857409417997011239732541484812239329959179914077275805698136295956140834589329686685719319716644522387865054752713945459234437308020983374994711175578297037005386304405000992209190982766831093824469451740223445438738636299829112645913130121151622852260971418523529298082725498604763769974599882516526441889201355081847951150286244329594275447823440524057183614383429963948914108492600426719860863600664922414781143981222059815408681271154605470586668979399266590901347670015466733512744392957287687852145415490168768627294616011053298330830524785981363038884641561803956973219404373223499811821368282624503114299528529967501108523827;
R[79]<=2560'd115546722739955838201736017003508257434755359998303641069551094497676565616142015403273461271889747252964039748628340121821880065251981710572826427443031949752678347249141731180748785257762203343334725748464712928306844004919169512435644332311121632789433343832090879639707579241217630013152629015581005944983620500135741693953834502714004888934545310889017470340225562701129951469677676606324902878992653177207066746190943034230152855037836533111637183381049977195623297187597202496613717709615106482101053132796062948744970311938163700178155937763044354733757122309895303843729627463977421679299464042595742117312110743043371591936732248115285708226068981438552579697030843162071766053976267316108554717087290930992345882950436909717750485501463653624447803889628164915;
R[80]<=2560'd115546722639094907626661245737804909532591966489781953084988522520572222864845856601620043491769758046278638297795353737255794604240466418343264751725281306521479364581765221306299608273170082722876331525555328207626501762453420469461543977334640100656643504890236585964141730521417102813553644177418191268038085420616886341725459427834928812510531129022674912771599794289563273028549085194336603310660025998747138877660475630809890762328290397353389498319669392973592640919974637355747712030718785870909130775201301094332338858540254644848166304599309797193301197132738002109096458674974852587276715224521188178491869206966392523707450311227607053647274219020873779213780553359525944119269601041375508583437066346292772058810941534049920698781146177247548220920000885555;
R[81]<=2560'd86772880651411118042356841401889421067330502551073696255335045086054605835356755382423693666379619922014936694799007400969445752373298193184674309332317308841794651098074706250031436859901107108473771182763113383727106460607201688663867874338586330943876970152824672763815484928233464655414222127645441452300120575414264003196335530427134053517372567682451079334348756323890519344323877843221300835198017266043354492921016106168743948808404961163608727732044030608428793478581220306846575626053874787450662937429900890155094163853787986100302283579730910700146259228824742549713000833937261179966475673914433062565669463281375616531378313949841745352354885005188756673977057621280339987227834508003209422679253782388712785861428676063871268925711104540347082415644291891;
R[82]<=2560'd115546722739980474480329526131692994171050579650247833373191615019254092427119445517310176276560891546743632092093093285297460471957598038380505136090695016110329231196681510319730670248312049778508711846805380962608222186120750590090759019560260036747727992059516667020894636350785014329245056643182486752505467281333498880213206581423687913280416709984382189596263465577943307389727131207841117367794028895674942581888499221272597476951112171070666938704147273405896324892528741294379418578395477719707866965282037934307401729339777463824313985428628216415009830348111539661592359085508868347034694030245697405022808567680052191597023986699605860803454159727551415786112431110464776622394206673275619777240706882131723136359522760392695723210934243806690037728191656755;
R[83]<=2560'd115546722632789559698307003600344956711552730380179684853867416640160677182585550402986558765102798430348498655302975974935889900171084812923433740653861655268576435497148481088905145795576118889098774356629885266987004743029065098611226164816719865701576199261614524345651292095177683408748358318177142988163880406505090030134346665875841569263558049920592589856309966928592991706651740118132603422198258207371392174339764892969209110016976108402852050416322714961852885822972098922305644467452266190343496856744582152305123538631248766425828071743637187810570657567134675984338450310528971503699837649795379077154365649158415770594409409405494930755291645012006958079302371752498118743236523765970167093120708980446106324188562886137861622536529566493538597792484897587;
R[84]<=2560'd115546722739980474480329526132034807767160513150230760675695873007655051263892547225604825473704876993313810209424888846869891899021097237122688469462902129448370901689052524657127397382164174266815572343777905027632394631168336019187767226608785058710162320946983857242986550854507095624842170426887561307795368280266674681447719904573561057305481797246622313270138006655522757633455941218644254198720074123103889468779781616381602035368768444375688870611228938057639185293321615650308473594546678547903954356191763530937084412744963914688013710399778657937251902022891184223941217750479217410692210184618722441273893761452411438952505388950513773571945520046608677100728612946543287190247161715159086299084557321793893938960584780368038407686634759553025936214008738611;
R[85]<=2560'd115546722739980474480329526132034807767160513150230760675695873007655051003325618910933535755320573574808379199379205032476999760926628059568277259571367927111757030014547292597294403259844586270847469326425300201400705052749329389101448446685853052612289783682089883639085086693813359716856365435355865648476312220880385844814775316821921128361409133133715126993320295642174301284851899695322679369632878291308452973354735448889115613884686904486279076429002027047458404692923316591844756621262174199540105500490264214513197336055614267812850171478743918822353537744577935447445833964110674590255751396197682986065236183756911453331615499336143181385332893707120153338387201667854469442813254529648540896785191266641125265208224278123980690035854537379058964365155971891;
R[86]<=2560'd115546722739980474480329526132034807767160513149935515132330253078634144980767869227522358556578761931483629438364557992920428504703971514878329640098936662197950288386386274955592069048049273126550595002912966996357685427544594431174848824049307127812078132197943135190335117955744973445939684014325680224682524603729763910472553639593359721390992480090438591615525260137754746361222007753170442248828528809133153621330024590212658336673249600541434531915655226077732205105635104810127927062329504875269617024218897683507474309997132380708231484771652947598801436392065017148481810600789017495980082699719177607018524744618867903517693653347731895594945438330271014861119800475692111153341096066910381113246604797197599456370251588522279984810689491348072000807496790835;
R[87]<=2560'd115546722733675126551975260100779040857778286802925929017572693996570925743012100892605849023547579316137181328429805206196121622105114828930292245291825525670842756428588895395621555674998289243305562824111801723012267170638613101915242428081528206282033422420116238960957830084757744880409654481563112318619068813498732108528237176182309669204476995215562436824158086875403236793702077412113898445326663268714764978794696499354390151965993264959044113791114988843575537440168675724220135520895298534872190657503493263850015581789518028448565856653437338274967229617683120556477007123071938432830126786583600363458832859516139960925008461372050122324342741232868878571329770958917450504036039734074910551667663301252548211013993067755865164721540222615944310897452987188;
R[88]<=2560'd115440936454945755581025183767796949002830262420274793728727853277328389909550471150102206324641010733420777309765417460757409479490560898787542382425964333052708911020347818354476630821911748612858782900190431809197250968683684198116805232445815776550931959671876209574141889775058271223768189111415335031434192706587925744932080121165943329462272860789889248806925685151270379665007037411490885357710013918497730733558513737938189517808493233160637800178501561366023193245251635478447923306159205930143444216653823834592702118151355256294979996613169756356266868069439177793016034046551588984137978271858425653070603823584214887931476828501204001630077753279468061098549998587914649162436681830052816964340606788438078739867700879988858607149844747169232748154285404979;
R[89]<=2560'd115546722739980474480329526132034807767160513149935519657299989321451544994279597442268315107011040432114759163771117794431124489707665092447732062328527125201011613521112007826368151318497042586954290815243422170630238120627428772259813048106444047674346164856050517890202126637330912956113488879538877091017933686156295651532484127143001348190715859477562748929220789193597015718357345931450694025060028758026248525313056602947289929125368950221277294938334392667680172923651481464810399917905648143484709011272122177543216050729053394850400421722709254071207849786473148263989228641620332467989080141636229125671316526669268709938463888083262083875246546216602367880580705678386058854493582993059614876328250196566473086790400857591860232652428419031183881145983120179;
R[90]<=2560'd115546722739980474480329526132034807767160514440199223063284829015232741743109381207115084245551490284461812829567083701948735255751623475903397324184796480187870748060309191323041765990221273236431646333906331843522337427904502597932970465014777386190628997154568610625978044862922875810648331172252588098602743510958379540967382055852629352487853166734967639121151870379775444749392554580833697697506431710091087310977158295527540397035920016417094506118747683535694565229978270594275734915551244526933373322157708231022087620721092635107506564907267135248059128926736562869983304583177732092985661834871736314911944896200516204080771410422063063137473788703492508252649637997851900095020450949796744322793793002089024244429433860699958526611220971260250011675264234291;
R[91]<=2560'd115546722739980474480329526132034807767160514445239315654714457295286574527582045795892392864981951282730967140309813909046289827255895982900747809421731016027386149839509354720351918455185670917861421388132121888838549041608085821626902064957801802130823403945266942305912448000954522956883824750345368646967129000436782207312187438805818010834205939174981362961792608852384700921999034232487571366721617168349525152081356015409887359477377939817917387960309664599037141410649456145894489271809351338085735281284087755118964563712082851089244117621916399570329598527010900415254902503255359441222908482064770352695031610908675284676177607171939597701901737449814023232751491446537614092973807625971623137078729037798357658680706082266804704297327367814270136684189528883;
R[92]<=2560'd115546722739980474480329526132034807767245073167305730277168628939812777834341317908057330522244299882100426894246954842433841755145637102101493941265907443765132621802504921296933804411247709529457209601730452476685002518090004936694693392228961031985759940704310865126460089856228762423727657649161077444908032672705242830059754554745052622732164453746947866126676387889710881459320066063183880108907494494407207492607453574835819701515546910908150877504360297428389496226887656980216571623806365976897361291705762681463384272658246682093601393113018552300155626127969731917461040913614770763784732859735409766636446068997260511728150610741895539411280825610460290257701122721879625485980542354453594276408595071930693178549484807520278809188281621207486165844633006900;
R[93]<=2560'd115546722739980474480329526132034807767165488482988723828040602644177878707693484547905581960321561829035076913330861309311369049240888737382203644851613525439239719332939034491975061053919746871998295306058132029258734070987497583836898914790808036360260254111312783358359373543886992682387782884339631473703748711559190143966510822175591603046301187003820293148580378532717725240728014649023098404103212417626119061263240633334079252660040393904666417774639424084006231748526588776381448808785402580764457212886754740208638419487403411683451392915081222972124535175246424520087309352933710456627001401756078853216665610684094629546253086997226834708827820820574253142978491185080697459488419982355199182112185578408550263801897359485604392797732564146987060861421695796;
R[94]<=2560'd115546722739980474480329526132034807767165818714598930853925161917235940977577173828490825478336596308664980578025390538837458796619209210749880825397011756114698910025979427872652791322008026506615675365875474273838763268146487472399171437927733859127588540496177539696923013354481748669126550641792411157459982730050865922983419896009498736568391909092659888102359226242469240298150433500616505606381146782673138844409449812204636357870083131673312597010216485956848779597624066257864452545883515685718674634315020874746311357270343408333396281253013563399579407550158755442832820629996771208156625769524367552254885729865788742513186962617938692839068234493483415785404393633101509922207175378876172709207017045204065674036423764283687746289842678320871176243346879284;
R[95]<=2560'd117239301686366907235464229640909611626777714585478885543984861841796100246526608587217789612380334697553239369725203069856406381647719925662112771961636012172549148947159257664692164890253599176622894888860767555413302883560725032384361458778814404321837428349247357439202141795166457138770999223154625405421310383462381198336146095537633024805827776284995976400334526400327715021987520154734151282401399434336579970620485543147316382260886186593181759072585709669146078737491143661985022991755785885661185717026485694108320571112540780853484065956280036896914936215457846779717050873561307849301547042833770897345287095967257815599727763994344555939640984154177929210186235897196418539620561430376407911060752580008087025436561583876161629545643492758281012542609503028;
R[96]<=2560'd115546722847145219605422843945967965334700497923310313381834172213292348366676753675077193410919697237697319405030479499143190657336878576568652339479800263231699733112198588583222529886736190744365176005975037684549316444622228801826092979977822912375269938720602573337913796858325867771309552249622639694765823940175219233013237181051884935358447198210422939012560603952953494476597964654955720118971760591409547486226653769984377492762268803146564411445125814724377676296314291546299106910381324310383918070920645222730221670011407957932069615652811861464825685287546657088741630515058470863213178448670858286752050736644514237640620688557905106936205195628555881942404319727479611446704126293660330515986210133454246611367396246825760991639581246160808901309230236467;
R[97]<=2560'd115546722739980474480329526132034807767160514364597834191840421667136677749563116878101643028990179226678281562086452586772609081356127322283193205296512809460151686158533332603986639936933669864568694234736822102810734228436226497852019349863049119496698375962585757869847199960558736117659995416338875230404764004978622417673350567124568454539381217555313745488912293411967216318156341592445044453886154851888323052826223293116233024446347115952578619638938037837349231077276349520101614219967145967763383576537263327517094592325833108380556140613414292326744953125237997065288066329577628846451349415060365495025251695542006532805235132063810564981033948755792658518295286713354695263672724008171034954924544338248354935106994437035024784058619668936215922855721059396;
R[98]<=2560'd115546722739980474480329526132034808093144645759505492607490535018219430356551449109780508415740113423485433368994495714470197997021355231629738858816017695786336462462627049574252664440500090710228158620003843579000229285046831243712902588615073162973938683745291183014504810548079294215481006072450211740804414130088095265028151995627082496574646383688364914842742363509446309576024534363452211057678368024614025840874779373644362177358745808580846995838706545344762272274427536056426598045914262327489291464807577700603159277487805894756600923041374805814656587748281666372701486596679234360878235491590403257036592144389447667103960042458807053978490220748488967895908924465209292127754029123186180229495206894092371003145050567647000008431127093061537577429997139012;
R[99]<=2560'd115546722739980474480329526132034808113597908414647371037991602900170213060117717930659335852179630532720298908904228234955007769298288550225240062224798463240731230418350483721950572565486904127748026986411020204376389154691030269433630448361038050655795032326293762812075205963493256871380311975130971851264663330368667658108395379179067652770846373717560015444393871664494400692991768656796525503500372063298405627611194144461344839830094035983680431523848583091744118077121234585008527396758799329498473226646030928353015018022739884875034557149622863754798637053068215262729017541344315586281559865891951052951654636243824460347309433736831948216112501261426700496736055972156617044292321891612896660660472300093713216310082471545232304728681992743650553511159219268;
R[100]<=2560'd115546722739980474480329526132034808113518323735055451393328835276927933484029269430565592786566020881936931725556268515992638496069618319878554690150868293213505296050671526628971800473999297645304959455240914839592511726069422654622378836566116880838666667410744014125324752769609852132552173999766124254911468560320609955001918632099749589279719642391572155903057397418487943241348763166633223533847423113283411335994489873745701388734477003793057788873532626183270312409129395686187435933096315933092265147549392157072460038588659165643430752376195686068450659237792126653983989227141147082207200402783530527842675998328880379117726270642863342482886555323311254447851360477930688389470153658693014840967581318647020287279951226493406555299090648606392622340200744003;
R[101]<=2560'd115546722739980474480329526132034807767165798075123292914807376962944107273801102489161780434352513432695057102991757746280351936769700359561645778029460679146830904741630354040346739904212986319031305680079464176356604911885059613132774733708741981582782925306875367589030823541539685215919123567355378859047481337767801842903040059913533013424987728803712275460328574768439713712722212014626056000338978015444712983691675004456323737275800069165043188957724305077421690313079465441564143643952067740588580376257925222523446184426213861414156317352787277966740136040210135632130854523430636413038275132777642057389641433495930585786287270112445624696064193458025287356080351268479041888471264945309550283954653082034176194215303877969458895249669500111601537050837533747;
R[102]<=2560'd115553334376489796483187516179077580145977358918222934262383407884859609485225263792852240876112240920704280388042523197174281245397166680213252864758774101980053138314881243186871233999346968714510291013416445057975436946686220642867762329159483979478719352815894660506630894530251618572733278343479246746842391291602989608996940577633905578311554873278753380416590414500914368205270062015239714363685819025340442688879785541438098203329878896705418411800777791341626840990597898642910170249919710493781656181324515484033395186375292740088986879627875333699151463459442550282910794854482315746135381585254661797587448837467696291665371677703923152999694673238023197933194145970508504677370772956977900976269400137861327149816565748488230161323197215149194472760526783556;
R[103]<=2560'd142627985882163398186656758819230554505193553130597976292014405741628603189146361726649053336938818653889077460289028236613734069736128282393932313794882913581432694977713523266023117019903757414210492099311678389766379381878741578394747346720723489450393191728056943847287773047377225170807890165207654139316413149015096673876767457504367785126338247716011669929186848894692322839718716775207457746566433104086281646623787906607298396355116719185961432801377588532878423018004790381315134701419109963269610829174930873573477807821309659287937631602701624546120063292549708302073423548912729250181164747637776067540542500899585310571544742576316064722280638708128427871537366137995915159025584694855760738618433370344658537422145018461869863640289196525023115449708332100;
R[104]<=2560'd115546722739980474480329526137868337807856828698470564803914481822959209989099126455590824417461061084271124328819486685696289722649030605633838544944257380633693445765830322164648973159608113501774725188012904249471331866779907772889292009828916059602161886248683782806488690256209589825693346063756855405763294498121717244776347993838976497502896306535540734515980339413384049839674571430454790444831967013022244292985688970213149647194759012103758583892484217204814147034367507273506017774131880767840533402610219908601710751622750204740873558047512531770835298117793014253174812883319349262197704340280627345223047375492350231195221258120382727416391101634070435612951734265140104488586162426890281796150145452654874449402140451547497452414971360175967520410468365107;
R[105]<=2560'd115546722739980474480329526132034813330532845668383172466323087411333054036379020434573307127829556973479434202240916469833906844901959562319486953251423896520576263968828042304015631493693401299381282475468950855878081535503036601357435736529858837930243690116739608096653876161577494833276739809490658611452180281130119400951198522562897853147313263993759619191201307736053102234834586214190395254674696499432576675320914972108809311057074906951835242558436393958819018874827323281416705783727679305580769958771820196592972251354533377274573256857619271176370846271863092359277838957270711452894271603895564137597863778388269593262852046046597257330416079299716120365991497694509469295375569521407423621287491156874358199014899211307018296788996458104594521370925478707;
R[106]<=2560'd115546722740006740349232757680016847769738627611122503933025322306276372413742789929425240083119925240553915601508495477545885420455802972341514810398782503823827536010459404797888559189534530206377469165730855268229950762476514875401729115137043964870486418710940137457963932947039069598427325489494762861737243507239496063841261882085202244116786779090189659880480455025832687869727138084670907765283559793893241499791255699765186123488122744890251264933060167171973873051631242953802979115223106512162596923364324311838717958687845114524513100661961612130046757923143774987084783516159898827840025844033223147441116775311278362977876070681130470582305283125207645788183974033234103172033139298887708540458424238760129960776337524369260246110674553608377959362898117699;
R[107]<=2560'd115546722739980474503818801404957826031202979563998549025184451467707579560696365782925605850506030826066347251824046713250646357839070017150623149715639699314939074456869761125855121191054444771694311591878632090626694802949809147994985635141119154405262911328541875641340039415870146127724086439733761741344344015921609600740568495541137693803706732498063013630977145794333008921925347538563316172855030931363927883901939628677179318893381386711952993298832735140868771363119170363270149310238422614856903511107918362245720667826977581105941691673165592964031367032216859726345736000776911965556422417583085113025606231572980491718901753654788340617200152691896887839690203327922188082107684978312358973519472358093591878602576829080464703869587331916554854339609576515;
R[108]<=2560'd115546722739980474503818777690934605362589700973338545925379247235396649416366876356707467572339371732264572444695429562748785855677053249377146927192772339727168669802815210531545318800654814227760345531220570931810054320498795622182941091176130214633816061005461155340389813793640139447350849543917079482330023808536807892915169788554718133646413600597972297272111791295420708355216570301469083634551048772170230671462254120104346079806021806805540497377170434382333818919542303067165101998476448337012803129136064583855904057582141605185287283943885695823177353904740579630507414355862212773044663408839997191041831707980923141865203743472670844627670996453859801916814269108438244806743752301762140766189821569956422307014050641856126680042747274057182417718713992259;
R[109]<=2560'd115546722739980474481797604354146930079881579160674152826335009961085825269435585371156013299819629550745441151111574592091367994879127497841689070576949143756427359865234249833291129279608277791772353833120322632455784246290983012926954122645945255851106875749883759631918177433369920841621925330688306304293718512187904397017113812880899461725921945379309080807721650405876131038761087893466261886371367480752667322655116042459103438596336928989776097960167162235616172749553058629291759007892705073927958315108772007705076529323513437964301072740584567235404038616637354539190664028931850152902085187229870273576877935141227617346140433605003787369140901232709603272770137674894275207554304595062577097663509449826235263751221462695565175044776615756337018956059722820;
R[110]<=2560'd142627985882165039805023042501880860498663422396791064203303160961961237334925993027784854852020654107635563599517490556537056245470469757695565892295171032528694219830518449703495305710995488047001231376780997525423666159134093932205262270536278019186910200201358296347279876039725731597052355172993434579670316161804333367368469945293128478609437339333566535106330833382189772332767084808178836576813246767250462087791508274707165072267043589991155740002917993666401976712670686975174677454921526802259888555418580784714662560996295888008312831068116843028216121647545468099637297097171459678959142105781396915803084956695645087383555644083304748953246158890474247721477910203264519129798819325898242037314827616752924085939911817125383059953413246664785712980701758532;
R[111]<=2560'd144426351019398421528450960115815473095211824883102038721252844377195040244912767434228808197389984824031856138632205351113601123726760202701809861994276133256926904490761163258235699001389548692706181722390945932993872766122921975633259555243425378820369820214427999317710142284037256501816504090232305156513408599961799718064968211539632834813638332281385554203676732829354061889875513179749519202298207023755019014537032779310663335631412943598024626683663507336631269907825331457405847535943826282072425730245254741772505836147613111483629037516189168960729932866689035976507664709202372928995602616260439744104791883325020203775647284595765132412622291239067606979641425750950542799364664151396830203415187297946204652270745349305792423568390745562662108671460525124;
R[112]<=2560'd115547163408162660961671202962855970685888308194562997654957562857589580848392093389316305235179687079134673333747495553632852951316531057826236725804773602375925958783905513945318245528559119067492323822857844185866119024965962256464156417280436733792474111343116316737697874178979206636567186092896259810998801030123362420465008308925498808831375119471974487797564465471091159783184344197315922595619117775345546311889505842110799274828848056540388393731242110245117751459003089903722354427496090918691645042324997254816661359786750448876346657926017636621284299350399817318837281083001236228266962463684475101661868904650870372512457605802802039258646273654964555574270521511065638111186727718706935512493575353971317030138812885064787436724199763725368913163916166195;
R[113]<=2560'd142627985882583754715213709887980850299487595130662115957630676454773297757872314649669352784309323842652991594838770209083652497251975745928287637886041014388125902339444242980023905800902594914309610952257087252465941041549288325585936804562459051572697467787539569471807292375271805769406398010118437620608961792509179170691828974690080577295085183793539218423087282079112203690106160122067814448460404662986932460295260102220549400221137393882062972213558599205254724575740043381025487542094077699426935799128778994932667967994831213229028568488275056623372339754149682203699646877313487242257870026604068053795452412788352641411433497599526655176318090257409878258591395729579029078176647154132829240508708678432110407424439314792948895195655142335166549113648202803;
R[114]<=2560'd115547163515327508312084770870077767016175722486494715799242805608997934874789241906798501978873595107764903875265879627774712914498118907954710239141742967195759431951433380057746832065597150058606032328167372435065845040905335516669342309267561862875626480528553161986798411524571676152838753920077830561956986810718429409311359276142883394140796454915859846046835073004337923464653858911666914803783495653759882917018731598429852552360543978040164125120563768577057009644655197348323425617349193740415307615856402164309469677176148505504638459045305571809142733493910424537468690521951081184302543778386954006512117590910025467391551030392565464991892716235158543330114712816649616823923907275565920757197677178400039115587735522372991380363426960499581545556608304195;
R[115]<=2560'd115553773437202448079301937109562422021819285224365559214495344754319147242996323967421518810375279384165408128453566129576583905947756148553911122547101545215247032955942976435823211250122552878229604866677636430629226751948282505270209588933112066683776718055439663884621807033409027064434783381094675930863828260914502952030788694331386711229020506039684609437577669222791728183123791776696166477144741060044546078700516088291560344848145603952421018728609615818269354093592305934570917674338622023537163402101473787135291529619670087683375417818332853162904482016468184576731042268069501199500220996781394214607918316373744672741102686907515628305479239862108788470182022218256890700373995790030854074464460033490642635289067182162432067682522597011411046927939421252;
R[116]<=2560'd144432962655934009423799258761913481817087189460724551378169454916430329537415369938127330238956957535350054307954980192057309892802731161955170556762950303702440532470395414545385425733340262308740911675156593772867188976114154799963050812401190843870983142402082506241235852259016627164486972770654369739574108960403215433402435546002207107680901664853480623888706199059773928451645671087857344532323815002005823024782270280262196728459027264314687290174999563258525269289819841557251949922141122025738919376762719433338006853006143854949530934096147259229133317768274103024610381091337490790876309292025904848206599960123847263332398992919826654558155436054372349557922982936118716555467191398902204488077551725795884305706872709317740960438116743624724114758183433028;
R[117]<=2560'd144320566550330171887573788464096764348446084982487975461142231043860008477668209640517901033783224896215823175735024825203746309506762992910959329783208661193628377684840512884834775869080416918001116301121929384235931063936934436709109991102355578204520519196079080944397638275360905565677218296086907733781904676493588815118124105254853979971309494881867286266921872417836019010880714299772647792901488222411242065798534031071188430043624831012435504428583460357469582880594068734362727126981765127564645203358986194189254435475305062857808651865854108132181457726094482149588471224432519747036729983006196227357509404296338235408752058442867331627000001741275959243672448967988776841706953578721080274077837766314879020699339704946165363758759868289827265897694511940;
R[118]<=2560'd115546750389351496842343024257687691038032807933014068924189325874721798118881536711082970256269851292054875374669135099546986132371005441041000846997623547888109046908988222569563185506400188399603945182812414258254050502302435657186962139433121135871317363318433504224395459460138724983879529055825491729686481134347915229964338182940514199403858089786277894105447256104524931565521374229666759489243792659707265031379398973904395011493294980318086117417716762571241574924283416408797787305964737019003876335460725575477206419874172918235277462993890783542840687650374104803224981527001067838173447578058333787357190235821492635148903923204358741060630657520570610259596955244078830016252189938603012728200566973957809277840540065716911372852214436886438656675368158276;
R[119]<=2560'd117352112741032918342650650545995890768122785768016538242282075172831471825469853540029827770640749868314166860716503918947175950551356297247218947690401441502860704171911465527624569589756278717513067807909833894782660849819437527880657349663197549727269335450697026596243233909429977792769896683511201110456885594594651878870253735081794871362729885929251421578120725499623244118291627543686927010041671467628096821195013081485484070946518245905349362749931797975737488226366286932697601513528547527281668719834214845027348705061368502038691188327184886045889946881477567304339625179655753329390984483730447785886277550428422353580269877218526170555340290003297536354081615294124130693873992327260957840850254296699080185451817326186441051504284349069927980166823560259;
R[120]<=2560'd144433403424975593100411907670875793206613286745847207965469888486340017206903177304158802770180597777086439110617160652345325937397807810600879104217621834972237478022690170630635019403501214652729094039533148478815802634131054761653198088880579233998826893722955771921520194097917714942703994155631218714391245493714426849352770897039413246579610823114356742703706851683651345874657585013467569159355055198278645371982859379683738810496742715524507667109200697066232592311672727966113136400641458338646995567474109860019141688418391869535550107733811148204635208560085986903976810969487815518482807044334629641984606211999857372869231576375997067640261694667434119862902914116922016905635991335615980200108612851326100087541224588241608659364331777250261604075600888900;
R[121]<=2560'd144432990298579327328901539793029225692417966800785526481295308750655903962650331855163168258449713116461076791358351573270824964479733829227653119996296989328107861458660424004503723513990404812871768661106928966802404444599628871604619381382509873359245133774336744165712573952013719280852164902150863731761419446575471760007837303221115587484693452386542253974457619661472943937576264501683408107703472185756004188233935858487172822102457831663436200779651847599810285783319932965286706434506931449440372293982484900273150658708170117933580055858516697459558393789822434722865031925625801877430841810549815732245664705565515577142810039951240978311475088412381035390571749719050660601724725106181030691585837308138360659883421914140971627735933598885808966410025845828;
R[122]<=2560'd144432964370988645936159619356819974937219550194858673509712004001447739665203201877991273019824126940310230754353483621907419182223891344657938782537711202570200420316445911806614605580803747208860591330144182729190186020039962032080327277695370134459453769295530637709772144518801768694064712137380895443482830746544043596047122956348329347267582821397297526173727893720468636601392465831889774797653892016332963067508102969162336499771175765834549720860244637878571584106726475116381473564018069376685322941250083180976435776120454677715493699042008138291927223667018011647265236318596259444678487001335949481055620114493845847747826015825333960190412646240780594661114323577597905621850031196078755508638019005786677661848785201448043276155609969186379542469655413828;
R[123]<=2560'd117352140282792669394085057289883430192559164799873108059697277707069248098626386198284940603799589147717747969332831042952857154440066642877873883900315968046193892227581435133936926462506736509442608424109085231690743010902568470275505793689203601051869087983161871525897077118232609952894485696969761777683520957575375091782587748663258673500605409588538888369112965339624506767919382280703594437032759171265083893484803153601768335997354164589545662045147454650799029547216323920290096670210656605924274127722154722685837459125411202856194212097300459059122282568842609683427297102701524830465705319713687608988393188251750390025555920076559699469729464973031243953857514210989057405789280314581229011533344894787564054232628591340167733845041182401631226425652823108;
R[124]<=2560'd144440015162370482357821379137659872103308310178443096184179827050930344109832846411377644850715563513736104363725432091571951481950528198149488562188233061471448518455722062153002724607077362072787374113916186730098438077450534505717875721905391983547903021256267116078812620554305958636410759339919709644178803655979833802873649147083783957542954645907724956647686892486052862104673970734598718710247834679439977544689316803021936317312778977961071582979722979172007698034357510915167111685788643365119840550092616558684601035866667210205084030210545605554682157319442452667578142202907876683221654065268573227692454432947856347704583295083037765651303241070245493369238226247729218823471253615861648636862995583568439563522812864793366628176745780649278434846643077956;
R[125]<=2560'd144433403525861166368205648961246794457169662129145636369355824071333312582072962332293219772761129412143383689544274757387352224000743030621791042762745210895570289547837329567835683965561243584486081727476828853738725423645963983392400008133878148935898197745328262891844338820265100010770853653507733656384413382605820219823537063832066572370246512697848640758769240626068230281527506830678739804518389698403192495717276290596554133211746166268950377909780439216927860236456111447308993778251286019079637830443200029750987780031991697056352182115130310087988469602540712608788000686057322588188062590155625701170307600808864501397007634900273407936685531745764868315393620642027373046362454263933069140051456024015158562532649342401860757740498719385992063710207951940;
R[126]<=2560'd171514666567158619432746897090015394949033252295904903369592862264929260578404221342165231271002741113197575773992929122405448041799060480443137379486015580276953419137778670956043851483129279366830972253431327859961544091838239532708096912420501403382071316625578281436446861468378686312964587458776097283424091712271333171732253831674357724150696835683424225251781106331076078637958398263985161317536590283814344947074736234100231005365304279761630697164013636173664611295339205163285640309183707715558815600119439687315539899273779059337807719516016610367302125518085506057582294886001694819611036765515212506825857762827472073297561008393364731624902676948050279074646940141106919165120926790214605318337967034947853147505235357614336572577027640986191506231320134724;
R[127]<=2560'd144433844099857314380267517075455944653953086777659327679519731529536515784270592549678741747183104720193382297907466899756203714947211108239033326360635634495234154401730217190115620161571912814543191873795532007726360658018887288726832445405555043354865285401603772093272390416080908892087650137102845312146628817657117528112737210544717667455895191450712707647290987756824948298983819221880076014723478587734936660930493872199997139870583157302516290715831512634374313612938899705431127525343091242047332620281284109072673629775238678438522868100682380785854588244369792078076911169072722916026233690542446010537886104224512986510146400399903346121484478923166813745221049545923277679493064352979912223071434797579870382283349917519521298660957991987657309300893959235;
R[128]<=2560'd173313059245760836192514000568621645237377902137489959777603858787953704555580786030255366373236039873552761904031949847124769680795920703237986340241073742596729746878036093207182763619102270655723582540412514370273363633263696003504330198101374882428403801824058938661386545038530800437143177746478239372739508541936152139116602575751371305174383780998475008875325956370843619917713878940172073680824107864733436704001840406076216956596704768241160537422728676880055628772921841564866571182062750947781714100712681784254053444020627513561654949078662062705611028029280826553718668743342875543100345615113999784513108774328964750780155038763227961112112994897355022280393104670994794283933634828105970760295132671261931049941156630909633219222015062062546160588842878020;
R[129]<=2560'd144440455736366636383125507215130285375329975355420905829923206290564959666151378932832396690383499103533859367318477180987375981939103059629437424527305090509231126009181687396351619413105865339407716711999208515820234284539032049617283930648887764873666158021143491173465488386602541108026077674878162624699951634482706335069665904874113907017777148579278102556764967457430548960245948364681649444386447884315542710850477870404188751321036642417525673584755441683472825252976508637238546801502683879856804537909196093243159941064788551124105925555237213105707665778836152105801223589313473430569487220872621423255591521307990987000163272532837588196957725055257653182212934900046882061940195681328026715230795050714651172984190752103689731098289455094770171387199112260;
R[130]<=2560'd173320084109970711720396799628981192934865035181757460987426158999377762725415753269057733753966743606982627063860151752543688009952234547648777942188891156743126990810830316002267676063423292384712090282897995031066728954361463065552404717944690456596853868817529051030173227063852942143099614979886345431520937095536143418920228015925095033769731697677465208663844534782685360763564445136844096822719838966541596116662653377340455138813434278154261582260216094655941595504543640187124930797253718979458550671256830021177176509802509011351023177524555883206660336244627418072161504159720467985600158251555826617913820247836023145321206018690454158809913312783667540743679892487841037728770816157924443627068001616690746235404905010577659248356329260879617983396079486020;
R[131]<=2560'd173320084109970711720494289198074994008153202260196325996383984686929621552508441955920515081812264465494085139967473131977906674132816907423851132346526042865427651591517571432043495695444506344847031033755116208399056781092165396374938082521403502995187687195133901463739816894763325125742643387672956901595406958128283997107512325861457903652394499508431896518238418955842407154572797271302946896547458732931479479562188180640440446027137870021558681091459482310034634408694221805935564877918049787856275742559932373576251611665215065085653664621840114149169937800508438942046689339846760119558564524087656180854584845157398318539131272601717151505126779670370880693440419259191401365367582491856828186135737510802453917393676623775059822652813515368057138072384717892;
R[132]<=2560'd173320084210856278574162545698167181107678864578412910053064726122052634834212296742538362384380440399396159168830900225613286200587859364199966888635088474614252110075556414558500770178398844870624250758796976288384657953765912664137383997137627837944325177812225368645524902528535042942123499953330226027316998622455400716097202403762934353187614945121580316592466746113863345511547025847140033402135466963589653298159988293448786206897583282229588008421238334004890352867775972994515826364595698567410668505184935165932489420554080779223890001889860704659207601923093209339354539349319568968884849619678957545196899663428423175576954679737558681095697227988064407765544498443166283386570248063179624115557611164707972701130695242552991770013871236874949290991190033476;
R[133]<=2560'd175125060984600617528270236199030682600872391078375281485491272839826093838626379473351642696343189420832235796534899981755137158486092679855825505578155810093650166547750066102932448756027423602461812577312684687368799896699903243788676204725283770990190747619868586359166060970595018726652020313582330664791067097820281015094526227867214906555704421664521494817613495847883232542220460445393373924668879194709910755652522819462991981790643895470010359668245640205177777322280183131521867790481363609055442579970237144934465434726026877785564621957671955771620171622764286402692422239356725453528513130353005986065193822503302822080137713789851496363509135946893235708040400333452493029307329110493185456678849769595614950853216985557430125174587976323360481983326340164;
R[134]<=2560'd175125501646475916688205496515813718363103045239186188284837111473773051751615462976974803588759400839522845650604313900865608879355796223582157169363901651953382004474023928015726943208358027840905489906008551728723731010675430563277281936749081635993046535564230472453460877997089489946730777737463013379306013288558647580550396410521764855094826930426560667327931327371678116626567286435772350827244903664510215482723590880850408655229812547546765897074251079501816747583762251443554572113422950333376104435275156377432084207430196949631055160793631677548576892427012380988675140327903129604476121001519301097893427755493402713713798619158523832328191551081083928269961388082332313772595009199524831089025672362818769518594605093290551435569919464503277175909831164996;
R[135]<=2560'd200401348967628628467732716463362203381269480250126773304218003278717400219152949260187768950452622300445165653164173028297777373925584879619204263558944835818646274112751909109620128551783507304069118965804451261723037152233890514538051263442539357575560954997308615248170028991677038830240842461451892753047477766794914789859206178913459160772098794995396658037673203446165641839039647136820794043935318773149969182735448203332442951484278424232704130951716250838162400195151202915400797304851176681083576030853622945326432741384464387128321913121623003198809266496346033726448936672079654461471136036669232242746201876922547758024740258815937898371334835750466689496128203733899606602499934148841965821174528620575268244736264085284612634868178886078135031777647150148;
R[136]<=2560'd200401374800218740820735295750230321733491766827305383932756715930686879948739587004942294816933040229547478833862965257738274929750864440853402684339600441588726133607357560241755629613854758249087267624673065566208840920161771278668707372845699733001720265203127709547612724205147924632306633545192187731451020084330882042284944239494732766606567521779115208533903743662466449079683575062025173707605741115817163741524922716626114019950295959858765557000376683727062452029860847830138472086892068419389233522856680259373065815451972386418592703715571203603701769623970677480664157060928420142333173497652070367919646408310570339961049128637593694896166725811210241531071571535568992899309263337417418751097000325188424944826687203306420093346972224164792954970309936196;
R[137]<=2560'd200514185747693830755262938299350315023706051820550619960365347801903497843993803698964817235690506007116942222623321767775921016185372206256860630520789958912912819920678746408511472084632206274997623235933265084223302447227695472801506286437949930676653810863869030773151756177736468907007244291784598999421005766832597191732827728852277739632209590180774085820214985038048095383576906927034244649516769715693465401331489453503417143263177518831799124766176219845471181145734518638339507595159215754859120874701701025557785037691825609325264907169257207898599835950088082469223912603806244650083244683742724824770648029448605638123699514775534833943364764202334314805454433114256073729419527325900247070914428758983138037504500424471077926321871539509703941229390349380;
R[138]<=2560'd173327136421361755003213623428672576960316163580955603374763197805823053999638242235390528160185084092225507335742207804626926390378668556127359110297022796064359361656617703737138794868679893620086666147172847816712873919479002267768025771599623492832730318995938505331567223022438608933889927319257200283878852279668863272021234349015093871502087508632178445908795565552747224399261272204465971430131443060561277895799565252879796905480551794997922574485589786284426195319193445766446298654640405714742653971137516971480635355265883474554411680173566464445567737896996730230474953328492106162380964180287147586775287585277632003675720670800702075972455902403851139010075628684041130184839996216842977918436844866884647973616124436588218572319993822484750400147589186628;
R[139]<=2560'd200408399664430245586692629395904247967357521980014679215149076614360461753894817144574797788884818028862250024356695769153854422924963947358490739454760106863659586451196687767684693926217939310557361093320806412369541241898765510962074404004868498171406673753005077617310014125162485019839733053363881225165041352751363848836286444428757772206867496901710312689619222393111961197500927113505764017540448714227360033343320197976225691978727232415613027206095545770868485896879902858895440479342215779833600773789789830711983553318170252745687627163528271383844440842820399057410332134951994178096320366167635044348858526437164247809254197277816539453188472547779879957561263867855237646804044953043639586700208467959247642808962322205805563734297833310887123504028992580;
R[140]<=2560'd200407986437148412938024753557508022563329563090833857872293383066573107631720508534235589789434306514966549530130698090826208561959107561339924996903009172048663654082928908866522060951637251101399620597593176112602590199413662126636870887071309514180443291489529562568362723171639625334320244786052769384801578545273241542500847905801213521227376230828117955421615782613083977516530485885019163603861669098168420993369682174309895600480178932106744150786777019123604316614396013122331958060569741314834215381913923835996919381023038288625291848780684310817897543185915057440392243299871844969118461489891443383063638680577366596214618223360825488708930418610006517269991553564840728063953134814627731202357685467724102437137043976145719393458515124187873199617409827908;
R[141]<=2560'd200513772621297564985220673926882606130787714869097518489467990658559594524837042090883479272265846730969959293501114540906331786891367699745359180632746959834660504628099401171465047824038548313480497676526883266487024749508467769130725219292537673731759171171656844109811559929285690808083590844775480558333096203541602481737542620016695625378065140037965524413815532256575886297119918462320384308185798797687508472806178511344338618972080050565585175746522509518882404007712507379657858759827126588636786492700344465863705270788644252802187532713001217631263662200479826846603597055105466070510757824178601813394837819402336749419585810316462801755155466842893825174376476774902972047806573864328459516950746688683796498076318413045716933019611960464893093653969650756;
R[142]<=2560'd200513772614992217056866787319656556323108012397043977953644306317053524025283297912686666436075599250092585863580898595495340477595291267238617733271829939717252738811143937759949743653490183179399444153770788013571744262365499867190568185164352251322932177174997609909990088300750223745902239736121393158580728583062824549373113098288886198742209880143782156788754505220123882923940753925149326791435420178619803288680548499793202899250315677803586178242640582169398398469779500797590454540216001959416844569864815972040876473105263396875853599284484879542583678270123869070479809627100486783527691077173002819343449950926087400254527552384967354861951475798867383656658498657551363379574082621134528105786280087378130618568813670051391926121086716832019485074127078468;
R[143]<=2560'd200401348866742965777924976805630368212816704232532351581111940308100324443607345958213553709102361684172662023645703709531840440380783677550653289315108938864317550773436509514990433933070339882679101426571834910774718973606755705206251785900899705337068732209340673399955265723348322729224035411525843407202048195448154929240869224925213783098151879576936623397760431355417735973655547348421941958926898955701229283169889160009403073871409561980526396499356934363707377680110881888152971215910363403693298484754581525942030684667659981823458424021956560125892477325211714697654780560377262355481095179320691140593188408309640720105179327780294208048788519436185240997552730581681236914743745962582609460083492982444945478593913887821143426516255289902308607868491023428;
R[144]<=2560'd173320084210856381176778921363167702529155344943423763233718197188477904055661905342755545173968698556972540426378951911753253628117869030485938066424601732026816016809050692583113069767688989031506274378937889352913504877010316999588693447751075461550887023284695568445828305665696770246672277150982774430080013564511271723932568931743910093053239393583328470427737702487220991903947274497870504685202227827321988917371627812999226041288539609584902409631172203107405228898935335387770179286074941380580446182880798388430891999826008710239438156340879176592696405802027378463739383777812645216950030659495475745375361706782074706676587861461017237615499377117527512728731650880069215014874144568286642553645319297053606045018889941814852521036527932224723655264414483780;
R[145]<=2560'd173320084109970814346599893922435566018663704719245323402356641894366784551260783104026938733051462171952834227672510434147700452164322940883621700716720271933754137301588502233228893314279912574025947509791369695019825607904712167958147539038573028393723111455281475378552404000928774393953102417151493164337021933672837208145110587118009734258135824643295412363909512561203720164417019431080043954452998894547837911526029068588012740497650913540188836988895686065064844060744821867811710621116686704878082092735470112783170976108992524092166109250250694566149014290246760710570768230252268572746516219302582521501380827295480193054742568940924532634478335280752800008334832050524321857538066742164474922893189509753910762716731779204788960069981672628597346700481545284;
R[146]<=2560'd173320084109970718134625531075792733298815691460631983178726589883017839195417704471215361514408003163031713673989893860950654050558787187183932813080739985397622153175372512693265554405312223991233485752060794713537384851621658286083642461888397925135754578107751476591633022589096212746859477605388788587976885735327151271619197373163304795517745797047382971550059727788504768337325204314569785859630230229961302993771557315749643435218294094381649990566300347362645114545971768545985449969434600018495251504272592753531725568432711204942570912448376407664583280784876410472184215418464201770327835081570053836780249102568838664942590019022590282533296349496167889463546841129255547207985687491885672143203956877243108060789100481382398044702204908294990991552059556932;
R[147]<=2560'd173214296311652490041129546007544938388449306845407150614215942535672371340160117128629715526315991726191476550100993344951558696135326629301181651448180620358020427138703390599775593814766070353975095507963043156998866737630118756881538912309696379314780227781530911939470934537001469984748943778876028832801824046074483651517105514097463270116988536455226513114028282303170394773385518065207654691282210020028168272647581411159950066601401604234774354132361107975537893115807872147585606282769174384306143142955314676154835106725371140791023966927487121843534624554212886983411256896957812175155718648380360042945634121588575802068415847512151334333907026284009336740123847098519247527333297899195608384116607627090268966403290681117097714554489094886130933354319856708;
R[148]<=2560'd173320084109970711722059880878247195429792390127949869287941238382666468414911119108615778059965539475184691547192761922490948515283210802569882700655128218655121432102787055499288065747074105866428903185923952399449619442041345462436761721090373821256015624433175101777080240318403865992325352138917674131507904968298817814668130718142972512301945920318941497052162865673936672011277503693195856239879732439805474069416689571379908132964670411962267010280113167082919602414337149430306901452086737605023350197715813730802823598392120473335168383982939942251539228415547225081973971275422335568579015954174213358510899680287007406237951418021727664693940100373010838385542913949017338263364307059641827668732262167231233399740649333027042451304130160902267050657158808644;
R[149]<=2560'd173320084109970813945808806104553961558041396985446303460286969156580404314533844458724650083954648390112433588120102726603268507039989017357139355735062443893343531625272278834520596440070118851959136391105181100541826556377098031022871060339774393203035815364295571269763851113300529208340154330544976422096475765221949467683204076994093989116949433203358536623735278984703004879833248500907497388558298605708785617497302137125411354737315076722809497175459303143950680821329837075124748468940726597710368961753945705893131959502785486953216209473728803431146240474374299069254400314864909678345184219237480071293968905806743333252454133996639158751339345686121930217570613603913559263106387425397466018387929731768574043146113291197008251110521534402519337704438907972;
R[150]<=2560'd173214270478642027548652531381583748392246053720238493498107370779531661049130598855672651135166585561294342651991855695674277913736894564336145047125214949449108934150023282637709923900490966041139893872965750386032392780297188436965206652149893055757687311599141620845560042392057487317381317143247283044082160311161979541697958883215073898799930061772051248228247204600357500740471722432107015890734688024962913646740658857109041940990610952748735295566031512775181280609754770685641749583047203647564774024963226946810573766908905054037215460083770113298009176609254054703642975786694265376611843593152637337428631642683389157484740764475833749549103450340591785470042372162772033938359539498591030056878774244941114210509030216016280500257069004907621304421794989124;
R[151]<=2560'd173213857251360188910225171821718191344796229765948923970508061133728845494493839774548343672079179986079993762654632804679473166337291453242751109618529718074219608551104973613763961839238913264654163618458162395190604945028680461484561150667077805973965308134854012289021501142331992559494016828087921591872606199497180745229884910696767826933565426500789247274897623791548781079377741414606927028170669467295163969409441941921306610777925589939366221998510955268362306005996367081499658752698290421260105400620078382246553718747762971110869110434835098103322705432234110456249840113152946253724658296518769539285800593722920687114700096513766604897542213119526360257999646824968637150129129867653971444689534594340783430928341937259166034194861227721232612948923663428;
R[152]<=2560'd173207247234906569607712495879843005206999977939594094751079159209325232996594703205596029005727169424953987745136601848311858713915234396677065739781817524673717571743324633948796059131315757360945894201791903144767807344725511558621784029050803965251450793098644348230940253834287504022383903830644736480215559263163552369104617449674875059430301281421851787221547438016804679014384841207425525887461824298273361208247409360614673769195958632073508362953607027769507974747490458171027339440829730458064660763883233055411140907068612214545636613519829142589619511681536797026991788179926503537760923207939712026238591992117667470858576111663691631451393235099007138495202307539481830223830336282338399185658391978657623183408796487937330106819998791542573048313566025028;
R[153]<=2560'd144433403431282577033207474102567045892699993648612780452111854615336952267106437801156732353709236607809358865141213817041379864531916934168891178896256159898208052939991267810752008986857885642063646778434900735633663314103517329428342808920972537560733769776532407790834196280060102573342699078369273566870383114233574452373432498000963737897413762452658687147272320712569482815710693667956816916921946892210164734892198165261940869459755359275673458756613806457660984877767075960724697974613225709201061332714387914470345841551050036862630112135866228757520170512340477209487692900781566017613498350813684262382525068787157810917529663047527462991531871154231050908864821879526223324936158849407394544289137365346332854258888316416860059963252140085226721346575488324;
R[154]<=2560'd144539189615456359342812370397341046218377527512121058613238904464320235322375943098637151481551602761338416560373245420339279184988381820797126528207983596754059569983102094660976868149540598287537085551768786902458032636907828938457600143056783901112180753250884822155050561821425191433897058218971443225072409768275791760548052731689722771343218808821881113133805482520399096134429783722238839481110202797201554889353975275379752217271858643563305417313116198686801495783102773170180482292219452279188693462397661012689210647109324898278205095420711532293990050358209839468441002893787995591603774529207082247370662775164480813982840905515503117217818532732166514562078931623405696663101052645857478673767145911615600994936104588222027788533087995823937242584340321621;
R[155]<=2560'd173313031698114361899135546682356408942311283906184218031978682263461418226310674853195281509253019889519534262096297795775228922681207924010369674700256053996558270413021029930535535577429640566479248414067786104990290294733752478855104389691658521179557364624363996953068648085954800518877377982036383789652189055792980804738046646898396229761941637858803394122809058346115581593631860581289585492621115211767063055576621497325950401598181448368808033063646044494057444113263771682241518545483718895529900102295043046050778730255817569477954761864323568637594661787986076281179414977738349720920386390770625474732150525502425828343349811873206952148341326943035349926572690286113722887600539342561576686890206880640236231166661271471078990328009681529431375209766933845;
R[156]<=2560'd173313033412773374774481449580121819229847374525074461276299045989538362139983133790238018926641115399312774960502459638902286673442662385703304281657952764929385492887203976548060644856089196050831258243451520585649946629942689756190957160661564022007875826471328350901456373395171966539476760364235465889845086992491599699743995524560051236460129878126858068020124407886866952964171291894317163775519438197569084597277713612910270380028992381181198225754565095010388743273422627820619291769725715638143023928795223017380336876291220802509558959632669899304232085238549460517949819100079329821624637184218312115409497512439325986318147110015111015997562777003645374296985037842829890808475516339946885134429622270893208760705828518025582481400835015775388617096243270997;
R[157]<=2560'd173313031697718731851017401598123323291987635240277169199855318346921654680171906267928562333667009149531924536700047755639106435216707043518132990770038319023609042475948952783986409390042758965044075156421233196539572516935646328443051025767993121698398631160818985094826275891084764427797328305106369634375993481551774918437776701409277168967890884673830514717492218297431896158707436123132933790137440872249100250150242426394382310266786863188407238987990326530498504373720259582921688411433667826759641255508275768561732060225915562180443945372163517228127567679901324713892071860664781733595595937886018400549446209020089566906720214317915355370462069175008672938798082665477020576951286202991235473872118479534704002086925299893795303054434380723490654768208368981;
R[158]<=2560'd144433403424975593100411907758039595422653194045011173311101083279919586568225187345136628646023252880863018426035411477691901501098598018069529481014820095735845612135527626248487460854535517217721039747945159246734908255049688382434319420476232852215546048995237740038899230324790781926864424811330006581072744172247429159429841437296925101608418878503488831945774959506596975783591763503019391409176139593557321454024020384072676648049551424212204157861302310623591960893920028539329179111187765523056089796227908349797967092305891915187218796255602148342377310216857979549998037188049128674502235996270368806443783338873811216883000994972706976479557555541504042757270610700608790692126644196659549012940020280244109150124591824814659603678976834783569896195795277141;
R[159]<=2560'd146125982370968044211074895202125743789474515880658610747565074959448935246242687794428600344488073909594642976063119646787933464495565945542002880974922190499465496340087389983318109857682075358259766840099701579637736419970986936066932488171465182193045986180789541500918595081910868869619124354688359035634542822742148918290241672884028333141990868620959894501810338283972883167687030018197142960826650721374505816962848632322709712422266383246127059903723315424767370811024221435458463836071569537471121913364510831043809005761131510899528630581333489760731011444741629050536487099974430897093185932190271968947084400907246865861549765419608157830979655753033026029617509952250047616476556361567654464264458153806992232543066792333460235336356557875831709686639711573;
R[160]<=2560'd173313031798579674850352455345015744002956392879401516759976890537605717820828697766572873424031227252724647526428765112065974818952915310937856017576767796039904582768369642129290118944835001334109112848688727856912320424535386746982192040446453308315540449673028147740108335994030766555341397582553659158147868997026926159623044105600043248868913853904783990081782548188049026837925420236128403326342361473459094522705493712744099952552702349368557069838437760606588875800595050940431968350649966284014448200466889175887875478240574568033102119781651484462760044079107709700506652314570406097047518636616666051055962604246727081455687035918560453193660976838116873142279245595080621927287682558241467958564450998691160633821578893311882811327200899680351179985363752277;
R[161]<=2560'd144546214472915906188216184447917083267697661374914236183806726765012903282706018956612086518966995107303719134065482828282725031352832013298405029756096106349485411232482599908596175618948964444752960326754658288097625936937715653490339693540524228678689558462070802763896790267995523945895340254850406958727910171837706633489454569955303434176397635234992528193960621379848900149440994961188318692318639934318797740209291987550226936397143813078432447810126667174882968672311017424707956492843578775411013528250259407150478744946022344874953822773699751200193921129674081333558236568295261400967509107834554252537698043135513370112051480377877458672904805123516779540718862270575862101205188873912140096676270128997073297149048441947926368577986478938816138341290169685;
R[162]<=2560'd144546214472915906188210449767406108712749415733807029176397498404465893902998279016454565788261122733269004106549394015469230269095197366971443567668501108595903952197662463938391751089441751733156170555749192084733231415116655948829101409494605503709983684189196662364583783636878618359421026894598322513809078505413493515761657061336601809476885471097236706410774928555179726417396792774063123980196393975455443659175426970896141925423108070099172779697944165780620789608322413879039275724577260995736469561543074916633238916647457631279837156838936718932390426446639203443039914407342606550580387009150619984087117844102590958568914739590746075248296794852674982928764831868478841212316778593724887475098932924874991263666782802360345767772194651540448710299009504597;
R[163]<=2560'd144433403425369677347402127601611979397705948792962051861017397849111114359466429641032757431107781046039574320161191557143067248607113169376988305386093989693202814488613243633248476872597978315209679885413676895558820851068004805940651286231397674509681589155188261541145663887477694211455326604031939493135485311334748805986554906424720212900482186635118395493023704359541703848240825016760456781884112654110109778767510312750612643687450527047203246995057622388133973435738779764369829049211565800258187614993048154856774349375926540861460929541205531771807785095480594288181004872215251988184184191555602780890030714630913679868755805011956396829285356438507525860846539493882324703763049415422673367179575108584526147727426709401312521655131196087764084567980725589;
R[164]<=2560'd171514666668464337562858743284225453170555658849799169398219949079883032495388804372092277886627564607958240351674115780730741725531988169153489695176591599802402478901635164087182020495216025592693801029525380817488162877438648659098922864539933351840285113560582187798839460263149891346972398383977406466344237346110397430311777943006282166811215862371112392707469783357164916479329204138732860125680021348519757459216595094109766358096847548980743093646638471227489874943917822476388655722681628235623275528208884800813208142205931978535703825688060924757062700640981716619865484923209572908666849117704071771236109585254094022346778405287626541821250831387636630986432005277846343396856625194584858489893982818815030156379143733650150333778394591909996058694311564629;
R[165]<=2560'd144433816652283697983570140008654153158987182761268512460212590145417612017325149494626871985292369731427016730550613411572617942221599084677548029020710547686349258719957385648518397636579459121727261725088042239587415159226911135944398191702095789838901185137871265435684324565789199738087464612620097947995891763401457293415090057411702772778427237011605341763485897527129790215173698469971973176222342364204809480459635274251562812911860170812164685480005463838801475995220260235232427971442419081650671460268361846501678592247101290402538009761650776902402028438754118073870496564674536480398973016480646708158165738183551593776146782622098312004796986270680427013675347919894898228243421864553973426816411168529657435912506211898285589793066222242981842188114416981;
R[166]<=2560'd144440428288766753741702632134906372114042709993845511007040384941832224154562950338833782783663071687159285604339854903227108300139027985994681930652072149493552890701269694410557360517822047461362693314749294563713513524576113690805468479318090681968809625713111939055128750239557637958879784048472349246840725438916407449885331287413994503893821890776975620299349391184396095695469836833140248766600974789470001406126787889121709365488395852118556715208095338174402793750453038111415747612369272613793148779509571973590182106104015981661802433601030982001650990256337083551398296968598562067523039423808163053734709801769462665912244287508660510683696321392813643429743863466035925065208129536452733683417625296744198724341445755102919529472691286106250112892449150293;
R[167]<=2560'd171515079794440349431917764818048133813697858416410792227615998636538846533899964659388560943859315356599964642081383188820108219977907345645881670169119903725773426490642976874107609155687036583462177356584767979502772363779388887524088024134226473187406691021516564582959565586608071715672519142733374433187843661727362072354985717765338162632654929693145389785649389425828590021202775831615131521062537323647897051869748174320984872823885731292685434345262384967375671025649726688152322670777454088331340690455479461883441034157325267659657931422513427456636068376339619879164821122216498849294790301106731181316272758777193938589183026099021073885959111337122158809908517821218068035146733463883171545810229673265502745757805506582637743734166662192126006303550428501;
R[168]<=2560'd146125982472247592685725616208086933110427240655618720147005366433949296225878942786743362448820075159665004009042066722909108591202641530017955391604595554629199691787929450743240415895265260234194793678104904484695959213416971936597950650683198629966879929250644499485404630565550869198906720330441288938331450002680116184478107779023840707473436530259825951493487050617842978070181313993770054807568521005992795763988077958218824653860051790870433647961030406939224701148198159711235860530316286276757563556623608257172035631846738088812890990763479299492439793882515566621183565370367788502567422259815216046005748103890565351673532837410369711981859243820712175810407196423895920198795149235161356024328711617713641413902420040021088490787896581190522365732088796484;
R[169]<=2560'd146232207609498125042037488862240454357760646990620652309270047383938709815642496771909542570575061543384691497706809424012309320223521682936240719828602433042205123965554570866202874051887106061184992032625229928245030403551235159576267554440120463230479300201231434971175643928415053949771110506136777199867315267623523608744815377699974098763560872201282752044169904354044987566043951448822963656568942840950978787841087967438976435558693957855509550706650711199914381761036410850304499816360039455930347477820190450692600299079598733257433784102497786823943549927395377847479957232792726359727926908506462968721336143970318375063293695472020637226168182924256213396879608592788321271520933698983027270507980017713070387645434576368678076264115415056088013359946224981;
R[170]<=2560'd144440428288766747728448522090027874021298136381128323939839399165382982315156219310310248927835195444329085511914178382806721415902712330469609974777285359147594895410320192342279918048345772311554721404942581009403974369809778152906826618565567067363740582580151048332433415162527232370421148975680408834897067318077633818379865650324577623375529444349927736140354061159001131266874159059413965223830873261961321677504970369217083510378053380643602912938837844165009501349161814445221395954533331125195363108626896603122384626942231682280083241324522231598390170785638040157104242105487004573770731002187236911052733547032248990440533976544812358610124495324928519009656751670962152183983460705121965492095466879154089553051848627559200193267586868476726706888064193877;
R[171]<=2560'd171515079800771867017201235478850071306248088221851286530788370807348448931987451848768641625154246661138144240485220747069912367324358912980900039243862276776784251278180189311889717778352614866199212647682143815134964017217583846502572737799176746152845122917827693948554393365218164844217150033801872478674669931397596449307386828212993498522279408714422341426170833465899900184703979414099684927446183359057494767469031015060695908752993158015267079871563347261681259960748162417429723987195687449386295399959519949414553514443561092808370972867316081391601725123284453562074408243752753805066312382561725727125930537315501251492622312733185381749794275941062564155558204838967924951770017397569941791338900943527250581932180759594239517358107876851903410989266457941;
R[172]<=2560'd171408880490226449199963026848659629679832341481993226099798801334938391680489620867737639959337982464787988686013060157841066211740882905428752205716912568589145210722299429621319635994128749111132152352670984469451829878623469037181543526705162374081193655093108650472308921599622612160959618428891049614634568343465734197098447751461590565290875795958463251272715115401783615158968521639732689895093715048297377788542071502078144786925750387952911972202641464670528084914584493974573975204638918115218055737964714624339226647491869779252308113313974094997222375731766155584548763712696904674622331297494966722764763676786541459990815561454161525314216775645051177480854948000783390048438799377894507417256385531374052922081367185149273700760232754431459731002239571268;
R[173]<=2560'd144433842579848107118332476368203441277481655266914415011360878649905144345951942799600684414707031128162322050403171081732655950882199741220656813095316865485763614510098700707564465880866341444552943999663290615004875136818362156025091805424774187782043208371474283382772809565100846852147114363124356572827822953647066834196247161635677536312332769978156576284484760551485931086120560484758402089411960346781671278039322012112417993395907910907678936785073414963096662031653243520261064676107129751545517361092699067858059457467614950270990005384965217534239611137973583916663773381053100155984310635707420678764410643341902727973397694801524216004650021000341648386183150049723704348808033372919786123900296356313543233005861076566691500450565461458189747337911686485;
R[174]<=2560'd146126421425348973372137693965814976745246505703256733426587419629217607338838258094809677575320983737987443286785934439581132037885518644815349674861906300129067236930302570410978307041665429312087438092482891515111543036624151870286070969862084676597561321644380336503350946524862174844359435231006645173492428084568513182391767617267636750824426140375899795824364331827251943990534642317093105222940004829027058888551495938399515170395628737698587113562283419586323088509363365982881664303204766991485176968612510620424951543629620194801417483098682639355117675685683498726619921480602879302663524469804584791258912018333479403847922738472298760593012100132485552296037071551788128940437619653636459412732889618336593081914157343945036634682748584740436913977583555925;
R[175]<=2560'd146231768561816532195215865223917002871826787930079209976062517995603291734377909320259610942822183987080034852429714141147170380383733267624660306228590314077297775413103962554315785198504177021309085508932003642948928344741417789981082126272264819270864050984872639494174826795226745392627045034950846260895307899815557049670368584140874069803722428943838700152528108971626310385988908839686803772295861541630297155411349640150122909501694558471266305543443960939787930128620509920345973287921329809604874505026643789906341213293914220375901968964941389864438945270108183234425637149221147606670377551033473223933275444100745300911651977908027082199483662518593631256157966481425123609494957094561047955958945243727058058340262662308781610570662813636215767698259662165;
R[176]<=2560'd144433405045450016700707033793565872396068793531616241346843684971733325307708074528770536662152971022363911794890850501935839505317449392751151118911742032698709272615679664317811985666573114681442189202633958913011886481575410824877920644998949103594767930217896226110928552268222415263273985819659948251070969065203134684918446926654972535081311578990807429617830622354036078106690923539550663098149484249429575588556256079960341870984515029864043271157516563772284994417646743790939665262153349309415654036281449398281949159923672552822040204135776997500691068133452879661166879345284680721295126303141358958068123369110620266135957277159757641937983373654560269682881017231863919917613181457169556438536518477590764964858639878377251897838103587955589121950608610373;
R[177]<=2560'd146125982377667380149488024564184584819922123072713163388101920628479957696382566711525467954726784393573788662415433291349903421840170395775338294053007692840677682654161315706713232112712834867424365669459094419580828482364025398422015978590144832658472774316492604929439075881354911716756201902911573409619692276710565009459738724236944210155214909089897232504503822526761499325209852483023935688509632625887984742842529858108933284631698249451747499653515265306873953178741386862728451150218739719192286523208818559790274811664040352085009248185029237154605910598033590622555051036335009758292425993070214882720821990216397235852121933636410221447714974912677157287950412197308562335526734392482734361760349819074948206743917943234862893085597397724097719194491376981;
R[178]<=2560'd173207245519850303880864343222191164668249746769240691338609948596228974501723249485853012113766969841076170270918061912041119914971084650978473700639037840358621053408372986434431368515506546303464482617031174262651603905806464341361611889981998716550199798254292015909271615384500866190862854800219477044914735912151614123021686769363944313151548096162647925538531812891307946593222017580536435332604742966579717814963288400357606614657229207490208206203701548988659092695439380442665273505907409852299413121198412964887410905172344632906999096644152156924942521699562303742023639629142932425893669599438209564515860028412126229900753836084679701421419093047426841636371097972859488848641668470249350504384730178797847216134295008992697200053880362745091094559518446933;
R[179]<=2560'd146126009913542133412048335301570305688323283698599916723338460615483885970148754233787057868486525380776504791298705723401218589902616103423086408394712218580686265279167462523777585370059276153178779874804988648652004739308051672917291590493347007461973511504731482903283454690872188101268177015501003603766135664302441105303106990224978165614782253300628155032045367168209338891982278160673374044344649596359674222677123646487928606546843977407284254345424657157326673146326718237860136133194630700879738026811565622861753228428203116996847576968247487946771000742018523439320420637781163739305545095586702672945636407063292361590278120236787871084331605708745202239687478257651025445703936329136626823164714400949238279592069769937349596362599568487292982848415679828;
R[180]<=2560'd144539630277701118497641091889174195954556622639243223635203991644831604716889961411955356687799885090883177863153357273632907967369113925470161494559630772216734204280645124692443513076553587830740752463667703841735998865832360962843038307468009860682888354393071971921467227717792020156001000735627411400085275514676478551020946735082488277416811363713845163716045549547988620582493751038697433915256914137633219367951982765703489320867765698117296807451088618744597999525355604638888545433390635489591109531047551684392371761468107697048438813334468397981631772641783459333217690325444884439304242466267334949000159663901163155998407479590305558791034520550936044634455302047239377537884218132348019481886609622809251793030549296453469586971332381274818365983053661525;
R[181]<=2560'd146238819246427803573446314478527505815181386211839304478886387738239865294643415080430412823799068335750800090102798109370240980523878111841365726357830095827953811541836261025638862155729072455648257425227278466305721369790477121015435820757173255155664375799521032125958926181479226927906041994397319282214822913253725569102024318163218768052247856476776403589657252077292288158087139626117269688440899959340043066897615301134400126875706216617667076947617767878056709510718894527003133714434001173462676906561445234188455928429135714031893740295656258199884520106791049640303207095446783120642052189035616037629465814471869638124261576616500671051189823162021505695965558604882093242950864939967908341773901133056338011131004082561638112128327625349708051270121903445;
R[182]<=2560'd144539217056724633800816733542831520082140599106411597678389114764591980554187172877656579903042914204319140747224267794776391478056229363822411357234659409290617814749727141968410905873696069216439042268793706164385562645819856308229577422946267721962942541008112238202303665381856824675217238241244809239316102681778017099801170702236119891366514899293347965144348922866106285298537276693534839853845155737528973406468371675766804325632056162698394636594432249289210742191641601413798230519176755738906195692503924931725126416724925284837563848489344362848028763590093794582498567726964441466772948137812282868843443134969045759740375756495734627029066586435898866881050971351622906826644677745311497095594307447287168809547168779624563042929108738068211786824887391300;
R[183]<=2560'd144433430973434782739853940050741776409004291208131793685619248817035350682958668546378141739796133524704857530909216945534931302659980697579837368463027634094528753101376496498421547472985909711380232049343171090267349789626883038902175637961709430198123327955358686170817403171709172435073530166377771033941267288876546126533473678494450256410441728513230244489253720364054884272766726463609060356742761290801925808561300063691626233660128467012160949559086943486543733302519803145570263779863063082453642338539168450554581105716570374035263773198194266902886346617091355286034193710460589760258597702129303100264310383100660015287859330735007847283801648527583165551887636558300090838753733436763820300490063263868290925934881439808282619294049328282023534014311519573;
R[184]<=2560'd144440428396378019015538744223857988127819829238411557027050780662998798293129690354306592017353065045010263282782594907718657232227350162187249611477650112598507211358538212226910289832111840997970680647318844563459805279963726271953142678257993950956786026659147098608667626947926220505063255017980250534259188002217760734948171226771933829917231784051566523048496247758313237561111532228872491010198328020954868552155496879713276508649673431918623956695574555476676968870625589004233906183663657078702233117858056123525963829263289122727834935189259323673861636674755572244392403236080417600542861616454884308364751381540996090443404779015937141201991740969195433954769584601037633828416975066256932829436235256242560115683504116145286825783886599938472137152206820693;
R[185]<=2560'd173320084109970711720494289198052122658515372603599642397637122773103141315620273432717243000144364019416400419618651223682556650883976464891746915247814524438646406020850361443954626222233086648376274847634417262639087498702508604992251451692423207296086971297530777340933661917043296398402193589008793277524752280407942280544505974194472900260482465284865781834148929429524479092932303019003349127568467838036174719864961552569899367787301514832176302681621471476224513842407376491767288926705437480951875645162043103187381255611132678083738221722595507353091668762524172757118170445140843436621049142186970520043597320708326400934755688614275525796524381863259888599088074161878165643403258887873967717484625999905631672795018023778223771763466692385812246474748417365;
R[186]<=2560'd173320084210856278574162545698144476659215983222750045244517858658223608634412594065705119391095953715537752061982471990827293916943276766978303014578323032402756400960304131087651002602389190991327330748116561746771216470609092070859598756482544691607908449131350366642487949933413723462722713683586222255412219265655139923659577952058013626889368779755695217789116677540282423011282354881423332016228329416039091412366129281564257185989699741590248281695287288679794114053233741849413210914829483972670494950023417461707323799876570602477616630963253068325498278851385874095414203030873771267485769660044011022565111107455262647891106725778629145772270239067656854349653739275607888543216773918390107935168164666300866638036725315233643958833720848059354537726630516053;
R[187]<=2560'd173320084210856278574162545697802668603473104194141576818797060828323519467341683979446571103357221299366829679977120362883560459545678717228310529993296221384673508952908330315156407903759902125721189245556657714128723227964884673571674262067918844123926925384359559945960405580730493848602143366806161494449517721841442061571521876416892410320255256237268784923178866937687736687752134768223964963133566072620045038194001722682403059766559476570050336582612745657756401969624981093716194144982595813598585756604917549161844851130171224245646700886372933020204698142375886945859060582395147098466974573839166908482217172641535910311827238994763037282231109480309163341100405999483297353629143116726772078306406658484303616752332256947305023065505062496647396800857462101;
R[188]<=2560'd173320084109970711720494289198052211650740769724901421685276251209038702342021925711395615016367082689950447673075385167280463643363111337012144158677146554699106612921750959259439230256088782095332729157391196905391257217807526622010709004588437296856857648171036523929692625785163057793868924578968517754970497990476174901885537259659305997942301617817261360358765232153192088594144676486067665103959594007136819177069430365352150310168168468980087149816202636372026358739343620276161744017679756946429957860959601136856386622415623877370564394624441436167429441908355887630288329980292013874866954832151580154352005146893799436485722771287281206755968278119688447847057046646316869382945713836211426791826419583361569888888478384059673754568418575752256987875457193301;
R[189]<=2560'd173320084109970711720494289198052211650740769724901421685276251209038702342021925711395615229026274340695297616382874058181544847273141146399452999920904365780999589056834644103884031514913375675976706381858999415059431906745875352628055033550305827676820688765416448889182272756215651910047251384328858633700394298108604739527752080484084903738718767205240592657930631886447366157580453594021415459423561755979176092936397289115177880305290217896150743027233839486954487452535275610813724464893988372012585461094969532723707144795896980108515074669060630998820688330346216532642367416247530739224916775078018446774072065359347197848635287677059025061776952193594718917707543593842310675676890661062696025874476837946843623476893090034698425021991874989787244364387669333;
R[190]<=2560'd173320524778126728543438681601089974555781345407454668744764204579998851484515655427933211469975501703259390263991567365084185945194273589957944376105138953954551706345634624431754152784111813277340589292299649453857766944042503157274718316710324260434430362043507849944081164519005822278207191498360466725905655046863301400032114721075223049271862843332205175147706575000050576009800942779249080761999769980234956278853676302417019911746878234538225439741807450577418820198454316325909089583523331857850845742994032266835743824061462698548003596649104347428373994576698285196699850981885054948254212874249651542871309367807695134907783578205538402210323895472216511092437716515747090189355249532164742813403138574958977332290672578216709084192881274747708850540280894805;
R[191]<=2560'd202199712281803653351994636397410003041686187264606973412797670864415967354259390041722998015697982118751680571256872140523573580233809908554606201832801812493427306734977520211844769251312482141824428936150955057582714009618253585845399365946914557888927495747554547383167260987337145497835628320604111358809564463310197983184007717048375808706364382837965324140197430778247059429205960078424985612688933514346092789324295067990434964590709515862589995736793641333943542423631813185606770512745874227200961785221438197333458925185456704081236118199300446816908465736871054448134519390769089172002390723974123641763541390022396432659881100599580330636686763542831935164713138270633561157065534239525371747198943599389472769182766156119548938845972725878575049383859279189;
R[192]<=2560'd202206324019198548596129204947117961654958725193827525886045919089470149186524003168970028367220667099761071851373270516466266998956841590430636641394501706626054533720889232109143420218102369197417127383681806267688013994437535042070019005420515400021271325759078024146934300336588350980096011699210098908546120105363063493513970137430226901524907090179815472561060744184988920112613053072268299288068650629552176901520292222827764687317838202266908329126341433628443510774328919524129704117989498933610281746417148332705477550035183556838037670266402233785830938014202416810016184540859815516683117332135065179128684931041532133352853564232110759737819892849465043888548293480010066172346880664776616749053767567464530168594609413949682501458921481235554086656390026309;
R[193]<=2560'd202206324019618898712022633942683804659179326937720548802019962733131372335114447527774197702305198972056617537734045765523109575841488552945818949289213609446124777930120612707055094950998667173052421757786641353691045857945519094280876190467846812939292185814190901967668846474487474554061468544926431625474758792426114943575903224133042110812648209114272722827189180381491509198930004363679706959928838683521719734767695221682154275432827054089902752270713737805800399220887294100799716066667721939803148757637298825109656813561273050614140592782881377711566912051278275579596140633548055085158867542229969159223436980375301169275227452885853838495608625889328791722163773592112277808047634880990721604720176679347459808717962935244198072008488739326430831658520630341;
R[194]<=2560'd200513746687007355205154146199977222683523948934375648381457558878148929343579751310998162874256400066981800789206283716580870357292668888944215526438733580333877794767937065270858123916367561480823192923616103924803084695113826985815295200982524755944500242342859314474986208551110625258060656808234688149963171246656068870513994376781182227755926486437070903915188789379148406268581210647808044299234564705130117110552140702014692278175921090391098624766402067063180813207233042996122544886414162934896273884282193815897015625022246040690653123650051408359624376663841683870255801082914901491743209425412958612469766675810605518934658776645913468293129923255042833709152723042398706685496523544039515477477943291183360153931760887188861384084853172008096442283506095173;
R[195]<=2560'd200513745072836740141635330736485021009477044527586253481070727969096995972172747917705737497162173397451845931195766532943262759903850999958790286134310497162347444905803915130664297535805000009189559578997346235336949374689955325885158969269135059040115226757255538726970099565512459937041381077403805950996991284209767608819880807939932557041452482819098687133863075226197786710240716960145919552705816761494318101628754110070449743642711684107592258844388661126820948275428006778200642957312215038212860557976296554441397798412579253788953014667181159029029345297960579844120715959031739805754900673636049471265403601721406982330047765674080896643930220613991195673132278701206180900066356628894424922552637461612920592543781162858952419062100174190933586217618723909;
R[196]<=2560'd200507133443028491929460579737938379130514333516995792728971986586778193367437087988753531183332204614620189336186891257068376760836661672048606335885043402119263768624071456723396663003738875128911587157180049530804294185765036571082835445831561558518732238709828089620565737801842280171586116684696325380991114860147609468212312007231522803218258880547875830643039888809484276333338115470788815062453026696328890622586352443988347634535279738224145821827958136730820627120126501449929886103128457382236267134670224994868852730594472224510921708585577608343773439571986677093345456360180459018669245306439747150132812563689943836082512710224807164148250586691155630161671799625686015962097790784724620376011379190604549599845802788866173458454353667163917984181182092357;
R[197]<=2560'd200513746693682253325665539934772887470333125319503828706026769696382692038672876101620391017743783129820488560079412378865822332748877874572229318936554713917303834792353583673395569895757050331577291412415098445688695635199238399270297959146713270132791186416790015873981021086851942377941874651547867380374807032011954840658943710630705013441427280809157227133951932158120089672412072398436227900894023097810195947839986265107613257751048608104823176089319843640552180854906938902900371432292895413723777780592863839557878822858778920163915568749669685106829150634482042812430799546075855902514725422824751625112654253321631288295831679656790066377006500823636238088528593801501427727610761611276809451709343189449479729696025317477222825899631728321170630875383419973;
R[198]<=2560'd202206351567289913469973394295239698174002001025897663857751342825274035278939060692284661951104096048452780342696197352183273173279059299321200793684146494077650555204786277394096374475722991394418361174377492468876893311768430134269860932290644063263864538054720449199433315316954698697801448908749723300550482101198748459291560492250755430873833671533130914100873554170121635399564530642335407045380302291689244203636368936927769558351041385930088098153667043956654295357360175408410721813167300664783761323121378726536799939080749488485426776958227818795261421830909553729927569317378149326876081750696702460173378469966277604929620138047974120266666148677974061894357028784251559144006750201536170061249900087711454312911823242203983534961020505174625111918813467972;
R[199]<=2560'd202206766409134900024323593984155077787398956223044937586523579378548076017441057629198146392722328158775493619911786936521159324583830722292327237275100344354223541764202920333753417506084737203281401276749054048523756556643558788467992369214308581875467289311046381292573273709699892791959884971796387183630485126306725216677596166910600082398218215511403385329529752221988453447773743567470043419435708147802698127474451003937501471347915229794940199396925064580300334550317178248085805518461171732248751336255941981666899753090639436006414953853972615135816369996450741256200706516592848274120456366753026104983838088060233126941805036825752209318888008700320803478373772866025606256503384043269068409112466703116574527757460929553242033856992523093237005936875623748;
R[200]<=2560'd202206766516719899451185915369384928085192955236374426104461190825603111457906252481680962573043139834343031118754856348171904419877820835648530357755086411815401668734489373727667452234845133751127224093092302721356876861959981820557955379217468977707632178017249952316442859261780119307019513008949217634579085638354834018495491523709880093786726374431184923621843173417799507965359491983242022866959720379067633723840511697778564399279967367972260643434048643269694473320333318763378191885096167185908487012751359654940102425132104633828634294883160853667396670775321080443136510022676857377326385856286495307117998030954291099004112181031380401398838037236870926168749897895616409578850169677017742426714152154667540691136314072655880513540220141538525340479371171156;
R[201]<=2560'd202206792343451285848921912356234226584986966910278940954443196802088781347327527615445456809617784341029367759907246260198780251338552441241176432092996549575688574191462916800594922833645224158012657657228166657033456667972596520800544603864405739405659892904940910375633832095227325177837797091457382260320765194621607778787155866745947322248552914486496674302521451257890840006273718078164207664217172300961731091496194250893501865037281545234084095635055634121326924230613288759233746516529385026630451395687605127768628064853555489081718646322801523880538526401298520347002170010961533471741273508561158089938497795161136924579850675050230995280530688547658961852101038642059751887499633207021666078651408800400055931488136461273700987001238385841366774381351880021;
R[202]<=2560'd202319603391417858767423717034479807361179269733937683751095823233507567241319699192973619204283765188629988545831419555714381916427970465888412316477806599720530974058890065756378230697864441002803797107833692735088999507986511888257119461575192074452377630818342520357239802474285801601259663001982112038484876577162664436110990413865847674812726490952056721384461846709570570973696175385652540105783425517812248313005350017315197694773329220280734410499818756711992976721073299809342478680744662156295093090526802684899658258484707408014899254652793100620784210054690102128327872123053872877690694905983168283497718472941308160231611533436756984572441244586581374932297677562055337561719535968622271652574962300459581074600341690305677877567326869724177499741694018645;
R[203]<=2560'd231093445480381203263993623621058979413425993388921870127831551738451259445594999804530123829691738687236964154332414322542438004518761865947288654448907492078731933079052217202600406810549136494010882833635165703182048063470919635556418051891640694508187581747609018891859027582276383783738673322596256567538222407346924391714254175467072885734684171652300133080376821977238409876387643708926138917717129106867726510173506423030546003049340138253598227964427809493508058750167264725910379139257173497821751058016573198903775370290278738933829428249295812098986013990371771151064406251452772440251562346952541398948572958551647788538919144499308139447429189188163507132770530041000857395545912271697025102085104456723202476464063118552606503809854347313588732233728218452;
R[204]<=2560'd231093445486685017814012193975899437600000830032229463762776901697425085144510391107474997392217010810952093779618601723346231566603429843521174326371251919858544664978056800025877897426363253023935338608417593916342371875392167481931458394638463340622099143904166485738268004605917568662911020393596008003864510608757743540691095056040917675312240118432768729643274119001309871741043753689148304907973502032597048660560339482853840478179459261473460382401185134131015725791139420401340895592666190387173415937317974761043610223319274359249413433807966339583014523137687953984269846426119473589582353066596072826443763220978780457677794168948292469553354987362522739218506320232115482040118630199374092764421233509127939594122337739604851365081569519811912247343693780309;
R[205]<=2560'd231093445486686653417570269276571480757192408376715153781166454000783438632986432318031193862789542269290164811071951724778772391116826738657837387514077695714632844604711265552829541280694487177255886690626805379867614605835239219709001952703459024749909854228017107275495272716917869674283367063362178420722511758771290676803661339474230997432431595367389372552710198778940755085322109960472216073611891434176580889783174226436781658230810465305826812939533838371281786240331452714842387127479358038352830698891189065059234486644346816720359055142059479198927676235214235428917464716993440962193970171861615298434639480817608034916975242261848481305749817808760695095407382190936573182478206769796843422869840177639726062653626961011912617140747355888349750994308257109;
R[206]<=2560'd231093447201741290305758653320445569939656741782839921620271365218409893227912346060334196738116389164500411640439184091006487581803059789740089478161466591771276377178028820096541302973204098599178786906364556018330502949117375831623232096836930486258714428826363030747477419229703497941929068776376473745423488848685402208628608679330065460543666470230733383045662225194102504775446922370130437783750994395821871902210690604887239493551875327790840221674252590751205271168621837697181172271539910883690380465393624016549075893154464490845375521812903667031693664596465063672883100916944772931439878975950751433056799378514244495751825597601568649618446930793157980150285226949612167578353051246038477485173904216632835184931154652196315339381503271111906479905151731029;
R[207]<=2560'd232898863022773144275199554247230590730503418352840988261825908378662432628237852946159413953120733378576291860877665010101019140907646676481296205818963101098204715019308656124003663530934036914220499007131459611276712815560359714756901375466787312680644452152961474367486455027516652241348898137180121691647089936199509817461023501703827351942386468494280752308269136041681849393167827107057979293795650313242562105099958238072537556392827008928510405349063038302264953678276693605162197754852740697338676320625422432191746868152981617236818123142363262204512216584549055089935768958565715365500448779477566220962435767654578787217378246375948736687809122602538157736712993470619378299307899490497689076575260285368581405276132362441223645228039933168292046092602004821;
R[208]<=2560'd259980126164956073971285910745319102858448164638239103743228011280356530852328700893664526856863315756677312570636786532780712504789148259307691276202814873997333701713021422996342863272162984962097988644846685646627386082152453067441837808121547378996757579450088973799508339849299395277783259359770085661775185482669715390140207869620458025933396162855251302485956184227096494423030048724803437079866673731696476751601023756261352962745897179676285919460904512766126755799591906059280906124677760924203195938031818685992334137958224787942821068409691266533831098516458308517809758598195523985310351483815250699421208243588009556736750601130013194214610104894557291850836297297435883065512767653592184699318616455255929909859612555612244254710443524302214843054381421909;
R[209]<=2560'd259980126164956067580741433797442918623563490787608399311008499870524785041137364878357473688936247053395408151968988989517889745979888136221371125897005172966288515940071934459576879097124891645019876079988264983043510889390860650400819752361127686704285741158478292292649631889271471830286492701581612548522021618813810198281404777991927921700870766615009660350577410642606773877943158360222236312300558586431287535512949920180635187953157388194793746508040883548979021618479719854089235606767522363545950312448978388081658255434267969760592473756949727157941480457372549613824745292473538259711781080341257599260862354344527277206753514005218887769018020833023467924016938339939791884711957230761278064959771271682435817851277695277014266470346939673688932556905731413;
R[210]<=2560'd259980126164956067580741814709045406016154843366523150713370052786860623909174897876281192176313342822908885306682336734262150941605961375304936591048108136019085937124686083266542687299888476663669102049843250843947859513112142477894246181428053715008771808408518660788716632386971292345877923701816958985534204105201327456881369827352236887587702283346530449915959022075378331699333739754752689643696322914610694812414649833004169803315832539072405024279792458033590157084621488770698211489335083875865318039608154839726104211285186726552490485484547179311114762524595851495816198690086323424476619878060038531339428547094123010909789010913204704035779520512435491945290367073355024561931740551903767450733613255529705103285668370232615590584928565239994350115216512341;
R[211]<=2560'd259980126164956067580741816103644878145956876960715041826243503432032175870694615538801825896705655102456217522980311475153206117430809467571139495401913890471530914339005246294744509261031856581234189950326926538420834287762515289177263221319435931676775473323566053232852396521714625967660819608160612913735463507838926117380871032453369500669876340907962139902881632259753224188532333516578875592367805830098716179537320236457535521273031070055406851128479968413919654831822767430196825227320688367707614726155014382032846596192194323695413437726605094931751206134019442326002705344835875497211348259219840031946263576925886244282893180541865978031376118466398936168455464115153461364255166751697806180492207024980730069098472492474752404299188817102754770769247819093;
R[212]<=2560'd259980126164956067604231067569569953397814060995491342011491160634224165084929923498678617974315052803978389820088964391307393229647295583424863463458128403079774820468606354392805178952717087165612371147980023979041654350425057971320900800170443122096743796054104685896900707677580122292812034742355159409018474488080698551284382148974547451621703249846252559565582427126049238954361364315133095291253209471704620522903174895605520141518491457649070957524611830929566321648844180093400564919201548258331786103758960976239701270116196216859330629293223621372359523405627929336227509012196261175316693690762665602984694098299389263377207261716232404183240473717726911161137283229917150231505866523200334021531967582676230495452386863913711162661813160991737179426852787541;
R[213]<=2560'd259980126164956067605698764973030098907314819011931001549072235361553803553833933244320640053151070090153917049522186591279188389892456615155667819092764207159179744594504622801667963870049709125620765362610568978993641531300440060704326800132014460277008487239217524217817530807289362338731506121791499567133109213941016870893951966573056931182211592628043930272789617581156654979336345551885524528155854268017401427077601392808589986486758914832918029567414589145557980297477918219731824310731845551870087654894428331307584519357957686420231465349331912864484512067027746885002691658054975327988877442351735317224866154641157443174672527642791841955654144248883138457668505789595594595460362217648870899691491922976666194656911639066685405801272096214870393190468707669;
R[214]<=2560'd259980126164955971368767429461309409077509466238789482946040296617717096008836424607579646979845865145343637015420384701174124411348331318392602433930369979188830895705590897952576676152618403197516775531492168954563134517997505052260401833965780820552543108573334715101117797263124078288976341920343584130065882167604024575492086822520602804518918920687299000338672227580839513280485597959157715565884644256348457679581545161886069590850155593926211905817679596048547387569862722875067950275731001479136140084752764058202181208243097313781252029249987951978229030425462557779545921706280265459126987768195146426111482729732772125276080288538531534727851178679819836367518121936495982422411791579615035292881030894610423144702940320690760196248251615293756171836430116454;
R[215]<=2560'd259980126164955971368773522559376525753434106105885465491424310522576070777690773967130273182672031049193662828488745265391280577870004555602801259157582532141237543895082964368889354747939188902604378733531212621005851105622573311843126047835285050852804799293794673499962118546509112488085046215535631435338166329544611576293130700419843642610408438307368294255337171958524341466619955412547292537821246300062995810607707463592280769161044200979707631132286102658085044350523082893343758170665183631687864252350753708476376391232171454029444250650125988427516869261987549443109505152575448300625448351588488960513463887096302213538539530472076150732248949127857864025969836344108298108246680310306215318209380377661891179595750374568317563452281317621793920137298339430;
R[216]<=2560'd259980126064070500327756284688296770443344765322255129896105215054077674446191986686434620803479214174811695819629113735079331175021438294768789313385701105536876021923954775322013385553980190261968164190404239662375285635644576319937761133196517968019542501089995257578629120044345991500159027012530884518413742622508561372889151046005753997120171787601750000244393008027912371380910086159498078655428649074517441309299493225778630478125031858736420924257948199345424458845169004557873501158334410821025076187573954077477867267992990691630265108878292109658436970079249345295973004198651573345138407083034431304908368441974036128119082983543936302495849130387653823953835891020161349590502388277929290281005382316147680026745829153158805648638790107452314373059693078118;
R[217]<=2560'd259980126164954431977183359996010877629421192244503329367372769764495806793162874606640499665065540474996085301961269426528065807620462978259196017914633807608546851118066112326600664798051300528833466263834599887572518117837387420032705600748461883822599604576809824218862243654548410942892422094778120903438423830532968157530915332819088622281438456538703956559416342855390223114036361349783879830938707681018474347897672177957002770347238935022813616681375245233934111447551911444225015545434770565002861921191401124335009039003211657414083312506049953527276084856173942318336397347374187848753932626387616462209596910532090375160615601772751053880195719654605526124743103640148595053006436104893004830394437953816911938830714430946905241054502586442810571469145527910;
R[218]<=2560'd260092964653770558452277774085750361431981691712236324700303810517494254196782366071859605259460739428365630057657772353657958753781511040553434627983647360372117274085621673367568406425030194296329018820293586616800862201872144488643497396808743121105066501508195995843937950353107280038550025895234030487994558241957856111462235429444636232612295508047469120145117678392949692441262487086142872092217142152345137589394585207782008201841564913529068767162797745945154761219130440230210673726564257171991092572468079465474728624920041361685054475656214045571581984256473784736134636615254211194551087460673284777978576549075856055205056878815477232828937639571916301355688370795983560341038702279275522618271314047342959678826556815352798235939753697446964928773005596246;
R[219]<=2560'd260092964760961473234392051505637168737056096965666500508934836268148935080672109974453136808369539213208988856366750408840732455753149342860490459305603026366604092153781270547308642109485615587577546609936689641036530673890881012999059129048210467216658085650006450843004825776578823948601779877651627722800265382622666507625438365234695449986127311254800262965192365087703829488807455922784721113190033479444116387824568838759818283352514158816570475595350042169372815745562999732822296550944878778013161759066440117049038690788902977922877979359150352323794924066431151490810034970738182971861739417576862513895777062884371037817268003808167807615585290028076069354857065420155885937073152403798318526194090131982356306865572381211137549728111270261572938922652489318;
R[220]<=2560'd288866806849951179811747416691804456111910891650210135222093941230013275430551075512040015027203316166889263745587429425862643610805056537274627360868283353248653102949154551608227993555987617114776977991638448842998626293354707238653871503284226902478435243539672903819457541539478522636882263761267500857251570457113190539796905848515743401515786301586907818752044785806040087061463504454170373849304659467424768102578455015596077864905977811548657173768743939869773435709445382621092004834399046484794780696043898099513186818689361893899067531520939793833965531355680582736989639441626291211950162361876241658181062395997719324473418862178152773849306226305178328095704794603507098002783788458893065006309086523733120721146402277639153556166873226234190000537247110502;
R[221]<=2560'd288866806849951186601609168560771520060194280524098096799299245751029776485362657104980773109842804323327502384825478792929119565744880778380060413023758057255008226607358271468892211564652477917475595758117213884792267785211847039885542496991055010042742697895121699254910786296136188213015963176130302883200761228612117900066221948855110602282623001514085454669436750361889071702860645658032129283923311477213703553783348371486082642509608564352192357962477008479705174344331553747132366603065339710935884131110819999245635683738556101819391720568918520249847899679683764285909107532757406208771794359359965897335263778701343113974219546499379001467809781342523037181201518069994676500701077510411884869634585822398701367361582935379375047756538356224584948918406042726;
R[222]<=2560'd288866806850345276860477198834781031691906707329246309259926668851178926335078966978000488631266765346253362653625733012222317850303541257672467204809011647705244129897571899624639556183562614815883219734292093863115539867913358174084152186545592821825084168019701430271118071600524624883189868989676058708644693076305308967644497145406595353646473119622025056367558246984614765409875188986721544606741333561916300130619345980596194861844856390357717452096022738340268333443560769552990713089617779270396245065971148580162783076290148831893330647441003172111863662817013543078100081903364068172332110657384654678914769442955275540066596947149744817170713506206296233977220085277077964266977318337262356323534064279197914864131796159226999013070327950479510488116624778326;
R[223]<=2560'd288866806850371548742629165476820992702587250880306442388068874052765453673619125515665958028427245181610143568505238536686391302359750906056337479631264508178347526656193499009964868239709803861560440693954919367017069056259283468087830608376349490592351372069567455305668290820402452945530084981774944308344367006208000208169906533576280779750662421708957320261611105305502480032366795544453203398776201610377403618830277132832605318375695221846973374193707769563624573567283977124102165533549379400699511707748970729353421997035594331581253824609453008219485765281006813790585589982498958481091982421764251406715879288215268417832382744361544560368680440116270474279985633017263167275466035505871890025094576281225985015374992654904566805038514067593738856525708227654;
R[224]<=2560'd288972593034520694775108629645955495889552051402080402061686394862356776562470063143253449167647901699458387384739900315611858247558314868538078722657212732160062564345104717418468474622266228593624662814947625209103336475338416909821021290985720562655380353081006436987198478173394231321178226176725773453519171359070107494122763113608763356595007230840293116522952390418317799955881158715364208730554696515336084934460332352249446343512468242758522915364939850190286561945958138676024275149064067760807829100637608147507050297838059103401744763432078485243216320767397242279612974044886479646249520267866740162944313270329049878351699338930764644896411836846234418456246680504856232224717354459522467015938071025364575678101980342569109809138558440903916168944928777511;
R[225]<=2560'd288866808571731527170095775243697348347479237754081687937993293280355524437938833138344238181879482641664365100050855828402115787135161435137230177253404716688368595367804727904898945838050769406667359075854528654198418697894123393291213699916853854958577453025160335544098116814604121485875657590333539150101447973399023975031603448630813498593399265221824055567007243490986722118436310074489657233368949880853022875344970212543455829736855269594307596007912999099903319646218498692609582641575029328791511227133572034819067444270004328802398805842808597377012503889949998906943822507026391782424099368002673701299981057168600783664367216967561651660572202122579593196689237179293157520376171385863303399868920668700777778294215877440109348064301087619247556768552015158;
R[226]<=2560'd317753461708241190682715757857929077792345210412485280142085232511938858113995079814748700851396477184445065885646317285275665206236621139928606289603745014436265581735255689383707325019340021025288083384129161239968896232728235119992076014633698922053399515294515993609515865915747875983005198472846596181811953529169001368198574672847671142827941537139296490832700353921402223713079352174335991623578988369074673285233738205628383525865588593982226805833746052957688234736197190187800229468400085971887179732821622648784962920942095904714513462212025573864267502345225874769307636705756996018869022888243685673479585943873791752841324188522739456689445926301933674128368923004565752814146588145019546101759182462033012437628218819748517606317006083878601434190535021876;
R[227]<=2560'd317753460094073762640830104428110437918814671191536033763068920764073510811271834649190867405410742973198387209777476264817598161610480729341899937345401536993621605276006289492648309794453613997106353699045008402342909593407683583067425754999321787414198242363244344541923241602058660585653467169272569003812685531098193644875076590433243872607455100958186040625538491868252174403629552556298911580098932232068356514545874128538981518521129373411407703083334821348706761816693942508027313344500505572761035544557045372175323312246814407841777081055767049952742469748764764761333484890008254086300365048412561488244625737091565951770236561406512275152953717732843591702841856053049588561517281949537343671303511072846233671602750956487833249323191057907152926467271644211;
R[228]<=2560'd317753485920803507445248902303416291608277572438086903782679358997949219473597823054048260535017432959417566769871018129864825108146614402582845626766841424045038507293247499070365118040169997139020850926327939299100022805044504062251485014452540618167778501428229925769623309842993915880125780696442787039102097163270416756034335620498399107196972351671628532770700856221300498860970239785690038002761339180361854541756842752828840339556063837440499229058191249423732880415873108112600173497444335715598448924767199102411600288337723334963005212827152800200791432317499130513672727295744688822014451183255065134428475226710031010508785759591943248035280054587645089523241361195098197032179479175636090000310887995620357858263366816336804785755250244550367538553640408116;
R[229]<=2560'd317760512398763731731977620729875566385882813267827127800869075824629602041568097705392795870452587379712346385105496464807320475974054211770590832137918922101662009914601694522276524368004702350004591898508001115290547974075574841709931007178000110806724869618867704651663951859549046996277294566269232037898888921946152228200507734520372687419590849791872076734552369478385796921260922435317503731889817044456382969642150774420859684379559689906760071324095369114024811058242379487874749273540946369725456409872307560000312927827107456159767959438863373275480394332242852008234512239098152505641041143277290222158563143905910500938020310749329901992593884593117788212266147891552088935566959778749138506065517071355227841016269597409512378421674818139507454278852105013;
R[230]<=2560'd317866326023787067975471229507657514056754706338078265587332643916376162997662236499336137929133595803314363541186493976207549592176863977963190959197098235580381014477577621617176920476074723797191919221359681094801250503164529476746583780416812838733533037436672603782897915864846470136974527444117725938706827521882514194464684027888752888464540300491764728898716691553481228445241123979947217841138590836424592817160452466721181577217685584255169755381789712632829698992349147758693304239404547204848899729855904484360613987352875142953442411362520275620964913696605042167345034710169252930068821680841337069133840212129350878470423186445721464645482808861199325827000453650622438409660557716300726942693738570767292910376994111822459751339072315514947366616955245620;
R[231]<=2560'd346640168219941423440988578401573441185677891353718414498080865611905406380636536481637617189009231841741977411133015367221425895156304635619182023321294562637043669680759209978464337098926956626999795712215428828167338954315955933909437895204994081424234401887111997329238149758784285770926145409544037258562911679829804700638097611862095441099458119993524589534487360636226130679761660743754292538190740136552503557342071617190795019456197270238568378928328444883980957107480173963775500325158058196391917365201321355157511711947574161390990643213096903331079263555572399016988920377305348012874374459881454112282369984072928654279369330723949769785189579952893478468163265083436150696125816475493747902248432633702998751314456638574392707447839374631787194658233607475;
R[232]<=2560'd346640168213636075512634312370317673931216494215503767680437561378859213983180955464045677203510228796939888441075445805794911053064076979210403796873104767911403411369908830534641595512731596310010120123547061817592294097220652806238556786640931325440663481316171181998336115682528183749304564848789650887727461541454542893336417596848332604350826870745034692644164974433911901949258172322500674218476564081791009525458905488759924918918593015245547287733786260348937605526963443656030489274128412299145770012158718909619696018581614500749253645764666215600872261340387642609188907804755912458421588889168146233994155178238974164532666234922148485349645904400791606821268435638703516751134355996932431257082506883222572889382513828137704710305405549002889646237305766691;
R[233]<=2560'd346640168219941423440988578401937953016199007389836268946267811580470554049938471859124309452907060889721301550656373323235022696392883544152659542516462690006060005898914736444592788379881482729021028080701829148763430476405175151246493154817150119769762244752301771563471069756380790362340784553214971661897130268165881832482283932933252527079830435507599887003008173366149049360540615918875990379376122564782206735259189951988025706090003957689611518263879983910870228369057168741531602085422613663192057101967977748588791076492177664709492002872213879564694436071521484720492164057532912601207819569571278959526566523415747112740764961831915368647286271163882498844679575486455191494404058127344396709801211770261524779020300738445898254624590980364228738262664255011;
R[234]<=2560'd346640168219941423440988578396127121882330137895166597395202979872110245050396659630518815617755026457006939835584069480493345207298704569277835815499910533442415138333137449552089878307507384189931987473347250509694640040991757603803327723395309019745177302692205150249949720473347859772471440644417535705400739136220121272286404767258130380439972887398174305225975068564247247892446886672447728886891104446624514890572173647426611827798894856493450530194701029170482292193850274110516675863864081445969648512322309910852178451082854122974644393908532691968190346229980513353679099842568500261592697464172501883267217568136738365906524584364074209471177360982317273000632388880214196513265138061598778379634284891526636433677131661697201452793269248920546999639523612979;
R[235]<=2560'd375414010308510779878961263126249810023043473222563632376277465812406393227934640416558362353085354780297539891240582719099080239180227344758327575341581286457632923469561611471706263574232923937689621864429163056814215836856630090076462973561840865153389880550660679530192550722235788911904888277988152190478699078040925751167259022279407749544042229153969327483280711197881875166195359647782900075379744978319863384897549887871351893826402277947884003358122305797535430976144643478325547820149572933309998172706206185174499928028294881707734854668347297209794270999506043136331059548776306649482026146714777751755916328722454283041344480254025094417336971702495407328652120630895088139081661434822165743675736505893926937574106501613767779403789763204065706497767905138;
R[236]<=2560'd346752979267881730114753033573771727013600836142968452719872259537860866669920231268764186648718907173091916032667176997217903813809589531799853860593145785372152384965171769829448106801681667896762274578730264012702940992372507925827314503207811043106155882763186411270683263636868931148644894929061118563710158335297111007162414828915403710328319006593151136968938907958072871020551033215438963826771476117755376706166864044408987540529975733183368968977642006401688214754619278239325135573631597126480090996016761913904208871498217208096943361230282395113210187619207790703132530572071500078284181077494739484797108510277717612484684130687393525175300590184361007752808147546805251707364723492535512445323620658142740234949077141100848129390747434655747885881414202243;
R[237]<=2560'd346752979267881736128001408850955581531484518720145318135658992372941514221398280997532052675476112220368474164723028240279658363697508544289384397690010260456353557771093499217486923814886482899099706000262718478882735792474759699681864840570292662855108920068952026950612790409731817636116274507548751322570993348837747157335266640676284072354053503501595039714557012239253269068051826152037210748222387720251174752947427642546441254246256464774740705153012565000210630309635234192935563377668192256266156401811410151964279870086118405173042826525039443187617790854534167037733914974019827908995465138211020852983859040257985324039402165376652594424871289308934182067462464167603020609511670824740602745120158149141587662838940054977729235000695685506749097438946350165;
R[238]<=2560'd346752979267881832339975413279699128866447205061029218773492225417117279689890679187763740326349500839323429788781214499368524300878386789659059002703924859691903322371999282129924105288102156819670871733326782952021120646337030686399130881816255110127220118072727759624565405948040214968520133488003868240302858425703558411612459027995512958505041467778494296056826116784682993099681081715981833231742947816957594618230154843727265593518838509545863227480037201434183443466203423058350356370880583124139251873186321192289724643024485656679988340749139195105582291084025559221969203144403388202371498823215305155700887836452093698785317292421373399005031010896810171455066390437394477070231994659969161428867415189767175497314924472125815496772430475080608497350951073333;
R[239]<=2560'd375526847183156297303773386756646517462077648882823798936402796929333504685096086611402442103545740025517529657294045910742877449674815286225510067995295685365271526936685739240918788500735468673703217310404066979512545494532240897920761917688920730212310835344370728052140902955851624680845659231844007848567702783109448519369181201082596149217669981121941422754927725289011694406196036420685385534048552319291590040055155592559565096177323095709747330027486440226326604628052163188706916573863079330057181757327594674053043160601916974022250024128758158359597088370829754079494944514210162407437985194245746702912283384434842260252608887877425635912592595352495036208206308580583109761459320757350618731805445042359952497987089606873966699837373049746309539590441248067;
R[240]<=2560'd375414012023591682260224832774341432186093865197398010940320241942362720154153961071935164833015641799541224985852731732429230911508687423077578251346881531034246359682208834407349408037865208405918173452377876448770064821394244962280501396365815375635687343343623737480358904048614727626737197096760116982439180324745796194409678730479313828286351880557855928476782161305357850972092347397041322595176417451452513901498929410614115783261055507607300786167271855648315358942085611510019656252972054019314920785928182806596973937684895917996797343109545177790245310315631945686183866341392599730455047000569002688667888469464748521148626439641488100220909542356887677661478832580647360044240181662088774571371473106406511172515988965889393897680821032911031325335647123301;
R[241]<=2560'd346640168327552592125462447271820826084773664378969846900844018080690669578394092945230041385578174169046201159586290676886551662658405419876056804979329405702440277444505891753482453000858821703842749495293245223080057521517685740424040761660015529428806807302058742924890391888359409814973059775733221887552150534045109221942978367736661677105225692966893696889986826782954381519261578132044158281893198059487283816001353585112469349349538776330570811233190633354334483718851052468962565563785511483866557108485320845254106388959447744467907521510622982111916904412978056648126796570529194373372978644249526835046044236947848761957594681743522729955925130844661481869568310852657933299078955993005997116812385578842241376526266395979015602226781898833569397353203718740;
R[242]<=2560'd346640168219941423440988578396104423301481540664168691521215530596532020320214926219256465504328123603277944993230241713827878014945816548538784772281203823008043340230355727922373748805171240271668878609145185129932532395609721553022300238814971960564679953466726135250832556613410515306744993891261978506951962239067605697661912867556342953553374938130734993786189468702873871815878768843425409621277733886857993397145328975810679952671763320195035950846007788349589188768982706267383307287990957130747610789382527601964618726349283264040762558814541005213849532079065579997703016303104140540545969322772083357833123020630902854911843843005892534375101167554306414507831103130093736370523788867819523405170131135796598508433482935271221936059406069539252101235402426710;
R[243]<=2560'd346640168219941423440988578396104423301481540740066556427449932931459321772011086682641403584071797330892669641883462085971192065260581406729869610551400716000463374945030304202391679881295816859551836664587354645135917971169901786736359708515092725250546028190817885553122566332115079741038386556453605262680486692097171004212428169589184212085038596758648222098033725196683094219079912971534376210725440168407031023881892996420870962409422906782467271186876768602622762785098344341085800664489040468491009442933372509279966240123066358087266500973374437426349942578362485871119206254324548050979953724019315947390538667360619566311426843819516911800739326334171382749577363823605403028088678740143054305192539950494576324350595462905114472873649337094989193213265655940;
R[244]<=2560'd346640168219941423440988578396104423301481539450099329056255358987018578857490501569753145881389538556823091392520756378598703362771203259048271938728907303361736039775599115424191606342345606260906801800653495800398467544714822363626343292677333271592288281379394204244566673821124270096571295241872063346207429129335743477395227629981672921642507750889869214776791718136942452759132200126416995955874565094280815503506425391712014604621508923732379226675227330252539409315248948537554222990771843939905259662920082863421083273609940366241217617522488887887540377908680591338215015498275953272610769438116140529853923686687763134059212023134448121571767176764172817728936993018346506910513062265406745632107803915252614103040533318796115206776420884010821662780923651430;
R[245]<=2560'd346640168219941423440988578396104423301481539450099329056255358991134014596825157887729950814840567191644553315481216764193635297293123177008761788330874507837511867348893734752859508526272974934544324407182116288839244844953223952011112299904206950660720857721317647779210306172770061492989086710527630760115125256852305868088599229289115457181608958853803330039208357475753149266487835078467746245912710533971629260823491208862367924706229349191061936369138921882032365175712960991305005753517205245632537499419072440980545818829063865337129752380977332620389037137282977330369901397677883197680031399236759846604571347609788851471174504648422530598435444038818380311980845182126984110037504056955840752868030989953771315012583662916625443710949360334223696976035726484;
R[246]<=2560'd346640168219941423440988578396104423301481539449802853021465380857286487650759585381960538616461536993778354108326053582830020695411279391354892743376928182121733169304164684145811969930785707329934532596925435500717735756284989395227554901626687571347057018973536335274985975446451186579738960490139171962817033845062096971095884402770898534598920577790373796751311797024990604716119118703339738899935516738149696791771844233130632750977144234982972164743579651776919616375432483589425957172719238219371063911418094967442000008583984846000687926549481953100871827430958612355598810956423000359937864370815240723219905685712957799968877711263951862807281429772588896707666512681014705196678032001409862197114292493943059719577725081893271450636608141294311714510731707271;
R[247]<=2560'd346640168219941423442548411501263510328487993179637824042434717669281223299693561269272373840162765092198665858539017124411282378308309600923934403297949077132998236916744908790519520833649470798322793075128151205710986185645114388608153922905874804250656040509929111008138475615707326093160542805901839428870177988140413475216918656803489845739762408829594818447614899794659847968450307411584169815163997569175980954774996827749297616708726694002762463221116263765987974104467495217794488998133054367462590381614488621082393260561784988648377487165971372020197099314097551516790761707893761025978909926536126733991690938029676739228681994540245964458906580566553245599827000284310722205169134384897348673383730893435952141280540128241241227521334430921393644306859140695;
R[248]<=2560'd346640168219941423816914449837511424493740794250367041995311433540574669379976050846637124737482801859805459060756792853555551204919278376715844022157024355508600600035415670149795419435383541576324152690860612624505255494501714010713915272221421576224024253511881988662597281592854658177985043837346852097249582380628548491155087884404580307479730233065584105050210448318382574061137596894221733378704446684616859433066916828255584369609623611355957869591579358597193580284436978358739601996487106669149345015433981014240457586451761892494960274560540061385566208385804499257942397557620703479004442260687929765254158229813213737834330793688590755198812500408834123034523488887140719236273395906551155552975298050356053971047395680551017725949718664474089842967433463384;
R[249]<=2560'd346640168219941423440988578396104423301481540744810172984089583077666636050469505723613701656642900787330967995585649928751640191056635342423168778031306540625089472260971810688563478533969047228680125817763231132322263518207713822077805562587441663777915422731486852853146967264561757173931595859084692202643957112894176464108834436900730473837761983499128684647481617107423073353886022286795168782318514851009682140238318103071834782163223288618785375759651513511786818627038045536930631371271256726007266249295869546858820753716842403375531783941599462872490319046333280892271952640276798872931671644970598473780663221849966141392541338759920838490692409370040646329331375528568438770005097148814539215395580426439717046226593354414466921835281566700958089593205974372;
R[250]<=2560'd317866326131372067003015893665959036601651860453773820427181990580597103168479708809591252460959792899450647022352480106934496344586445573979910728184975708004766906887654418499385757449478570231847337172390413813660959312875614541313811671587009149686819045210006618574526166517375515000114994153659888260795659117783855648883744355925594129739580635784245275891923675381903747265734203373228574132081370798749133138721175544910240311079122646402235943763350028607787175481551887923163558424374274786135100425529708114724117792472704553778950265515096769161298503243984277989551355792328565167091713011294640923562987012115357672427906755868329885690001519594716809072602770663560426390230403527671888696489041894887957320849177634735460230101816662409929488268714792324;
R[251]<=2560'd317753928310713592954430062866231906184860623517346588897287348537535536440914349190523847233279096277183259356242109249073790272779382659694526592491131195400723399521442498702458067228278218056755434271344232027773931501690098403664978130903152780840288242113186711826334962581860110272769137601590013791285605419486612824766678038963608902264228710861671961787491859432886624016917716029402988548026296637624289836821431004839499962327952895858049804058742722706031170188976284062120680806952701227331040442224439255292494962846309984295219320625661959483257283935041454195465232522549626210018962537424045065260507924418754852730294865858117494170506177828506246883176417141944848091532377715884618146108668121088720536892074693637637108916085750244692378261035103017;
R[252]<=2560'd317753928310713592954430062866231906184855649398974233554798150025926295222090958630954009424383911618501074202085463163259531510988125115545518276667966119024895609992638763689429635520988842017079502891361843179649883972404175177170418527358936384252446907254807746436633785953051836137622748526967826502922116800690290301404245081872838309149457517728091045972394892505217442809659997103345038647902031068102533274760353727975321318238265381744714134656521880564651408327733629107280122309477987618293906019011852302822380642919018697275260617645810520542787516375795756003457551223231327033315846061186113381469886758744836280957151564950240719974524942452725814233994672059938047126225359009056498753298318481606484561052732803001536071760848522957877495719411290933;
R[253]<=2560'd346640168219941423440988578396446236897591804476423072381459814943617731880785219567729902852851297666906412983414223674875956366531466564388402286067323730830457101613036638499421089399912468449519092639417597816451786750947870374558491033789687847456652031368860595090151799924516586387643164752653043483700253098216852089083734787440222260990608482582544859366084956160361017877615661476428671907292693528339371065065350714343987916879070921901970187195960366076691867597457396953589014281939255673533418726046211800829126164065329284284080934498773581119846982400717484136198913921411639027848222668052554535796108187029276766033407910425042215575341268691324886299179383230679663325222625255260720205213646496989383849053405821942040783735807293069263054871790327587;
R[254]<=2560'd346640168219941423440988578396104423301481539450099406263555797928604699085286685704155700183589463125443053799153322378797192554154423873363176294533308924109919565820666660490291489171502366077644978386332783662099048354769975383360286771000443511880431429263450511703027601284176831867197189718594785064788462608899094862091020870085353803578190242402317493420585889826532770931210368655729148934818785398875580520007253529838437975729197750443660618919150691282768572632580417586426151510071930683066943810540202700410416169372516173880450967306976329100083089241141453493760306847801637629920295757698111835369892334423794192937941231440095280891161529444733586500421709157199167834701740786364920259922358152881309899717669437768255557809525865663297408472270911572;
R[255]<=2560'd346640168119055856587320321896012152751365916607385772363691906503165932558255657593098072827561894805854769877973028264784505679840867025868497603920948253313631554116307334556192029329430152167700189592589369377879519736764341896177265585603977793525686678197913440086458778297084729974950749548471404303581467517097981555051722461303484242565959677118189631088800880084473024526957006213855488505570988943760135033845316549712060945863306523053489820372954468645052967497794337048001334423649132706798558945259949182444188690219834913464074151612519621857188954137698952500833308194398357458013167805090190645959561545590964839819194223831840061426939657600183981473776837300398542700302124625728390689115097789085227954247104919214113977686066687078928206229177570613;
R[256]<=2560'd319558905077758499734661345708908765231053294180287005130336638806846699821861687082859233781557305103315102975390802456067302611928537268778892050096585108684502255712305283503701507980342454362877601604714406773583421284263420220462824668067888499182649998612598625682620354414650651335605978913832224805451392992444103161974203141044778677661304552031020259452925633370411533367356450071726530979896246040513538997046847907632282846758900214733233590390275226706092534419896112191745167385978891157149596111723565045324479752893113525508108161851891558005125724480518023438851272445240747721048274435489173308654842500573460781770160476055677211361784863474418254246910781400444767596623524015050681301510998344064973574498504213411635863290582468226544466098569626195;
R[257]<=2560'd344834752398909569496505007151866130152092952942419983009574410394754862076591650713762946498655616471001756310864625577437103596013672230327700391901177496148444344947452554669933720019807752394050897296164834535832778862324892580784089488709053160083832129597516194538820318694146979807756042390097057464237415914211164420053444710946408438406467834762406734353008168971566729655404247621958646395694857970934217021971324626633101966331713039429818845950476959378852538032796377206787999845208001402972193835440673360699112590834974781513747550162783183657014164431312312691041397653584781341925959714413044460785113828817542467128736368608647556091590625836213651133461822326553156770539692958805900445656793676466283441778829740750093027744267999904398261273620787605;
R[258]<=2560'd346527331345296002627467734115542137695067288429925384942415688143313311164988261005874703863726665507281898541677338931008558265212530831439626710991673494520544808182507976493038577835743885483559650818140715973933873087538471276117260024327304569658693151953971029258882512786664211782439828201323532582214689552954392001164939315775254585790758464868554262623449817064234518404678373700674118095987095677130544565054642094631687310914694599259296033777477338381854642028942308206027515561828572154776715130875616169554079066038677482022095521444667022462790004872352799905555560203853245140207005123906407746780615940647694454392150275065056714359167158857636805701791896667648015813904375457874072037630405075672300131361284046861419372129039999341347959456631444259;
R[259]<=2560'd346639754992659590815809954018164250374242902493492066808991471967671609634816252704171384903121282769294268400385981088695138508622740234549717508487202569712794995349737797216897115252946002587178663525085458495919055931779792887320350706960886472469357557054457250565324128636786865263217091181637074704363883585131124816580814444580758470493247852625595835464420331470199360098882625163380040813066669102060279791831707795644997951422429637655327754857453576497276014680884560643819534394404664575657326793729288425330552329164237972909596712769459656129441610069562015072577160725859841802266529558095412767013551575771843575355161481752301009903646220811707132153856050489627274026527313326121780548181194669343935469268051147041051990212946303169908667685750202931;
R[260]<=2560'd346640168219941423440988578396468935456713452570953954374605331905678270040827841887686882805640261629055024316367123695012413901429867103507181483117186262712989058236037905425742481426553020372911639356188938600226845142865566690050800967240112514660669470918729945410790499817413537623241274882923091640535132957305379994359501949865607202979700119007270157474511503196088712725526686140353522445207348818950457825865195399282231283864545248607720830516300174179545859206332098937522350237382556380337594974905708352006894488267862905497326318467838482320233713991822305542846665582451298495648592716482748515382511758455349803731611200485416922599522224921564506091903163452662894187862827051234319560844155892431273562463216690964200356244300403455112227661369582354;
R[261]<=2560'd346640168219941525666210958102395002469637075059692229665610677603992878884479689264433871317288100800609409227400098169915240241945251583963998287606754324699441618742948380799998992012687556718825811032408979869046038569316185988505552094686904897759399519762211594454374614547470583573622629091719667421162933867801016384918921896027648937044694018037088809545483639020155070557745629568430462702052639150743654244648115517090239142289539574567767507809580978820941332938310875041362257210095942737780517022813762098951747949443200482374719693828854361416774630656632751375418631436616515861219180119859265493483339297626678785477921353796867014076815494936207211141190090927446792953295577855618991221594272840490037146439802521001445543909926906619651799674547381300;
R[262]<=2560'd346640168219941526042038981556833117873379239206184651105860292714730485270951161360754554777264516196773895614426308072460336810988995026797778461211508975947765576279917422673893601814298396719001333370438442490281568767448974825856902070072421065750172397640296778423154945519056963198360492191277470061054486174002430694906308252023247828674323333948617075311885472368171293441204265708184639369035607602933136883034497898792385735245339171146735671622779658462289783294811402032988408499437241139227717680949553225639549352540676380264880915740508076205472417250845440447078295878782936824075475263664786341386860612964210023633853197402004598676921158610310328298503414431542508035482457531514997563273990464401274871091607591915483689735632773632370582487013120838;
R[263]<=2560'd375519796492659931924689103878956955612449801074922459583807820680529429944065937547164371518790184775380914054370421262248059151490795606485150968366594585975344916122759695389410013611633961543057518962209404908495740981385895881159423471859940915249027175420390450896173020443414919670363849215956925161504530104308738987789450974885736189641960691372357128918100966606742236840033063543254521834593349313210996471279771882357356932463262451030768909193551902355126717097710251936931546740734173903045255950555498315492453560918869391968167425501614667741250151353100671465368273109194187499229206188585097096246287367021174413814027918726328662339483966471721925237504823274250207314710270442632675076217385310898904464441729325894306676842715495752866697181994256453;
R[264]<=2560'd346640168219941423440988578396469024470665468516135067705844012299696505762024921820213269354270056462395364231976543028095455260452211640910563704682439370937070337990551218780008943061288792276132708653222795563859161402852199316986751573259768854171922382688571835718750073249094294234115956944947837451695952537130786342492888952835910763455987228063862062113397145988846739697943215300976697228934044319652006765663066070493113828956296910529646867339775856097260739890108289860138494924311189876143123667370671243376914154555318810868925225101081367919123548228457656894576833380518366768516316835127034588763760690821379869659759462542579874911220789863567532414012921581170540546628279938886159758203244822796354602053938608139467286591613826570265123009207040359;
R[265]<=2560'd346640168219941423441086067965541467409853352444396337399752057404929482015340881470650229423754210114080212966469346530464279422347782588341819614535274894403426242816735944380758864370089342081589791651581018026874132367380616466111821286159425939109964753503871816416316501015097523718650393258997404784014210727659506103293249540170587020377278976579251379294510655969807018227797312043562388873280978675412106453095254665599354709825445710035080870844996289021128183134570740481837138177944152753536987636497677627610857389519708612697014993564196880717614687076435403989791780812961435093261964071194242499209651278837162448106766952396608169325360714874380117115708039447101981714268120956177265505340843094466518359298231916982777067718725853933787996220241237354;
R[266]<=2560'd346640168226640855616430936152042013991380831774920154475346350080875365168619692892029723151421497078485303936227836728583275720325975516689755591942993410380756555900912210105982597721594211298341622931841671621447561003202012662744375410682781715640834923492402341385225409524010824677242745485434968366410665445588436727953110007650508149017080357087270509969114599829527198608125416075042688289370756323284629654176805889016906370153688182317997161619702431685070343724967198003579887491563744402884223895344143490196411178962832329974496683939028132637227038548603539070385981833938440231869708540912726426077854139074815614662520927787846215053205525940759153314505223025505442510731292921859025604849561782081396257472423479074852861015146758034855277262719972453;
R[267]<=2560'd346640168219967695724023387837901322330270632059918143010196337897304302099973974769569402716286239118281391959513111909867811035177906249876146656078119099001605133430363849160849321463586576732881461655392928802294311250227921516246221927513037400522764080473502807225316407945945709504433244729046824027690698173574309481630184908664307375395762866103159632965803036373898066952691724832257901718753735581386439625025066406045929989813706305400739396120948199229243746073917322105775197437187316803003078186568772368334008877714378258640786813809147051242230003159166846032787113185601994659966501439638076133556315814831641026738014354505095846152901118229160205757509778099920413106894036888730690742032660380748623383679731791915025401320096265468966739965625668199;
R[268]<=2560'd317866326131373709020705569256071342791035737463972512754120581260180953104973912248487090412693658973698119485052389126730321915408114693447517541964137001876916986879100316895249544718831125774667537838928659843114593275346046541561270443015770559574229430607567049055285205816552018972058978197392324045676314710223938027720523508000218412316355348425626915866702767496997090061798412156111966829163820511080308321493531552024146807450640850014418133023102607900484661131489312684008119505572341377652342245424184847264851559240847911740976410349715125628764223047437730776400845520510432123185912253026011841024644493183169272346032391026262052074836214833024480616490929136234084130648508070001742036221215121456761954087348903343666655066123188099622204488056071480;
R[269]<=2560'd317866326131372169629121498390341055738567626568848569981339298389951892046496115004356882737688589055998903270657606190163513676637972636207188417938703645682483444834394364722585965776988060468320743899369830133506987074219835578249421631182462614616708266436014230465984609829624717937885000167921955336587567376628451032227460720024559105771843780165248685847936334463326157791382625726603931309946166145166227693627379257772410171912449268351556723628695626249120869493328870661625671963827984107433425468703993520529852233472311282272693679506875421850789874492649568568730883503527699593995230376446578526787404700523391134977636291082700123132904570453742502693992010677247706845959746446911210506224372810650782885709686574592630142142818430070621860730657215542;
R[270]<=2560'd346640168219941526067094183120486442460044670011671209123748445162772901709143233992884231559792232401213712773681156733321058968668291373374826935322591310617546755759528449269275972079191769536278729910773580764818623220764100492753879688106217933475392077176163908940988671669068407950577317279698458944214578591188069279120783225293551455851372445754976797059000878335845979464958373628854440447687068270106556536094455097962092496310592783076031534755830048116666211961069780850045061854595218190496903626135270896241214988790191835052127516458972768672940807975921207619765195300652816575837717068807309412178176700573345221184221703017274369348364618613008729308178904727731185604394090156527032181436101913417257810207853131220492415345638324305529405505688692850;
R[271]<=2560'd346640168219941423440994695388673674970861538480437742572954911755834640999677859370017120364862099573734273079309830555978080254361301302454799858915400500694080217996506126974020534749002830786850960670707935346038938648816460456413020659276252177828726305657014326792903421202708944826372484104943692036883251152148729822891576343403009659668970132738173260611618405632461647333494866086665805238532288292699559622362976660645775315482603585811694882271581824381451802812016984373543546228767749001330322636902684761846793767298328987523054000664236572890784735906930263137645038140819568494002797483743850899522558251917286438263146109494783738933432826148928853160993305338607921588837727226466871223965708273646183298552369817602657386150157954289541985826494564419;
R[272]<=2560'd346640168219941429855120178691379718157478282116332341518685644960692343958946307958976030395751752760495613564162285873061569569864894338252876610634171077147950755385256405782169690187035031274651970417045622035183479509786633092115102003934211530264154399232103328132909786176793211571149636416595498816974219857648635898233769469642928300995276876790785987778456452209328162864986406740948000055823008515738518620623291939154700078407654049433747566056058311476615557313004241819883869049117899086193747697224933478238583880860203342608423678508761344830739397860081520845201672410087536219956293736512943361873463539741364629472265484127319188050357392002362120167561706655043686391771932815450985636084725779456222010653679717726416352204390138700923321673549042994;
R[273]<=2560'd346640168219941423841871803414559040563734786353701479427516430380958370776710023909231036352708118859362960048527409719703492167418760845613875918122509418934288851741603489584840401440520424916489088288072869414779826743530768901587257603101409340147502736592775863431637164237763319710321739434795691793823246584612777465541296265255946276384602297945714315693165187692982342161714417127330247528815026537206841553640521410999960818004983191595435716918992182096806394203707800429132394287144058471525502799536282859712274430817238598618201313505877768945803556386301909397947230222273678186808064902795038024780627908445918727534414871952820279933778330636078893025994271535991106758235390847493389595861974191244621786422618612360190490810120226235092965701779773525;
R[274]<=2560'd346640168219941423442554528493832761650162216195837371228787610107897164055741749848768909835793370228351917014102222296401549235537070608137678544614061035056009340656920640978058369793007942125711041897883746106220231316947130568703838504893789354381152385493340961641265413288694435005024734153353116041279606019028173383921056465827028635277937911816473240024690260864377474331848239091738319284594308708731671779827227271696613535806662780481490245167827303744980855383615117131871108870877539979919245437055418308241569862042481277287327033840139704678965974316737148658231003848654813416995863359367142805220413227613662054800311663854885887941202298855349536454189413114628699363937400936683384517485459160749488047581556952408513270721165539747881510901419523540;
R[275]<=2560'd346640168219941423466043779959757836880372367462252932057512650323098710441307137612860939439260998008591484665461952330007766523381650147078312537097996550591354997599460635126256504254276236320567261547677870619668708558184419885022471639782072894073626547637716027768214289712155694880066482827359198051396560678078223169015923276125939992180440938064306292323824919536594448145089016880329461320345487146599584317409678387389784708677081443541111396054744808007387106204112522919907870646930052205111952110785113153282302659447571427117067454084762494379003776300913489825073316698693972878988612815288903496121269180834761046211201583575328316391395491207055773408083566388162078226852189150719726642203947818450156705974204319592174761743095659530682010332164610212;
R[276]<=2560'd346646779856450751857978168738421071874992090557683622324565210425275210824902107483084426232168323000418237538673577926862829091447305975004234738975272672962007157307755805216826902103928037330185670953137955312625427386399346680032636279188940785223628658084687297921614266310723560844979225032463221870856430857689235671777869826206202762767745968297663056418962385407954731809166460001515514576017149999024529491556362555326544465242723323054840639047706462391104360163183058179681623901523631594516968194026194396507001563477898573244789836890746870540370901034135044480078587511872331260520277891031721827833121457155482962548304171923978492749828773758205202379331033063279226959217487262845878333640602127226175877665589749248593555506393448423453685353828149077;
R[277]<=2560'd346753005101312549110737914697399139191476068817335459430674301700374147417746109200476848300060997907357385864042801900679764472376356220869380239787398120109603967606963192266681130674934249280927336694072416654930238810052509985065311740851759647901859185116247204536499264916341219726560297961751718618645262461846986089766860208692431850682575168378563573389593463147989485637597799076553766115362133086260226984758209663620743637861192329662790925256979937900191107798877281357396690140405254271563662852718467632246016212293903260805564389601588329439105189420643872291666410873369347553251668584594532127269364084083170923120928890516875753134928693648067075650120933917031595245641451134639573461585248047343832342830340246705301223176125174891534938743140693909;
R[278]<=2560'd375526848904936542061070959929113125243271667737286424408178202803930490995287844971989714220149860767566764421489704351953446053639879187790372014223643969715948981547164145044843857816035041842480247108442207248299442280315410681276497170162894489448953343009515494897462500667772871280565618207090033629991508283636772876879884438132367938088160594969179820330049294641820226604151101614504897671076869059531353715558123214624572055853501411550720390292325759990059026058840115196175379185150351571696399540075118847860959896885529761906655570018114836832509907012531845653993422297274358545431632051578409511528860607101053806734476550002791250115147145313254626939959595440106570453269535609168472278351082246586744317867697853513768900679579740803581754791698038602;
R[279]<=2560'd375526848904936542061070959929113125243356558062184471727556469815282639862125110714749944170053562055519536578148746815954351172453836391371805600201614639656413806221015631703404389589966066499783793091037316234243978585762600812450467054081537582666506969361034581233065856581076184976639205191211771179141350362215794119324234944626159935943372824555028088486825481234783283387075694420092562555425979101182545093399766744762687790236148667594564401481933433012127005436232854943235343831589943567212530606839972928961232075585952349651811972251301620612259312459575200117860814727495801586456759261726362072270237063985931431684423693354626862531961591163706666570047725022036941474113539195629417550911038911364822201303578043022216002186650253407083595221718969156;
R[280]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494853594973324418037622686313693593358238051170012062464041867230118212483527281286864788416228772874639601852980248998821199082686379191084733823742999823656052126846488622488741790480602482460006261545693042112718059375236352043337112670844691002800515041085323731352984359013246360278557436737379394237687519771289690459630515509745233421572971695529101187214911111841472825924538593736903265524184422899911093116161256489101373512313358725988873129685561943375946678911072101634962642841521818381033463991759447827022348103285408113136603412568772523979541130837124024;
R[281]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494855063361131593037895801483267854389997255003041355006999126353976370218728310620279818993590975721927371185047246354939847082523495707082547002584755880644674922467693176241950503125752531872141825561385964302519795291444193158007629478790612182980570581024220511078495508214967756376470973080474830453173243363727256261740842703831907329384490362157787250249012900539230486787103887151972606759287571168994147128439276273391586815657945377932731353745965955578239523714695665480030991725041096918461508253874229067344378700784221508071199078332483573573113480745674351;
R[282]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494877175553992581272394017848683528875632357189770533725794980943322421076844486279058209504834063973999053813282321525127532605613062140456722339123253829199702771355682227955809910237209825411559259303336472022448147416922761002429507537024922826379787517886068849446060909047039765420767421319700906159391410103493572730010552816855815295539070104458412992571153909747604925780042204381948401650639319522959325497489532385042146349269567847687988228631949569074680560154813355331920319795927511663128775987844321223226763957890026771118316853488811944545377060095969335;
R[283]<=2560'd375526848904936542061070959929113125243276973382592552082898034326355859084751492702076101576883111536787880956614534475375287884279663331308801642976860726454542344061788987285611944231139788827592494877175553992581272394017848683528875632357189770533725794980943322421076857001336697503031653038868716243434050234203525358684628095887447890049855679068587827060340518995435530845556785934640923981192220717886397523854155240364046246960885172841661185834369497533908589683788491700555041500200469799356172223100232742861828169960256775918733459861669754927482479591731195437587015241057983962472110925595411507102218322991528819467677184882413330145175115580959336527665133649259570925767148112441031080054342233862335869217504690995054596056326689228916579854515215010;
R[284]<=2560'd375526848904936638274513042574841585385939390720155658278129085107062466460973405550289061933033461629854640298297634990751872741010575431502700583342397701138265397156626527586783838459992523631222579702706463348540403118359670849941038229269338287636559792358013101001514962560101023381525290339120222757799010146001475316762347664082567115526842535024904775625857086810839616856214176069178972814887625036175281887941316563485488924599294999855526243361610523152242576701370517185613227985363356266553645845212682348147101344382460447759609608182784378487848496863842309184338579166849177072127720536522904776871412693935903890858813951771340582320337582173247940678295374674226140455826931501575994438224997635101970788891130484307906553103497467597984044905727035706;
R[285]<=2560'd375526848904936644287853172740199614144856102681427696213128261632665700484189713031357621256769955389002239107995907746991765745071346083533367056390654680314511931023935078965120736956280927588092261406964856636747290708534894661258092120183593800494161464679249624444017470690907951630181418347394686711796292517121015156438989369162518590241598547615056056392628121169123314926355737141835083358565723079887737236454323284970885854774148873428864839809947895686897307647063740284422723094381147263814585899869567732793203251145445230303917618378716497522255806002186604945321590720988247827257924476608712912361194022415293971172672526994295600462900263577420523375285833110604810238983822570348281163345421266642133434065409074530824607700886407595725747878318489394;
R[286]<=2560'd375526848911662246517982153134617052975304416381590896504923851151332796304781635856389027283550332793966679240266554429603083007597096659450916058003011348561872845159795094992562156833156793872937272872301359058512886443561627221479831225149912647365361302336533837716967547142678569852959332098967882693479709145762774094466429997123318803274272410096659593903171572409974652135466483983750632287283187925949530151983012882033301375766536535641232878354308158945295794185660977257087236882632494274159454151658712937593602219041110994940542372236952199859992588977185824163478011033538955858558549739284102028501016049533844846347531638563237820743755797611744334201056690747920570013932101402894492425104098979764557730484378272591698995743323063675389911946208177286;
R[287]<=2560'd404406917953422338678295327520918644765738169333448693901246192958099761268385534562352411921086031334826724184544445157628807384759159267423089530407927320391442142725679662140427581561749684960693807719528874284810270623158308247948934629463036651489843851814143475510170700392618020734429135306178452932773324723480878957476221233954478965472168072254980925851572435637617322648423178888072247338887011719777440854345857986430647686244632920796854622436879686220912320364767151529215896313615876748466984432316175992525821023686569894942464055092259455111535404889841644334794284823618324530274775855406100732914016245091150903166936494249944929442676210137180584586619866231882112019515461909341298583647950156793273249228079725574836883395698097604821267972366440551;
R[288]<=2560'd404413529589931660681153339969057251803798294552882071480317662181396680631593414512921025891802237229921890829520912143143387438132091166917410186123206365618983733026977927446897035443097079799331147974738889346152543296373643308062912169691142721569695538994623060524531230847093599000205146838986055434479816355706378535943935117401811853623858475654717968951389078516570809849254673241613551774405823528382888084410886775976567595696995071589211699164450181334069603966757953211184340697574865791002576247347208514413290913641232809548945503087350498351613490302432450956671197569473613802907147993888217705555080633731168314728409518137731291110802092177364189240660673719034388780967093339207847786681769709336116665307868756181407456649977518465275700279391467671;
R[289]<=2560'd404413529589931660681153339968715438207688671930850276148719930130964996761180373215478956642378300763593738147011417367598189972055709499568907053452740900893048967382217141932486495272696734262801068803910781558819925499954481574867164776370593874483303062618752119385049767915322959482324192601067304652085081435561852229586872244882545535930579209298304954394129081421400756758874575884476976607692363963428402784776185242683018632584868627875166860896160407242500170798797879343454717859425718251482352798237041084811452126964118395702430866258525033814463615471730422846614352540319111451645646523209549835983345762881790419055108276608730618968130457334899592726422189869199123171773139236377435543824431924269692732665243848841591501848427138712595949752926381974;
R[290]<=2560'd404413529589931660681153341462121827184982211345178075547046525660889453344265628440907000880542374244759382731728703961258427277122136380751400891741209860574247691838276737552313492740479798213366684542976499548679383671903866549740177015631899596955149482697733717303652067881210853607779269548930283865728105598045612017444344079128790154766612888744906274003005022219232220398282974919405365541198896209064383904190641581182195561577526556834478569806260991319809583113001872630858597779015181333837461920418339622318965486937997636860504591205032914603565875002590659253550809338374523998895462825553177761925770536854742206013667369524415743177262013714217582986982562597358488998129678933277748039372657201744909472254953817493332324041797580987939467521100872295;
R[291]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161632797304173338505320360264687648792156264386749475057482385742176279422131287517768371354204537469586621447702483005860541522903143097493829280059111038401930075963492848979250059492526998407693639130213459368257481439999469944450927663258385724614225000101666458721295390321395116722785825634165992356694083697437296228089626714022808571889460093281516487842991837958042466605864670641134853478640159108262083624156593887025680011282893368620576538741271222416735161634439360933634529764924346172150418711096566024701490607207823264589050862751628250571617184000450575724453;
R[292]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161632706732631379897511860480348034033710810823793173432692340833814553048585908025066517617754971832937943883007598349334823992839664322615512264293028367242808123676638357649479909180341909490090328835571006317978425332954918686811463900739822437072601074878560220462356132725811000458850644128372768568739385669387531225796056256381514513982994977253909854247356884683186563232523161081071310399955543150575610156681558175646035157482786663716294103326535245276798005692530654105447317256744918871339630037141154454285420711957592097414272582845067560004784570731198322356114;
R[293]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844676142733623174940827834796563416718013547270614521238759817916105108331283439886616553558245742860461898180278185985465142785224388588716628434724255262019740193667104000193024377774961497329224485621471220682326505291180046918897359852794380948366306345280520167420503641409945266640313228756897370876384303855036024369114239965388963490460238977604448809671178230844407620804690632092610986863113583368508804442343816595200311903772140995375140705612176050217293330779210475253642881166681136915087561905755358628676289744768980096933487485918956873881756878499;
R[294]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844653736913811544692612081942423866028625065493264659036889871519715438371601485240993626306941381436679663271277777485736367596314558173820325567892604219160749256865726952466264160709125536926886936575971917995679237469213420309335162174530313899817110737947230037191794200605581120715679079182413414314975448749131520388966955185416991219994806043812127674681138240798391783686864739504238546215658569680400485547358388880751006896322416388823125330623052442086298591610554300011778947324319130851030758648329772449936806356543306337760376015633336958614426514903;
R[295]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246072931639215390443848271533286048834924596025928654661783643280296215054381330893291603834399348136915163182286185759461235032146674305013893090033664028443071675825710842293151280235025867366856139856005672335579022400805886215667403854500264178505191106733682106482612632688337485785140013975890405545244281190809606978035883853798216891837892603529666910396820514811438333137492392068906956670670154112913797422316986089801411687345746609574264012683292582380322783314236626150809727514343016544167582017600491487222851065024617417635661678692309225368551849195947110;
R[296]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246426640349237838960509550446830345975096606929751977480177359356807724041339168177124908860167697287170178778982387692075336690182594321175979117171653857191168333357378346917526828941184638801538925922326899800810784054115907517498103975445475760335368140951674352552864728184579919532538239630534247404131197087148663516348606585023260962098586928743765170855990330363482903134206244768574089370720101608846867668523874076682853969251551209316354369042672782999950648470207233866140792826686164472233142526528019326394708274321469717493405359801580429766756753234975059;
R[297]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448838917852190430297572083107538019587064486503949825140062310809595008755341407523250826429426491735622845468864822380140679601098802283362650580983060204029021490553945256118245488681051596068002975106981513048427293811887830174721385931332253857531363996959751079882980199187785035333358415295048666220592175000598059815572658397745234700449115923626238814766517131784244210230475593092993947998788878581835396027901457227734960998591877988481907966512658270388611285543139947224815968950936719889088398949182509394729585307514976922430579248362122533950491407740724;
R[298]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844316336775632503259831559940060471529686397760996388758986123723960539895947616719664172904749838482759663600543969309502601039572168779708238688985330340554455575577205547516230874362877110943701699304768958093763791228025320195062958053733413185657354192572148800684885280399326397066358230292564180597431077892713156012155074289150236342508573776445522460934827473506206260508101036068841100135815888625837984504135623511492624216850718482219884081354793607876137723051290963180571289698774535415119558016304478565194052326189390230524514339607314160597773278612;
R[299]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844674829892618587231283605607383497904680299009768927568811248048903997053833185832604125789713988795172249935638794286551859051928974624350949694873637555454977353646964454129466334746320573493385922572249893927569605311366339451140063271112796979829846335666379983470351014844671932590818978424320050513793320605267599149265745189732100905838274925569399963343115827200167422152865702361681716298393696339490448596499015564591251495399931194950407318063245989670045066083790190961829692016884752710697747248808273415318970305610928661319757696753427085360148026982;
R[300]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535541563654133905800754206988663969067049801960913146019697728449270502074954609083448231962077513974345785184468028484289379250268367429475595505293878581160075811266576630711683684781921785098796244870244225628583825261750181999253968155271096271460772895972753755295761793806273807279571574173842552598508530817312029542283414791206787015916304316716760914933574152861304574526432528183985353591187742106873536171944595916593427511348441189116797927941777803190742776981946900590269990945014936980366832002032492179577767255364757035265949655876982099774098556889659171052191790897781;
R[301]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535541952655944566313077403875600004954645149336364241453498937755187716667208456536884651027007902291689519079404789068466565998593154692378926880264162728223744986394398752962113521719869885249051322363515342208021626983843012073333218370413186730763026791250575931239347412779968060258539737308075348116425753427607020616586340992432151058776294367380150743163907205556764369915338169117339504056060586646429755014655373166214539121432131776506937088459389847201664339566253310517478705603538449520341379972076208391065245867481445098585280144369473802786691889188296032177547243320883;
R[302]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535541952655944566313077403875600004954645149336364241453498937755187716667208456536884651027007902291689519079449819817789316740407910720423258757347631126605825200585407029541898255443844294811222040611150727664616701891938805736741273562927055820348013134799549628915464347276415986052048088863332730650600603805666045050863275322472868215442530973765524297454878968804166625452077077155193978544452696167620954666989720043868545223045946560376915297582976312465802062537773272989354887750076743894104684632080145926526993994408327371593237189888439482413568077424952443838917198376882;
R[303]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535442368192415475158339021907805228676352188988276005872525238499602416995884217956468028100870434580676080525013723908444438088927202157052721183284266781942399023806495100232112856950176746455734626668115375671735225134862133450728265228556486241580075413057631594554915586915951959483231511073902325612688312768983658526538923319382770444743159734128301207212125225360993263307102420253161764574683985175286934483670602429568709626885128287827893626280844729843119869206164497911755209380730952764976736895240998711785252615520826932643787683594531266015623842138068934709523057729433;
R[304]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884786918772746607248630063638125591701522177586947813585754063763754119526803657654198388038233665292022769214421311743688426508558495535451173978779975903949971957786458063996055333194229874637484765107585092761714103963865951395485150889251432732140175175859506490182444871042385319656985626487240037775155384034456472467210791457117291804199833082825577587295172264959555652468120986492478922377776573629201414219642458551223195494021704488755664777542795474146682811672253774138269371973114711125909138662209312108017744008234265230824199820566030134738185355146330487799426904934787643751;
R[305]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675970526915284467228490168625416888505441888996699767798197702261641219170657290040032549711697761062563939503018383178442739468219722906316537220457078280513378718184247729520441668702741192181174309718808179863229875514513615139849634486853993223703082858185040903056651581375775934442247606531352321116180198555384837762945870798913482241542708356182119994038885497856500627660252751848190410852340435378235915724111359650951665662219753201861111542572063044720179514719793476025648750940747870043830567790327562662519171081836105584836992003789689061656157472726739872046686530224952567;
R[306]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675562628952669309858681756085329484869553923410930354858529430110763831716913208814646062206238745260680521256028418760838880638831308062801231851089586049189443561434854342949528286366516080085752767401756087043957649476334537181793978744266246397429071335757943377170860127453678585926200908943424929143604529809489095642369962512811771198504290340357855872889900933688202518531669736943557659463852381278293804927004084354305832616264357369015793586582456788822319769382271730064119461525050633526223236366845818290847049824525417451021957841162924737501115310027500470098840917456055238;
R[307]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755167965559517919196475625281290551872680513179379522030123885103672500482379145671718424229056075155498202413012573323302031836317168123352698286565592609570543656776157225222983689259941952151287059970039694941414779038414590882965184955264434105330885337288534540578996387938028590730333441960204576323107197754350364948204260047779421750526492422489894097631570377003406638009891237305352973564661956860761999725075895176398380366877275306642231385177220918616463867572167202764447156865863003994010847802920469060543092400737812016396473214839426107974666888693022508868808617;
R[308]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812139508572253375677003716853745000899127754906748380433443460511189065738091329848456795018665833920600786440269700206694275226284331302380107852731359265431820903647818783597571951136860503942982543211022443623062605309041959371621396320950430829374619269505677603554630189083588661647807036947321086722380781837777035217152538715462488553605089233959226550469198509035197323046384257489364191830134214167270826092636528921197630969917025546996370314445777129028334820644793872536684086971224207113948031625439012192774077231295043450107731515891772024841476003106313158829085760625390204440450580560363;
R[309]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812139508572255150848937018018618407110502215287371764859672728996302502058491948238655489260158715914224540885598980540752505679797955387736641219187677682346200013104571035609211456457491277970825962791458203330556481177602775599305416065985448719225145333244759887192089163217983936515132713837309498412937050448310623989133632675915873779188269701242610398402537875057088611847456436007857594336550773620951325665347424328750263687455799690781352815782679291787177974497140336948697187052373617179350164184586129974440961334236409433854148492973691172910361767176876073949755602189314994960418901169515;
R[310]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616781760445790646618040839865459165372038106739100361418941450962204717301885497760834754816512346519394863179203521381114723037035913801363634817494907872434297995279201274298996159444093766275729196060338852896862374770582400413243630151920722123612327368949584681219983710922798531328996284609923855314978922612065551930961798510450986946949382887384955037431016490627578746346622486951467998372090395389751873898398749291169747465077592831582547575358148934597579751785521970781364073527007553315486516097533455910640517262951824102085786791135196053940806695101814009162912655019394237301511975888823623643891970907514240040334943;
R[311]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616781760445790646618040839865459165372147601014696432140017732814663290498104341781313774052165590006900585471873725661042276522177816352662397657932962621343939996721145478263058040764099214063599051126673645006989337860732446277439783636088613217638013153425357216929690004644335100804335469183304271673727769662034715356700764623240752357140142767637814632733730832382553406435502824472505506326977363687196559395420213840121245048265260847974711885292013428095519315024871179355608485995703307003024342698236567750050015845196658268095715874214029928103385896792262367569543291548229883499054788685003458076556137886616402883663144;
R[312]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599302624438591986909246128863467631482100141953692261112452278383727508082112759455340313904636544104148941974123101011438710890249284387064694837438888345228445060892796927760058461083599318802527780713105705423019782426119238169411820451565317016103469735053499552426109768074296257964114346522453177306389675039277500542925866826848443877266806531417001610064095443968836669023508344287560849699483247924532267792703320606525527255702352123871401837176625419157093858891128072629753970584765300449922276457317628444955816050502130247608975360090221179912201691260532443277467106491185842927077646583700735073516446248844916185947461279791042794959080811059;
R[313]<=2560'd404413529589931660681061586573583057359943787621700564892669300699875961960097390194786178283224806505599264804503280588086674922657743325713196909931691566316229483773462487293911375321863444426322534560611297044187445398426888869199527686209227041187697819197545697373933634981122225389284758903164504233284399218757951127125295704850142717125550802069696633508274554777737870032817120502840331569999358733716408135757266075777176319033112444318006908757956383516661132797053426987096340984911795823943672452816783070548019350060933253294656358833249543264191059651590178981132132783905393510599979629627425739840098223582345637903165393777142977340146131796712761887229214853113245234103881093450211446604003114462996504706308202251482638507166133903735901815550225860;
R[314]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891333810565158570704129969518314848697015724982659879427559746158009388013601955764841113616541325795220701273398285045762641026734870647355774403996779829187578179413675872955426357807525529716092268747229050198475310135132741863480836042958211061239005971773611120887802878937606145157391085658988934394112569198360798466675926547108767063069102947289009410275711110880598481869944744252569411832250103536446211883100976687584660394386078852370044331663572593532672070029623769290963017469501148977488560804313771305309390590912716141021513932224152490978148100733027218185942583159357889539857457674159913416760885256260563514521090694199818594922229;
R[315]<=2560'd431494792732114584387480574149317485255490041294284684974500337501065006291637059915277668864186200872780094386098273983693941536094621403663692779131675953962003668961977645849894000378519049692837155687305256672635560103681728419973096542336738908224044584211322424620156784375760909532583189762209575244450287752245065469035097413306400416931705946637759308027901621823181819086661737450523752122023926936423322830818564497766882774253010813328877019084285737509485457730026280204382250212817608719936173247588114356299450890096777498377744208455986876650857206031323064661852789736136050456799010627912458966191767635010852721088598248585939415870829994608032169136028143693977998040385137909160309669192182401884474033764391696778074615539807693521214213139913145236;
R[316]<=2560'd404413529589931660681153341462121827185061796024770072398936659000629969094484870217245482116916839127568920174112160645243664609048268820276378026849757937983240807293048600774666637599040350154898055299663093376195362802633086577109499460894835153367592564536168319377087537377624311717682735771643934632044634905481065652906064632345496543449961382145385033902918956043428158319171798598348799483685757626548952980316418504922615497481807602218642691005360642817284443922254156205167105339976793284302220085086453832112259180084010735418308814792344701163555432982815332005618861641901514419676448461800001555929161099775570892629515263702903032908185478057376488766233672136066752768958959000685811208943389411478172906051863437432203706330212970437498810548184561521;
R[317]<=2560'd433300210274926779301235722995130523563559176473396597794481591035129169500099323929517723136182285162502096329866484160812527451337011599712092149760715004939288387712093087940495231132312223870148741971332835985604474502680108873760630159979910139015963637591348460756405824472552388577966140010442107876030975349135730762317010315241725053699913441611952847839293538285349846843617288321542930872882963154494063950126855438745928308648722665250910306709219054090071216608646464368580396170717885261272742680932612692339920264347658268941325936221610056360058218695147139690013470052985540534492994458221012664296595899995712879390150357215998323918004242660541317025263101393061308980452171706248094261995516460908883347006242380798256561637953593600164617062116966693;
R[318]<=2560'd317753487528640956892551930832204555597846079656674801854503038627670948137425102346775266764593919889881439196463828188569009415156449992055026111409179918129193292070290047246652767743838143641120156126220495202066788611444422203252148759968195151615068063270793035105727439671611945222186511189885028335094983780474130707679377286477215567416404086318905046371037656988629815706555024123081718781433786041377464058996450254394474917104432172980701567635004566952441292348845721692593123063773794163916320272677173538071098184515040124107099156477709750783618749884739421796634188491734412672250358687464094006888413905181596019549491099833695218970062338770652615795141162503290313933033636300745561320470797695384050839268631641632895154618000231517191094283369214840;
R[319]<=2560'd375413597081230582857346831035717323606014621746355866405339981407251057172005372460804974842727197084480530474266708636934391090156766453127377951635945976145970367372055955216571093313714004428295503381572485332940164859848030008368051020364590780758230594008288413724944343710124723809234884958625725980294811584965055592069662730157728778404107475034254253500177240892335111460551882273083713336707857725687318286941984276240140252306072741180074175735889320587868429254628572366403596001258264456533866379781835857952105451355334061309367284523169989624078340338183379260557351682256984019471129631157841478009913006988541473502588742079906435968617857062709960177028282627093885268353788032659750757799857682598899234024759868006008922400270320720124186764285146497;
R[320]<=2560'd433300210274926779301229606002561277805177390418715604256895368230825532602404728680887210441346039035044260345808895320896412922180909825623743111551747626493642125548271651736680456922490183723781949906467190077645259274783764180421810750283291421320480207428155737375132626619475370156652748794020737066844813989899766333024163011016530887560502685983564690564059801247429965343925316494628563140430074819702592285028019317164497227218233582889483207923813043059282630262902820949557523279690141046623468533709895680384890921497190544347637608085367561065695657796892375275564364052207306777408069712719849311964546357005726969942538034253270554924315261997683300485322773735605009704394857306304011601299705718780024737279501588532256418657404541616060207437469082021;
R[321]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435781088756880804280279923529145790718604549205254747513074568072283939335739006254484424971263740371889830938669363386336216259277288819111376472204431309589508049294954013528240141627611476064957959708577920238155587186774641304951942043411197260010688980930797275062441970370893991647265950591111515319048998863023670834804930375905101669067701114647583134832245506050880460561782853684697102747207852841245729632800553020038830415954321357532951421464701664954747092591697218761630657446136534165041159080940443405716857182462394703129492145049084857788498680674543740167370155580;
R[322]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844676230256356814121797090160771478476203783411205689585342738237236733847281189332292116696557170201411928063451682343754382614361736983243934457525582285813877424118882692197441833432945977977591114098346334725988351222500670390530248444907503436657170202865954295909086951073675598918130884960278905050930498781579795601353509813984059071195833627820920477091454283402556328598021099623050655865248402985442155412059739903807327660778834496841024040108893366511639520865437445803080282815197282836465593281219669361180579459002541118353159742438314786263891432269;
R[323]<=2560'd404413529589931660681153341462121827185061796024769995191709275443957812223050393615352532743890175416995628512599301891322624103246120616772095490476161199059776841812017041414884675535435755161634246448844676230256356814121797090160771478476203783411205689585342738236416547811820651494317499585084651097163474719656728147482114369411885251926130637118315677630288869684722708618691755935655559047844656849999682519374482620340038182351769171003298699284489797428841724780679193982035394844578769470321916699678920898091105534216551339962891533730103228980609650753756358729286869348076652347034742308664589394490373383404804902441402993719647453269823973640100966950869153711774290479418118439174283856417977187907252791874312301339506869373325035763641844684300891172;
R[324]<=2560'd433293157862650169164853866944951571924229416956714629858109412911574428452357581147698874498672371781612625910044442468278646454369043048511802016590486675310993815989266793517876318014467727423542942026551479979241488980678095210502005116288850174684288081011110514707599265376504117621948428190105467124963507294445189025304977928501759177009081728845681652868504440009419965434965279436916830429519355545416058909640581420102075135127222215777686011958702137675438704128280387519957566911314019757473306431411311101321789080285849392895834485544209734551586970275384678268979786929519467000678646979942857635926066019644218379965655029227949324002341210003621182130059175033525386662533945794228058477238246599239480246131266216300772678022921386751857021485399737959;
R[325]<=2560'd433299769499159491167711856991994344301688017602532382750661244444877454234461360265723679064092422650743719544979755000462015507105105988628958542809835193048230816212292720658925537712837469175434404640007914687039442826569721111583822345721498768966541224091977579151484308602565284149978143570089132494063307272327845766506530090876693863827658601028390516187633355938789869743237198519711591268102409509209528965144842023373107386521683794035492315036925606804395137575433202323951928532855951652940786093577553304941349361003562667799348982235013527747793603121773229301764042365793611052471696315632636277752138251546937989213231391590120038685696210766011822901881351386734244097761946172319329142025436306680204791208798171073121551520992526513287328985958128632;
R[326]<=2560'd431494792732114584387480574149317485255490041294285843084011235853151415720129661044952032704418535377955157207639433714402264110159923336645226884927689850782529755326214611152488560057897970909065111166401239371018535685781308503610491652312494924716289418145608641564997215128402364017759026202885841523535605982263142281204537187461813863178694965890085178921907757493233899644594694902699658274407781653441854535675669752616965724361475257905714581923073874249175329668910693463982344989292622335143599821197798185210112589169645007999945387846464794753253096948521008139888352961123179681756684441091016502730063362240320126364696175964941316416936183907833036645667601255845084405038962264586864934652575304531222046751514135671250846030009096571842595378949208825;
R[327]<=2560'd433300210274926779301235722995107741553777928745607802858984053485979536310116059254498349561236083454375312419469374466026939394958948285918738379828006836337920358634704735229903905102515909142671425242865458276769724983450076238905592143125877398299086793049108004784535997388217522051856029370276247348463165011035225557159015918584822849725971376838685423051840884836514170390340279023580854256047312744530303825751442650705870787519107908472402567870045629861455080108841985359166614404378871357870852082005866830563449590535115355204397567682801733050354340144484212330192399886947026129515173632460196850416725111470435168250544285803719695917427317994181063606112717358720176255169910606106731711970962728461250611486735475247684987538732032370024089249076334506;
R[328]<=2560'd346633117637056425584457773547598638740955659636760317999214078495307508755185739537016615801349336167167624635431561527572412018758998377300717209984330133638438167447416014164857755545574352134491051417548732356282462517301761596437137128490068629300463371217135465075530036193901624986239499706257176134535381004201649169291840327863378763242298568456821887036008486489332528644992805731210202923011814586600885683834358338440490982508834799900417374963675929329008744745541536844977933257958479945863539602855437354090969584839412637295592648602300171226151359620281182664177399264461744497688028135792635542482347077476446492212326679036028626303647897637228623807500801894456552106660132722006854193085377627093677665302358845836683321606586793021361771422672935607;
R[329]<=2560'd404300250325349881676099252256220749038061102658337381988131624134960799552582350829667743034241355011108365134803152003261052131281094648306590775475239958778992832510889377272800566300243252512793286475734726586530372887455498045765117668034854080166097891423394301800476745539947630909891272329210218527152365486115603927176813130176732215816647560249208999197049777028802221561675514320905990231403820344669521227040001006531531677087732921571207947048512073873998706788288060685546823399392261004939220781196859006021929094442199761185651112429603770640882433779653415223794901740219609241226133326634083783101718817861117976677867188059139696424327463736687729450318796269978408207841749585131096460792469776046497880581093796691061787422513873611063850214196005559;
R[330]<=2560'd404526368186357422863263038264985142427021913713392977891260533612329452237621557229627661075152904778704928643397413194404098324773048374310572934513860259541973991057769197030268535220083502275894109504197116097017128932315453966524343079616991968565875545965985561369061505947159942268968290633995033299003406730405246995734488278456053804541313673778444443495845244596005261484546370272567958275883378970261116157118699204472264839587269264702803908049374436715851220145915137640401635629012460793710190541251745418436150840883752516743596498592791597172330920859401025035240997092001687616162158864731752436671766098698283950380528872990674233995266435055324262100649564531131978486699956754251809047330552624418715528190574867213357974955642579021543647524372264879;
R[331]<=2560'd290785505486316415470037835398202284671782515390475246505358521014301627001719993215521777430072429861685989365446030565084872049594159725210695773449283756055331757479003589558066896629085444056775802647330529619597666905761601133694935334786619503668706795631430643272417754787921396730361606796439182279779656694170031787888096664461170008714395650488065022722414379521860058493249137209969609382938984540618921133977396150834120275210056202468602478444193694626144652645260150081829702260530562831243721627892495953776735121798834637117168420029037084208694903736239283039513094742843801703055962723188385607590148774769066412762809184413775639011220916147229103964593836705615731908456999454972636878874500704579548645483650022366630370779848052528451424992300623837;
R[332]<=2560'd317640678323124956900021618486922458200352481023900943273916685812111872287193094724120787269541878999841065511572321029808558266361611476126582137421668100020833020015596031277640273626451563535552275218791149969906998398148222759667253104562543734165596665098400557142628969247226153049122419114269526497195597457082733090386168358559298886449438422878740983992090814201865503982969067469692131450304319822198277513904041878695871501859116893657576897392457109345345355210234910182990856280529931210844376258722674526605156097864947374063547508169124476221138764187061768776438234506220325271973515771072942815033464223626662928018096794579070199198998195970903270376007176516109198607411191625816968327780255531164383242870605687807101527274597504708975043594058833615;
R[333]<=2560'd288866806850399463467726103192287374466697981464853208674740201937540775869884007675146556869822565364305878895709958181817760636290311378209793481012373222343186767959929838068296256258626848052641524197045224947625433037473236885093791913133920511476395276081667597833362774240064161912184987892953703095705216766501196802618235971978479137553512411785100917993331139337464083624053544397089720984367179660086856148827470240622706844826061707225095232431391813541717152594878442257934807251964166101911700695754532203830913366495810279611802699124005507265552010371599388040506259368779903213854931141481155129814565232977844587042097136705658474655644266130224059118510642889890935658019404775163008658754742516926687152650012618168741834142274399465921132306522168063;
R[334]<=2560'd260093403822096123426765630247844189281134270777768526159257553257896958867218650895763881315600523574864283395024668976891861388357379077026601999692080826489696662859456579353475128368153939861533018529781919447849820841959485312309102312454707346552887459017405871711440750112998901228005864380423046834942417942131050494563843516295526308376186081773252784929190455108510798467716928423748416038115473069355914574395373073090611551288102978855465782684192692043194881317911902500753740176727222564146707057742508266017491568994876481309935085958416166310614844364930346799289820492013297253536393392290149913261327979994160507790133255138127905964651312718547411538812678702895645865698813169330004067422357562522831125437562463430391747487878828255240217826976307965;
R[335]<=2560'd288754409036018423449219204706583623081419355215888099173056554009991689451921694151949152253947628383924743426385907892931393712739648496387270321484383995062727617095431984210361923806863870728983103107620405282645466776255146025184273118034239009091624724800708885112313344338706466716527413263683906335097540291951960737389046912540326917706069999148855497136588294219596000054641152839357480801721022378666447460455958879397171608886337709346832606482866851230146100760820299987225005533666470285128703940330366280377807837499826331467249577166208097561167567742450583797687304278041579714188688084703047857916646937094241790622193554130217706817969201822347854863879606671475761113136855289818682022120824857343648066818357450331560609883549527050425775458032258494;
R[336]<=2560'd259980153713467897998325343683154614318625539291822060800258100328369894236466437075483257669647425588945233608829916564358337407779912116714301128389929957933039248374731146392144603694922320930884199897335158568683335054811681980508448420554430056243973216332258413862091341879561781338081096391918315288356775730706790043302318079302670217432617743079043976242577199794115247228826588345386140533647719200938422446173259604238318493427872592408308697909869409977146246386727473135738180802000931678331383579138761331686719903870146848668541854565187848955490565531719753908631294155389330913114656409349404893262262008656159643746836054557889975704644269022767951973024544882612129053345238748049881129176372869987408362803063364445264054846506260391403362821004378086;
R[337]<=2560'd259973514535172450036360634841930539436535949338713415576736251562922241288387574787557096792719197327813969708543695869229604233984118761523826483202934971927995121941033294318571189588143376364422003852385537021369752604827171665940380225897023397160179900580481757711134558262703072274469831773690724275615148073266940153608226036275958820457697603033147408777194022267697691171424966124765060066301345272997123769965345884505709286716040109858993875152081122779653625485267465116805149121336802212761441763766096556249900232266431597897098595262357944404699878124959568268327523238595721011973567798413312587366285869657137071120643468069205580792967894144545778643578748651349029835937011910210992050720033360834544148201135790156218496488647081107257843486779505143;
R[338]<=2560'd232898863029500490347449143702295660766718213075307989304571907620178717968721413006862097667362099000486504160063170780004734270411241772651284431607345934137115471501546733157842482522445793840702264100243907539435764173160108520177734765879481613577421279451563490030810503096954133003714069884305135827403395738162133205887108336476064548560587963504542046520787302057876877984683186119803875260282105772230856262335922448471843521154471127167526846184105657852561907107644324719834957978318636686241660694486185782553571823859617206048000446865754167936962935988637701715999841491863629534397163175954027003620399679846618404804177319664546947002131821371286220200966028050222152070246968704739263532071400139952031045055738493176208335729853991378126231914024008111;
R[339]<=2560'd259867728344325507431996863011170381769443598006806237404419437838238401031893336509151502788923019394442898937433483375846379113496707447092368502640747668273746054070290394608814163744748222054454082372822806671318944463474638097965374149668218657107909224114312618430982957461357642283864790127467994913651648079884207566400199075542726157095337181961484489794020290392154110146488017350941150553968167022897241140353290091286729599706844440958353575314049466747746816617568926967522776460170436899007762329726260316854507257894261197583607893450209406967729351534013902535709245644208663979109146912896035039240864189768018164756176991791168838561447800960481307406564141558489937806389674286533912376502472444811254869227147201241588645094938261410882348688242154447;
R[340]<=2560'd204117970338287737194651345491710339553356400652397168817675059860073059502727126619360854184715202046196542309021369742474238839827875013972192238476913700885366996409855551509659826843078136987694945200801485979718886574737802866795285467115341198239828852404326308395580294911162554084047689013969203760807550855162892649409912179502166434188616473856609519451494969545033414760165657604592391393594375181544072220376645564424589285382687163910356902356162462097178654097976628129329561581629282373176067320996833099662047844229550055558468149291405715003623872118659235711942775858806015217095840979590248157239775000973393399536302772226537743056825806417758126890462699444851952135253934193388087368937173886595261470443567257522239060951942839487866895326632607595;
R[341]<=2560'd286948989771425881125445867288783282356096571927165994798579090108828987102778461818987380986714960616871496602846836737845706378469120129202391167183506810220697614983690148546474972668138211800010701348637827913021836308046321715879009268769772288477931112051564208978723425426844650257693804980465138994102649858809002129733060392870014643120959382581665117700563931473397432250034186825208367279196399513981958099816141405371786033142921768489346416229673627345750499221727936795117988507509427503017805777950722207708992451955739740602678125308969466126468330551395969817645946481282182303529380390319855788190678395578062962152747616284323022441754470204681416677545664001896764072536750665514926025409674482880107906974248461749768266701965101502082584233951358890;
R[342]<=2560'd205929970260374510419790256314965470537329742921112206748586067058316465496242435629322036930471595604751637568910153733373565944611271139775728020263613348014891494483727936075183429158702263047103154390545396905060927176606175222649504912277514229438321698266702270824860668616489753597067664127929440546748620078442213704991577829941608219113854194768919442453731286596958776342628602716288403218313472438474913985187339240940215182545192783827911775737106391777777748361132734179348287302556817410495984036856681443027211186457395891770065975982244383444783662185081353019433470301100519993871727117901960186375630339217986147322103383803866955131623433844499345869366880070071369884141952856050803516295434497983577486776286860285232383391690410707275581041543937976;
R[343]<=2560'd150326718018552426306521993418130752892178764133379066002736153074331546964847293620299066757736753079035432245652916172024584729076936590860395661302454573514482156166637666651052380832228008738236707486834684192515046888442421370299377442912647414283296998292722084379855543429179567976082568554229337372211416321138571420085714543936842362635603277898377313439601893473196186986540085158277625231118638095298257378803181076612605889919348189794889742883868408497464324592752296518702138687950480351070709601030513031831030127490734287889948325390700995828360250832342473788803856038749730604744814527735436935964547967278818041776761218837724415795618282698886778404454860786079651022512266115740835871610657743109795884590442077419976306678885805123702189517631211;
R[344]<=2560'd121923596667169676294134752798367944622349575864731413946524682695792054026606958245036083315470579380851136334436796503224518191758071348909317934231211454581950351174363924050147296802746047941804936273071360821177840782591843810015060847416297791880886602355693100958896567100030126692749796479277641347696872425818687199463438953053368600337608304478764436528882538207429474269825362413774705564938702196191855850787405982756584274283251615877939048663016184828951185481801952092512439204168014757356296954594680253914988770323431118239125953197370483396474151410437912359730817625247700383348118863827860430314703182175337273677444797538702402624138899179621940279063001862786080772103530233902494691132745167496211316927970830119019079689664232606195073861578;
R[345]<=2560'd105793905257971206008549659007166801740410365779760926759815880805736673310563983523959714590906496315108523129381797560699087396712681600283321562502120989121255685528237129570451626998711020095080305480190139736480064839200667258415403644685546475425724373264195072399168780706683253283748863945923002542399573876544322190505461834774051334961433790602504394754948719543049208129152131342389963968071386912793097206644402818042367188008254194532427040467997034029675346313337716759804394415230518373538651059412622779367174073607996594519567638850355317628435444662042472677156545144545026154828017550507893447010326171683413278947579942069313368646386502057271281869747560197049293141271886021949777113294619598598250951920769760111688408896604815131439299949090158;
R[346]<=2560'd27081296589112829943597442389342596363143422228314674255051421046265733304763889582351055786178196464799564804695240966871862658634740541764212263140518892711866705319165451685451773605387814098082655255986929963519539799951746143348991242007385502358143889887603442057507313447221532312779345336971050554394949094073578225376112389846530207060533740598015642846161478578342873604647487974879993476614046637242334028535702614360829258334450459631579497418640333077034439276799189713835553793800838438362699252505285258507838375059632406959435587414477398402988354131827765795177938974635420884827734117328225086568025780696152537386730138071027896403698032949934521126582358909029084601318654005749672559102664852754255818190781429235137148937960501015701019853510561017;
R[347]<=2560'd112407155962532525955949135630592314026079563088828566222804073560207152941579972977704623110106087903863677400258494528635702927381978334228071899234973568451870099941931277922761803719202730310825743045735663668702075520885910932399272825400508448742059236896601617052259568074721360919814159539132757953920493285768298741572282198921069510988001784504105730617176897028704889409491364188570984983629583637596322478951566991038394832780703667482215232405196743042097213427648488100091236101585107867956038595627155055918021531678861657389548798126532600380799265013725735058994923526797812185090410813408551011918469951609367872037669063531522717635782776030136921902237370837655720038720951084897874751519128833930278293735867547499446815193872844420914884861382601;
R[348]<=2560'd1692999895198974024582285182675216451853470162127153238392739948774396004441260349495150492881494428127993793894014548039177669474885185195527883098588506605391280686650780234493292803655414092480686513055273683690462604406896691886907575094702144388530394459039382515260882920794360881678631151979930218693810155293436353883466315871297103028723494117892325402234615253208343673367843304516375832708358322904001472254787174077206019410702321528281710110078829236020501316774123056794046411194777280619277895239899543626110084662681700371815358162900315632898890141712672846285114180377805748698844547900150686132058732724594917360042772820673205635872547001842085508400751948482360492843226730317126156521489773933734532333555655165312442442448368094994753196038441167;
R[349]<=2560'd1693030570715009888017321101032297625663912598853154232497189174803026698255680171823479133095638557460044714190301224621745465452839472710367658795851430593019241045278092689726822046979691208647950100499090539952534708318002869766228017193732797028535813025221159738061474948224905745894501442745321248806039112214655265003424229514378949965211552785067740169551785886294214402260945070054430685431084336615713922124683773555100141667217137399174092116044346606178560348852636115951831185194220537613825543845526699766096225470721260548175096412978606422928348125340424935635713891142692788232887816542835456375556232715155858341642690217766361207212055131795518993329084826061561297935834802948588889262250508945192460337780361715696479713906679833832813994702198175;
R[350]<=2560'd2728813343598131202768395789201858794592203856432392742334877607836741914047880082289382250000241653722214710388048069927274561104482750597799115826022796387383655302064600364179702717947932365043965606676264058704998256376876501136289892712552011972467593283768868766364466061972313530463562633587945761064623675782330077107670115699686386926029178270570142122185562196239642239090296373153945137886495569146361432668732341953711771597537394599089057388360432456098397645966590086106075112243897657014238223032857906591327896691638399587578447821989095620787111442883183081240236250591687916132631225368271079064972713452107656144401327212796953762221030110447844455642664695331048036665229794726512567275363108276027484752101188627116874118173909901652045847787902;
R[351]<=2560'd12333113002719420867311148689805955433277406011584327649923974803810419353893496966109616116807410543280069855712838669120222928735306714623817553762237985758985528558987382953912836898684257415386114097449739437745927249233633755261186076190675955155228157598757497571538096796351333318020083285458607558829380742356226195460759706082307206702475648095751807863744263696863628687065923191783911838982001905034657752166931160914551023089972415577780137888870461202515815545738780713473139045777356709210727729288915065292497759136742380968623016123877529981458350616277854380636809475200583928128278285656046954720316947474702252930639515606787053724253393560381903051291047642656192215191684320453689044859929281329942285389171129643730055359736498459449932374538207;
R[352]<=2560'd3552133755258743967657990599909009815418084399283931847415206028293911493857005480281605188050810709147479860956688611946968873880802730525511572959780051731882170261191252447917544744726946858491021056551589145515712500469415849648204404506707905739358591634042019230040105109940678527489635432957425234698898587932290531789704786527659226231435910565698406810622481673850469825796445487320132778926030222592399411695284286870304572905368412841214706688432844746609284360386427489603223387689604721946423729658563366822474184530443161266902624950116543234903457226542128090889019337691326295479632305647679399938954134075042040662430275641842925484847759669921427797557017458265581886066228680454656016892912713516191985445837281349198447975366389736627827032903116;
R[353]<=2560'd3991086856639054551689892069072562890404150853676608834715350237876460187928713091748839426486610699227357923313795181845602609266546859954021689791375073741451458508802571549906687649203099420141461779431851416670360648781362287763209791942853925946209217513837747074675983429531511614501895605482428305461143705753167837114057510370789666237371696169106477350976291015580210962092345752202788599894283809577381053495869413434206234058381377951398292508137511845363534397160521636187897591838519602918968951269800876711309866793178606533468522030696925945175281028868134156660088254001749651409497012966792438057848624196878625813692734087536995745650352919268260631576246042647509086398263332781738788480072080124754532712347961711087481471854229174282471670135703;
R[354]<=2560'd3991093554435624772174268834097402044400750834298084221335477856287645773781682497286360707118748081758765690266778746916881785020284247994579657335826260232133788871881406891260494134018476965492923962934478283107740480207832668700476765512037504502555861568583321623121808790318655008951331828852593525172703821293548197883884546043043355962666944426873458995046078461344974359565091892560109130352921020106169806349219557695809893244217145272868499191008466869084461636355775975704566378540933337427179783630197561360764700229068883656514810431734138142287144501093700500745988618254443855859577048006988896189213519382482825573238615364661617580944434848670301207376653858976107195910283942653954285681348655770516278619595576670242440491236952033352969598269340;
R[355]<=2560'd3991093135721113904874989031694802555432236361543005264328962763681257021469890977180375116384283851084116126292781659514106758795506504167478869443854842473089950877234066495288537179719461331228343283747333193952328021111507457821555532563205013702370077048257036123169275774727313396378159593395334283140676528606971498289909908266434665588167762213804758708674002295351378975356440544635099344208776788746826283663507443249079985337900537320825544512280012977849456341008982470511245137935355184847210138590100272774553056906653446012279788013048847028987644616511214993283930691865329853946797824971189314707648718633939158806976994403237060542258256176341333114380499870043791506260463494558347061894186378991204609924051956166147784960274400730242901105626266;
R[356]<=2560'd3552032843419607264592048733527003984696903187957225618596092569868990384444659438539224198841467401255776387351755051721104938945531910162701247654605865245717774628608583244287971122699756584194134576470890709582356920874708134906117516995772110301089533568737328198178637718942389825974350825672801487887051562281075840106174488736121530435834983509282843296689989001702000145625376546149899817227854350528842827033634047432958455479418956911496798748715609484426039966817232186308459146443372707687531157964217981421942027287791979771156210228687397128615613543458023003563790983971734736411328235785147266490616057846760716249060539593880250184058945775164509731905932763850647697937195298154285211673080156561383822762090059225634875955040180566446162403749219;
R[357]<=2560'd10575282465504576609102472217361843482831562499149049785835343314671257320094710523831893176866457229421240600153374347519950230740965696050800136076542920692251924724388338129695510033453929570629616555345269981474862892215663550849420107263090452960757926948488597431195004356764271539904164541346439049037109871864004665151447905727995042028515844059101486840771572215925039919332731230468883322960180188482379401254836313122316285083380446235458763378415298200227570138906813840712917070886850691256479727812654062133120189060532396042804131242307355447112267048847446141596708767037564902777918046945781068083173027431821299178524799283592701965858723650075076430995489520607468904201385266391561422764890045822119347665671589788783820267234908191748531788482609;
R[358]<=2560'd11015950621521399553494875255119206882997895760082377196389239781316313535654072772286279616809591544096861818343335591811937295907441567545521375556271195554917874838820925322262193414246882090280019542290940644478909899884280619830470321148409008803748431364653228340272888185009025392827697118145176539792537476068842755921258009330789029408694248750780197547667802413158443311197256074239534474222553894208682294286991591498858269491557095007328996076239906520468054067411061438952055841131465888769419933563095628248560105834195302469757000658081717122076244589187841780324872216723407516407282417905575977594607170036497965229115864636967461348807854660498212753256356631104691331344792415835735258823421341593787494774121761859237105291115723919209654005346852;
R[359]<=2560'd27085252614844220819152009135992921462709273855885601210847826175405970846285970291921076609328020450685225419592886915154072447234832377475807269751335703132050180290488375032488184771013700502553179889283896041239430115154219552605134503085084901526145778550640467060564290832472820657254183077783831090796129987090407004516845172010311424283435594441237816953629552775220560375988282880727124811785801989438866369034741260990916860887765217004629663812266702925725218326623286429351321707169028747396257448554011685470796408181390385357654330043644231505986833164814501301013507410356695391447240228797172710716293941708283966642325460884806668176294199009328178204486452213245649127798402143395526585929502973944295357590555260998263295787886568881842207820499587874;
R[360]<=2560'd1696130979229865920388337671782779100982685860168081108294293922615235986252124766609714697958163293252141045976428474901926030563411376556517017771396390757760517291193169260506017052715061163708229876925871913109891963017907109008067984912977126374145665108746908789599688889339442742225441885627878838899695810859482087049499098598520092887737790486540357796375663200161298820904730673715038060052213543804276489301711889175055420767883678744616384039046487514381452782720369128428321003491432417228187324283854673646382995356435219675758282794068037236707578452201056404015533237812001946531022704206512719440612001348814810488616640185436519354995433884491716631690287113574707687615547474226607391719862352640424520594508042744634015964129168628237476356064097057;
R[361]<=2560'd1697396582020772435414631719023780925733831184081051268360904331849888164764798514516994023875423385620872113832487905633464489215469907573001047297839990127345871068751790740782631645214720227381445636190905220081736978413312994604438104583448356147133377223714071638954887635805025534314560331483686034538438038224771718037086518091559569925070721598157653421961624831193966377459846578515390329672475431982794037040574622863535824397461177098760659216189733258524111574345821364477563035375811356496855205935138962795447428548664977898110523384979220648991729602602866915017311463914483311784248423612213703995375272484356261978586764316486858466794329117862583168652622290471701819621273664435932797088531211759204223626554848051632171574663812062485097578457215490;
R[362]<=2560'd27099250696153734975544971261351739081224006951389935491667522640594009020505444347768333015185021366445626570121629606238536921520263619556489269725474568865739636303646844524812862910833152606095583152329656497821682004676628631939996215377508891892010241388691716927541176151325780272696370018105288718854566161238888331241812876664662284601494826180801470500645456436136456845754330514519299081280785904876831865941274920199442942653888740942926541256017400810241810412920088380906124688234572364149301679514197838122263617889370571965009082490043719758056225016411811321847235464432635815615434199566785625819832992683040799240912340045078060166722047665177669681786215687665721216705635809402895229939294531786441193435629073772188134341349067041240546656694378769;
R[363]<=2560'd28897229850891864504677625664416174121045756967373023518626907929436926240375470720627237812686335383666366722668238739722129762222202459002828444563112781381486465192118798575818083514396303685671779950194597586765685524086683717792825564886886000265574564091659631173756051058619405607992913462291817509683494046315052750987989948537437170840711030138774108386591498122481528976580197203145975064537694580365917330549340132510906702722434336636024633545936710494953136290354753673249630443787704176820460096718171240255821371822038183954988143555571333826334857773127981346024512062683684836262076557095943224277486078192067113902732467268309648039916783741916847061388585273390689853763673745044392131287790728462367790733440032233473766104105354529604160119665402128;
R[364]<=2560'd28785192685863981096640024393222193783890901479067945053108968737868753406465801739360140318938472068559524128108512973403807054181188370140784052425862154766170224981646832807103758064550721305448109806521994317529597815781354810675664617000553406812144860755752473555381461714828198076297526477993554888080853265451785633735260579110133668694865317989421324189412531589297775241977784594672403054887110750033816283941097387536636008590766309633678227666295371147571914950889642286427592558421880976906477577834994881870744622521329650394261248560735940745700984974739968370818691721043799865340471552647397790940018151480663157507484033802113504712518906923992847211699433132371866450990176299044605759984746865231821765388556585209556819036208031580805749469526115089;
R[365]<=2560'd122593517817379262293667314481948975122203673457545125478520527764951318122419504759913074111587743632310493257981722184687858801584659757971370083711596485579161892634544764662799472616044047034337891742305581741904512554168930685266858643522971268864252309356058228497860038225771836553955041893255392044136055239383923751503016991853015475639061276585747693827422636176883008140050368288152373571598685738224230731676840157782742063423894641258664152565867835102452745957873595995677249965100124090671595869569298581308279984110190650197524679214281872519675340133675016792712156030293370188966320605073263044494189326840098595667917803996157209631466311580519492026163291397970217955175290586613094799693603723072187286166476534079259329273545394340163951752459059;
R[366]<=2560'd1718463761589019285729091327524580892852963064205456388991918068840748961118244534278610868731934350131519342836504682111513315950961257308052527576119685100073579550034784771293202810283605544365149270200158474018158052457426252296087643249698315899811734864078380029508099610337391722426152499201626714360023432033149698019237079863928035122465741951557218853442403995055684765708171872505675878750436052789867318989773651351776101379947038255654904953703328638462162509341353122486605256660956002431239897815196836186743024107370208710207173827548763168222130098752935087527133896869112218176829280141112185597653132198195487845163170718566670272175521715494128845477476035430061707828261648991571696723873818477155783915005099907884827814799035875712735935271674436;
R[367]<=2560'd27110602279193046108731751700734888637263113953131959430871538148483242442973003303839845075855862778598180406313650679607040373545712426738293722368353382301164547341374936834598932207091712404299665987374168042191176937957988581233129770144409332909359013594879389430399956348301664645771536130170199731127898629833023045002175143017918393234250561076669939830758990627065069797909543373245157422201081011589021367066610219511673102268858789996049021951951716471065446148435728638524072914336488850387243898245110243949313731567846038312891149110399679328001005213183651481408804703061232651202194709010746570668344037000383770454390486770182586250141472994201172442372756795847370870392049405124239977437675776538592612500698865884900014233944011906066228437923734052;
R[368]<=2560'd94207886959121087612490858808409470463415229070019286885506377404589579189276117698990446946118091919106683551081599138653899664378751677461399955760454573429903431786915642470743222672141900989395004350388173430145968759475440641973486809448458232431889774731663801303322491626907871087033372854971407461344011944703823601039313664367989595332007024372255389029398432262968525624635748325508395051002166327015627495038395366791401232183874922474281471828253669058062852897691234771535060253457197969665647715609430629595499993480776127302677121558742581693665503744504310626141244759833793643935818453172121205179655787687435824156103265544208173922694292324247197119915555393397500534004289198107859871820771619332221905247573066727955;
R[369]<=2560'd5563451585595209175435383911122505377340840879980891704263285051385445040237878840918547365722310176808195909369303320235739285325123582671947654049980668718972307103695274465441780528360902633123466210737150901657679156200796948958747573141567670382746192128175966099020802640793304365646526822803090142296118922223617076332087143958122585037619015712800844632901773786894354077592017674107008225440165242641760944326955840787819798508522591056400830977908448619926103500257890317940000821831778142471218248785412380557486840775699929622114579672747202305270659976324062457604590174035757640604423429154428573020717853968208254748496715219130947309526477609308810197622191238977788690938596978950622249338207319503081365171121062827041;
R[370]<=2560'd1363860345048262215088241904927565987517441519791352188830089625535351440106251729818539483336794563664506017960506187224398933614358741730090217646793946695726161517755547449866853335010736794378881882009399394687886686478009974882680148152696471432111219745404474174390525725761118680081833816163983994324792030758681292226132684574337126125322266973211249796002732639751509738774670967162113959602467076828531105568735917519847921310503292287319453237543115557744693742047673686076276651227268719753565197052831508302470626126007843530001254935120811861244428721319530038242327861375541928434023457772673862171633745986848903922967731854737318577256299085219066788545490822745547001637916168133199862789465611458854759469877961234;
R[371]<=2560'd5349594597284138893475397197186395555973361110600450335076854512773477344679645313987519771398332244921052194331467701814153627970976630438902478140780131912142564876930163183781502326076060100834419364422159857317109320478125319429182964222731586101129291927114046549836758134299420457629018257672362209628247710745704347047102201916911202607360024943000500001216127714210025272676747469141733574589688633707073381383996516784131798886537289380496611216307069570159547562220796411152626746969955657420965413200196388519072512870193554936664531525508371469752320000146509084162671974980990986212184228709837027459799358161813046546241062346432418850578298834183125732690434762831722086341751861414830244170024115068555717037409041;
R[372]<=2560'd3961827782650652179889815946075605491022814887794528312924726310355645306566555434015034027404315357383913740762945270014543983499219206422241742974407426566418802632261314387074311549488309921985303195877718528090698343784612095161133069469634312268772733375650935399126461817696847398743668579895631440419235517341090281186938289140283827481683041001395794671262067695287389612379054589189557069800259230886241186222843457396162547295135271490456519406703500159158215012252758536713017874643922642134337413039642688054757179502442892373817515583211844318799952391261075460205807451069617025614298905265018537328603047547904131086414630075205470503317141894978643470165601955468955481224944990317179440368703116388362327573298;
R[373]<=2560'd91709760534535030514494256056830719852714058692657605663430971258296945741964085205583275306251942846787840649253468771893543538884370494485157372716096516653721929472774860499002539334227515551957087697163704973610612739509871963813161622256206675520821382439325080150684029006646743580017201922299738995369356893956934592801664859645481614000619709717687682556161187966852043626403887980804391584722836001544739044797007099225516636298188092989108365396036383320586141241340249032375446468273896449758092074154921801296470172517827369960326893593695315330143902686618540193353305608217530733033481428396090596406290208457068373826482554692502342908927972125211579513601872042645175868936779251338705343751598526371893289283;
R[374]<=2560'd40842962414425793178489861213563373199150557815541608692936472885052228388569126184507675075825549732779869605947264957489667885927482456189515787102638794543840418025588025873706627725919335038363396104988112882656168811278458550518243260996176613295164397319820317141532587058930148956546240163799853232670729919468963215646480040377811016598538374244697098309738559394194777697670199945770263320704633273465523525580166960699585047553971733532461796619480930520347123199779622896303213561709731624217427446225197822403198584267528639445724719728139510916043336707979049107551736435435592386844318478833276811229686664247082574374931025804068057201829304027005580148473443646313298465127440389289469537052631778479723553;
R[375]<=2560'd82335526130275352263614557147058148533723407360169169932865026235971525594679385954020681535080298945902562814651469200998008206536276055197043406139450075480577859793957530731363946605083756462385771589590398562613640020832159700344846926539538351415364366528728350295598219608144659746708859220800527139816371184713245698282950350190151638531011662943549267081421085857249506084600899276641741984911816922055303824999771749257663239741183134442787057676809919718849872073964015716501391140707207776976067751514798455631434060940538369872647631929889195821412361849917757714527889997720249210249749372456402346935355691196527099945994688510335144909964759757008223777585980205103417050767324888607396248719809636824598;
R[376]<=2560'd2498551612493125614601359651403483896246055022017652562287075779514148421498012378984664288631714968753668874655584918182644573339180446314776485358760457803285402363226191540673643483998395234351341754929038339409632189972104844754064084639075854983442952794566239833083015205124555592251746851218349248496221137721388155305335652467785418228801754358984614534159392655774903895683192179937177459171704782402626613423704809916143481363272393528225734654621631970451514119307462345202431968560000281531024357653086379608612530174462090918780012562478972524033247726994476107727080583576979246039231410857461530723920501469103784072096613935915369771480977686080986978271040688989122958091771745335381331125338198820;
R[377]<=2560'd82834446935425952956021935490075385003572388016321394957728654721455827533536407861031502691714001362725991976769138766795952834467334052828676647239878562170886844926974219098855024498890685380240099522576067633756318929147767976824820025814449299732139428835748490889620756031164721605980735317390369522627099010067046655143901514073693818927014938428464643225538583761920947587634323774519615601193249429217913068059542443264625159076032858942918373455002781472119670791994858586521110420640503862703901720111100413397906125252657566467424184697749664205011361625020479379063761425183924616533683487182652632386835822999578857579071653539403052599735915286999576300041395787962935285169043558548594439703577106;
R[378]<=2560'd13804617961815594851711014422846975149431661813725970009524827363918054724839657823352773314970181042135024513402737592098135298381621867629666946506351001126525955687150623805040307706666688949492988493236478211718681295687010959175775026372731854385507819029204394248453950266411529331620520580647337575107188769061653274163708707867970543797043451174100932901885817211289344003093446717176105495687909947742179366123752994032702763229069567324870868615803965858663349292943507633535900054112011585841729196284380488084915591023799427377308370584365609756005351007420047270529502544120297494221696656432632868152547500490676118702072689244857588198032155611123526970308334254634414238467051257203353188305019153;
R[379]<=2560'd306789551544134128376179870511872544839712287498930687371273659833604631214074030887140863737099472831959634831383389491244189134494729067213346909160848834228142108067419626592216768890743219558492651830642827283136940668817624077713706301971428375246785552270633250783528024567853385285198322802958526690858656876512504760333280328802063769377490674488561950919654531022180806794581977673922787430455348899035621030274069447686715358142680500276171584573733643706228921959433299522855386284066622330343402974991420671470733755925111231660433689613035616485667782941066623987809653265787931873406381981562903168500898168857656794728531854456308768601187128213448509987767784168891152504238967647240792289837073;
R[380]<=2560'd19170232540008487334980743797639608646966933268054318885744736013243385545150267180281705588529782649560046735853255911660257501531194181520520809008320504879197995657814554995477678768449510958974774462213208839418018028990696066613746231806997800535610180764434781350108036539176285058868795625191091443484633540027919985262110649178108224059761787299416339591755928355615713266173943875724328724725091783007794095620738844679097033237211277005512074996936719194047503136906471861595280308041882339545308557718471190906409218133547450017055631026668793265923729859081542057919300603984677737520342137130116269774194286490918766286018451554326306989329224438621745523805805317112856402877417041678105379340304;
R[381]<=2560'd4314298805738624375384353714984128297022971238399432523585413023510232134662943240093027401492130279932567363536682429498271044334570081340949845154143612903629045667507449211561485814058595635092332794543339805338505582803963730680125360824437819037468224392661156239412602714701348058949160998915613089634499116643974130986573201483879302144930630531381455778255731559315190809799509496861438665701972557255891109526578796302077319647120090328214718710030046652731969080932884968492687269736361177289664016320888651359024742193876607438795256597236014351309320818789957355718019449867761877308147762277386282561950409768495042031399924803438019177517129671926895209147908894389256971143167447784378571154259984;
R[382]<=2560'd3214660180265199683942863227724612352812027439309913366863429565282644614055111148738735183287824461331287101249620239899115708420123412900466975926237721776795897989672644617778005284557487697996074336652667646205785845086332243728438011416214092530227396298732343381162590504275522754915097853589546136270047570874162221445902077674629888232419179348803470141524083564527353205935120763514819212737868939604480992580165709574071926584052622068857649683760205852845663455019357745601308380381225447823143711703421718112033014462514640928446420333020688272523303375791919848164450692319973225579502139136731513084822243148137591405954115772648432134920581203018846702210098894334313379981546808705814528;
R[383]<=2560'd4806606856755855836031652021462024729766552838455343717960176765150119940817917220967891254182338477040435319325892709523289962687663981566089902704372625750864358873703607420679952687388194676380146861127304331426530584073670208508665160244761483182732950692498836253470448071414040057147947913523569236832556858852879895717845251542290066599722248691598715448460415418405765894065267057268938102032904929901364920667543436503658305962052409801449840538216049580392033143625687580837868920067867779323417407118570701992414169669492592153519616278258545829677246406367972384700349348414569576482813042533077316475213178831083824950676510004811760968926745185099853434075351539746196521516987568250132305089529796100096;
R[384]<=2560'd24630265345133851684592839489774321983011982656094776659580810676134317120630757126922464337393195083771347477871669559170065977946530026190729056053583745413337322597566514967134315451336490925012066512295580573712385970094756990757983002982131592206668138635543237685589114019073817189961247297596245511322310985361323271922712839619936854038594363490225020395533397008822907767735569011066006704709814920286665635391251075601294063069613156460021122199655597263251684712746378603476494167122472326267555417187644293048756186036899448661932471918244320169655802012659695482674829346685203089351643969443920698356634327989861039724245287717519426138990001667585783099726841965245218877141604981543964595341847837595426877036081990342155323751142576164438016;
R[385]<=2560'd279026978889740021175034252447841360769933350756339039675642147474412079941011156945839486219141801349000467911720244841805384832603022901703601097550459815023997025153712571377097684305189929517755903854717461858697578987882106734056431582840898518742276540637679531342880924969109987104107775885930621726535484166120841605256798421979955768790425111808800843281184016497399412311104056456958352706831089164093836549142473475249129843208850367368169447685182843160913039153994666853488737729091129898875851948288670712761668554450441668504108990584698350655908088730804440456051668456454749307355972001718666125899965833016912884153165282666452404660848687495740045023464013928033171249541534449664;
R[386]<=2560'd23489251465925075230210151185774156554233534484953667317186290388030343354516627258288386761202685744061840848039003501143386996222094433729614747770654120170775727249462034054381434259201992264517972882605176717825714646454999907926888695787576658860618023380054261939908734877287558893015710077458515034355865171322025601518433942722552043197182108751657368265313598727613830628199103814786643941568975440579950756786708546644649796728013552696923548922814039276875858246382129362512681913845016639199755613096464817882145581185367376268218375908000815789261853428251026622897639850369745650033331791867931409366186401276251950685650510862860790425935785654252953472163060080539949331404659226789857834271971470648292520894212682540578830965687713792;
R[387]<=2560'd1635603558075294838429993247367826069184389473256293762549991815096569328450350072700812131654348324725781875806806606016262040819261070973349527915252573930261119332768147461760123255068895278659784785525184122607848229849693896619606936637642811461773176272226182997177689158152694834959064271159807238400467575218496618487977343151339727248960700748594313190464062819022845731242210689406846397083347518918466485294807423471516168781792616454875311629669550813884623582670594809822714205143139031760911448349148290551736441927676691372442452846857587235849237516105861606836659795530445692734760467299107411041173621425494668289603880960539757266697911160099175986189795316420843427217476175974607018896649712921838003340120422585140294552182189805535232;
R[388]<=2560'd1539391584070865730287052468110895123938248916005923541223521647764652063202442912823694578702582639360052793702873417721666200745689061724075961408386008509324890582306957034595621446479549127325686859562583079616327493881997738770669671372178810540447040008018031065210498849687322326721202377254371727286163776208992933929881325607555046561280813049257375941001302303127808740571584855974865025313853908115401464356511521349287083350887654736148820978901599300253155775016700576242156525053810961848478918351684005401645570232717448041082625791356508483687833784840280107266141959711066487036973218349459476403443163828546496254126532340894401724459496500300599504514373001859960667225508235450034745588101841548980548106440404422210946897116788477132800;
R[389]<=2560'd400877108025885365940578713010340976505649656893603798842761879947784953318807136546739696439973422672254228801221841912582381771385705937706316671636594493784934245280466202412304486714616591754843792501393463336470757204638944226096112111100743226896588923819753474454666129511947096424156551994128004253024847775418830670286191612593840438967237197304467159208853712225245271021179206804218994118438582569604773745486194747932848311847275863346972657520567760205952264127554720206749096325338999611983060293335696287725162425730615490972380928375367407841047535627539751536107205657109999060269823798922446012884231956881529943225802891486549313473439710094490961528623226595708619069924954074774482653190892806419383647914949957502701782523399110656;
R[390]<=2560'd12828159211716870479923636824733980678479828995339403413231333377965392602570632879112481943558852024578335035761536534278655355822061708991314485877163540465962606460062375901904140239619639110929455472687041757876698122688104732467216790540563212432620839622645672402518116996369839237308095190164415941001630370393218148944503035083373772923200052696730224933287921000971965932646529420612885706852938045153806453124256538717667245975381221252126754569102660499530414517436453199138554809905876769582740490575018502410636488271292435704913782270454599318205557426966697653289280965889198909444885334658529713837361745173298732973831956543502739004007204792247465309603646862949671362362767623343971484831409777070694238217368460232424585056021066547200;
R[391]<=2560'd12804767449820017847632614557476467791618325434020036711819688469167638325137724914983293076976662464497311728235654519401837777034398591633013667660254350530768239919063457757671716985810800004144366327440469693539400421699665349840834639945845655196787229467239469540166162618236069012107851552331837040909772703651601340473212755083026028174045055572423361538680234456328242839963397171154483825757389625685747009086913031555478103499840020709327095396809769030257087901526025745790126479269398182208412735690022056777226370636553577929319310881775613937494068246836968062420615029333109953806004429565639077328331527756014844634560777292271848538860133494985702420073189384461574849248358922399611765654597898500128942336056294463391798157773109198848;
R[392]<=2560'd109016741454249125990573393814407413037758882684390258038289791453418680385164906408454536446923713893169002161254291717505139997631423025915763689967991506043798023588892491056936097975685243233743461009925274478744007477856735556372894547110631535701063348288845621038183598472641465736649126125566848738447588635296032006011307147858844380229676241548111360694394943965946090400212782310570218281787551445771184210196026849764441330743665064718356845309773400266205695462042638766257532720843767019038822014282080170732395782870904458068837185199611242101057991518295203915653425388669031782734364802530614883399056096078011039142116592494788374483062777103900949200926235825336273826470086505147434979868372724515535527453039458963122433169764768546816;
R[393]<=2560'd103026982330438231806869805262035003116429331390727072872701442756889362787260865072318596875531930564472179625991520834011346412588262461766095758435821258577116925479467254242424669104344709190232608948172328207804724808323501395909139482038531545558580527935415112293257856213453520487623678298174523786773991292739336917671829606693309044352854053164597458082920673557387107185164933459248998318172827136196159829637950993435742401637118836877534778640032275626503442708007360422232629469102330197378154007639095555105084995743272318621694462592931359635826332872068806782188361820132467684016730207815474885306031446189801633134988119083314342973781474362173768031418570005231906700368924095286720570416920991142404063929552284360804222813600902807552;
R[394]<=2560'd400877108025885365940578713010340976505649656893603798842761878908342338019578395599171169943001261154364073090857214126229440830838361839267171135134143895173650757410363776319085779921838852367009585124128112942077242709985907134021134956435485831233170104723064208088126563185675100825491036670264617463370543961490609241803105294061725325232438451150133444509899222492226438202127833524082552837204382296691626478935632809788448687478004996951140872641732469791281743417398165031951107874335393308654796891081825354507665290877591211394159536350417870896940692074666615544571325355457038380134247900578463917043965060279880524903601312268034948494864704093558579778573573653166516012627800145903485109628451121081519260560308829910928070006001369088;
R[395]<=2560'd889962143836803409860214085938336937524937632439794418615816774725056656318775198274332608440852525886236077086598050936074074419370044632552842147519377349269533053100930934812664946312670843904282324566598407020381678205532965132548808417147267835192084815490355307508287501585440057935185916805168009454441619698909114070436023297143264985422254325855561079772390854903858287706165823533928489790682217936796940739474496965258036967301095893871571832956893652905456563863887838579097198296702581224302945317388214298016538631746451592678548340248083588036655800874639366125404774276910344943930746518214877085763103578139280690267172695884663608029519129330281742223995305984;
R[396]<=2560'd3691999855047665944681715133635658367279348177316645925203759316108454721287977937375765065357731741479875239491876424521667663861264409663985883626442970852268330900051242641934934771527843969312262084645835916140317163241544066951092728012246497248530278496628883934217768894427354325889977499977859351643372280773110253590492807351095489506271765124000299013551660308479491114954784982318736856960234311954907601686225218716286055022515251901508054900500002436492473714851013415162611560703452554279420894110828016399940822402736691511092235537216396387883380552105355171427157311093082084052363764245668712311830686051000296459932802855337105978513939253176170486643556352;
R[397]<=2560'd1493041787808189526630419137355951764459199019333429443015935368902126370368334481384194930503113682293592218094954706463693390243200598200473840473763043808188974951247761901407991991418980598606605664084166742841020104185890570271520658114889047983179962053326186097296200548425492480945175684761678070910009508198118348716442233277303853387030339626162590007727950257717188996632396659238433879878760217779517010591564193697637704051713131663442031574496232157054070891104757114699605982816815042359826092213259135009509921239560311829880111396123519059227023370665638957144654205638995799347967820974734673546300481968343853137969457427286562316590674144413097151517862173027641673160814685086836053090878675823577629364588001736737635172352;
R[398]<=2560'd1493041787808189526630419137355951764459199019333429443015935368915420787724144570726446297527503732743316380166432582085205754088147784150913365327659140111593708659078172841215659883886774776425902668156280046165390279502624733830993464747575991993680916893739075628148551641743913689173545402257623407543481277382719120275136217429105135090642596103902953589422858561285121251586103023373844150957912563442542937598559943235513585704015517284861301646100177582165848367334059188351219388514647971174372852912785559771027588329980890647567169062752639597462057995442473121023944723496853427327682067181725313224570660581744142263006094323361921261289522934516955521537729425413093332190893499600336494986340304709969704921275519941719017652224;
R[399]<=2560'd54454047507783025985260790972171027364175609815406330882763344710881619338936320206682374542595760444940873714988481614793592072482787972865565433942356001302813512880390111042513568996730519186474195380961310303521862514361688259409650977636969818764173289242949196420071657831768923236053579460026710703151940728267153153840321984210533302680561306762446518157630928179122167976048276744492891480075407788217056300658459716534112776261687620246882677255440061647355094981939690728568233620403334332740020770641687606910190386924582657762019247954407854685698756506915234581252937107572799037195149462594327309247527318232130269439822177525847187742463025700491609126791902052483072;
R[400]<=2560'd862759507807732459914819944468806323091541822498361678160148720473875179169591372640270118711054116335522799055929933104777825257482763595817077514405379589594422965713550846949705214144378810702260907338636827241089128948007745669877946238543862482951241689687796920247775855192157142378430051597069072666111452155788404007556627219388847256847343604728702358579760346386722521406713792616645865461446781710003516847543751717113529280482966553755686205914893916696907659576289162632296825412938304628887111685466545221937366337532551369276503103593490808046200984651274273928963779428242484930952370486910640189330958783685543132334981913110424357603083197324722176;
R[401]<=2560'd50785961068496665862285318833381157918816222405146543552500652370625313065206815915662253840157389576511623787100448378497509971940721310108915728621989669538718723051922537189716677802487694600899029449677382583974142226021381988780750550098454563665663574162726827602924255946698104656117907762551978084500716674684859957290773508417988651372758850101492623825160274966459430752902559391084328214352635182316126022696712878571240325236389994369622094295164000403136312560381433180793863110172708951179494454915996914712538948479124733345794135865597278512721570559830685010972206477541257311206203418638120384171967983254747969242340659192760945091693511092207616;
R[402]<=2560'd418191306422039143057782542486874579629101109224944392151352007812340413620777106036532495766203927556898522360586624696936826454884478998599596606311774307678612981477121254878418924882689198249877580274322024215874057931606171899492640520084642508844321532916652329632419601499339464958888692720491031311234700079208321749252798802065819175604773797365483715003375697738535682461027957035233995718259409492164680850377824983660653022311768064802417194590004293495423122664250289641107686776039917800796391594621252981005042325041641528216527394950700393345093728542594935056680459702222480711474080110167917807640222709921502196640205060216204398362147694837760;
R[403]<=2560'd13888349039301993794746527822613710493286943598119521299381781665099834314419013698852104199200754388545497678739107913911793757783460774037928208893379529357130343673298337478018316395196330634375285990621893872540179646080753424106420697014672505967998641199719161067404506613838514805265506828882098251982926786072784907687995883869225995367644320430461801065548778175806665203258196856322322129545037509263481835850378351035354147091113831801786056820727015578902842036799036147250173955087157171031423909898164163052632018845418216349137502246201867548226336670202184149890108545892868535868930074743566559569992157937418724665395884703206014252001926316032;
R[404]<=2560'd13470981613970287946777546274048680870179544693219978897365995780840469016992491223689955797689402617172820017365990198222965796828149111871482919757932782227759396964227241540983889826529819125992779852457756249816831210504612148504074266679074675640940936864907615489330760398691342931746547812435160478735885381732704737443429898064793480204674316061817894132741935360776312543127632174195142977244977174035475254104887932135421474553436643666241226606388862818147174267721721430196611493417365524337815982706241800745830937563547451141679652825051230832955608431270736164871266434367344279372843823829942179482837962025520621302849631123451477753344338859523467793924096;
R[405]<=2560'd200922828540406531708023638636155799731906055247861143214265263602899144235869690960584990312468273432138450134900234478171217254505431413034431120707351984320590816323906398131522610393906461905316591332989494397988275198051106438361421969166706358456723698079677499762404833095480373839910348196528677748670096527088244531069299811296980349131070203331823853960910419647870216912915426945314471351177661518915209311044537963344103279586969647770997279133656939696043421819013999412719944282876299311230583878843066689845253596881946046695268403324513669790959108619477176932910709423527070396931520964628645205032390488224428099637862670397206074354565120;
R[406]<=2560'd802933073877986029794809829903275455291981564479579891214313998630976590205899010302523618630724225830425178299472034270304542302236196679386551079829287533633392229716598261063093274102580786585760331253599802816676486837952775814670956868644686606144208858679091508607347503306534800224763701116317416696486164088572140812417929325451196432087051376197852111353664135899245693176432557328114454972723203967683056064828698647313090815416019159965775736703906030157265327335308984653106132509301054888008472419937844482958360575366410132577013477540225190390757163136600657041951909120133817126148903810715898080221983090011510597167471571556581696881681579968036864;
R[407]<=2560'd841936350873139605322074738748897311010086061938602061180165296926450545129318685815930257953638342795963536461510736728375899923053680205862519440487072696252716854557095306970634889269169748651696245021783327097338764182959660289947072582144502056930645168847140859807282823398579376749828353658537777775163902907105070489216912972642449819044991522417158826784348654986557925903345192161052356915870852782036123901662098003037499650917604519561987321745452883545796345653148586289511329066896715107994942653996970626847728327926124923532916310199661972742930603117883933434193837089565637541463798349707964097042603712326937948737810225593230678551992211581617165041664;
R[408]<=2560'd84558727106507213883799924563964108508929340679810295926805267374410489302158343503925779238882858406087686080609727924217147394000910682969520538194262284016478194769056234162648664909647894470815951513675658958690432275784916180932736239132211311870047008630195409987625074926418772854040599512077000669117433600246928129840158824063045852965050869650091386844284063728901174729436601968403316003469623749823201527237797581419611977513588993651729144840971679653266456632900004382657758041412891385847123750891815655076030202038164434261597044950515775576661133254601423307265842485281585775702686938421842479589263675257666873110623855129939936258650552031662120863041431186683329087668817587279053776636648149277362818553741312;
R[409]<=2560'd84558797964279528688573979438436999816447336957011071081169898418083663619122001332653743163522442145546993792206617518320029541597480900435410689587019447680659428629987530202224754078110118777479660077897691847017924768310123430585604951172068304866228994074532415400654119250850254195409003123267756103500651174090183339259026797842570467700787056169759561367165550775297997916566880788447074160057317870474956172271870912039761518571430130993154947322422672832511035886694690495461692094194288154872079197392118520208456821209203469053692123259021005504390109521217350255093944388497381192810762793110205394353913882338709794165690135138261561713857127392167390106054320248551709293767000618131165724200840917317346095846653952;
R[410]<=2560'd331597771775338103801301767564449254427565619614151679007094689846189324020044666722814337666795324616983220019045094694719164781994775592256315503583526745633181435665379098409622494907072938522165138498397149606425090747165560187051286979103621599184814185527968348861897202131276138374622545516201652028148667008040546340415626799875892491049721109233788417815230167992214595186491044634554143224377301838991006384776065145522588405735641022269713734615661717907923581926539891988285812342806668421117598836388048099915404050002926949002946323081765875928222481187179360980278371103423431201415265033758032035967678716938075443673798628895899085289123807085476972208672350193729287515298072574495007830377979499574764301713408;
R[411]<=2560'd331521873910431869398966839258758146793226510980685404875941772773667879908344038505959572156456198945798954632102234114489879118747165966689797643815972108664282179362444285289514636231816012981540443815121201000006687676938459155914997657258013482368187634638593718065276531170890437854650961726294476459776696591333132732597652448454915132705025507380543310628927647392172434214724947572392356924904670916354904839200948376679668063390407826592544103779116494690442077377334039624341058117451360758399228403184788078871091533864415001638516267445827768447305243763454282143854909492330300886782743722674324947256854256393164605014137852016544089843869670460269890003760724909061453839982865665133679258383138994212888878514176;
R[412]<=2560'd47208209521469483066006922156132956292907315117999206838903648761181888818001820156124314677916569984432460551879544012439629021079282215503144657502739898986253746163250053902228920503499695699696628249984989843478709745754435933876100357742792649839108212859029389668910283012062973959022172706304904593618715774863454545635860631349448713125354066196548458701951279477164945653184254159597642533438261752842353764157185683887751927858493414345853640270344843258170417513421549152732566319754213466378549415474039602802906876335906922984764050320946460692687562061329005652981296435594312684105964695405185270597572940781229465081454002176;
R[413]<=2560'd336423515957514694676592972830334627781251583854633120954712829221390308448031326253513382987593393590096022240712920959244759783895891161329187414110195423380450735059401767125956196850645217017279813256794657185928081933778563450013353388428215165434188419214263106485067947836268797606029617765653996863205390346587332961625675055167250299097731919176887801650585186718822470268662620696765681387153888148290071537819560237016436983195711990096887521425443108723244212465156412409018840186882079244941891622751725856572872206087832792097548357687255710918053802533790885933021148355795906430001318766594910188345736834905747016237711360;
R[414]<=2560'd310877654655936111963866340110776870252988962677858841202348329047835081525773164313268852057665717712940947192670611006326723001336189939600066686090719677669203965902603179247932260641272710482112228427727299167315433150974884719941595383066936189041804202475661291518460500725929295721698917932119268595153118573351828647122506920173751974873204887777011165422598925770951702754608944685257388333765296837204656019852047541632424344821849069764967539749516947271929059568514127265136922328566199462178278553847877689143497863344775176039418981985270064975095257796833818644779056575051850512579163919623201922649918237393487647095688216747548034357731407426917659513179372504254457120526080654461673524044403907752713332457472;
R[415]<=2560'd330307508071932118961607986367700424643800772845225018777495099613324774121133987082848155299784281478585075085924414553926531319170398469407275405298939374572672560776468160776823315853077615096693925611149726744270189330970511263406050615664217677063490183384940429812731771850906183571357156405962848797971882368705732356965631484044565976936900988503117733260131967570554820867298003715835437443650112650270113067414939538152075065335839718665183326553216266362029764476180243485658644540211148748706586059770242956014978815439651070267119639722349662455029512111006564353524028792148191249759343284720599527122868262042652397679074822680701426061780471982379485080315020251495132231061528288554260139272377824610224823074816;
R[416]<=2560'd16071998050459114315688786864282501165077657772274693713005243883014820949941526882057136816027612695602869299714286425220131995398093613470582610047558877166971970174724115216551943161194663713388961942141701818079035970502906389590215771236112803323359471257512298036792448828221064860443484231929871643466455162987996672591317460568236441504257811192398269408713560942319409903353041673276579134677470651560177506670258679828954580942655293443660368166364503262353207179468709379111501486887605094548580845431721095672247168238495995825863736995864985046010256903837395276439050936635753854930309847867275735783242635091351997832348201533852612758808411630221862534818412804928470656362469788175302656;
R[417]<=2560'd16345290347096838832583423010815392501898857101168451397308824882146827428620176752916887510550373103707908740165257566824007232276896602549611278643507074655326724308017422375604081840849930875995539321857394396045229353097437551388564910264611407687062747709809964869408571233738422060967424897948566394700663000559354070591208918055116030652687936379730030478168307085058134259312502499110273610348119688235752237324991230269503015529793502003745745101659264351866980741202870160055784849235957302760299304952472154644818550839856255014346261698050076679657043121822386217585366046372042073150594683339954059853761960086228293593984176693388189055410590771575459455826153755869550701783365451776;
R[418]<=2560'd59872858414274134917887996376613159347614861176441213909556135099441307005238951653136895245318122529193843673040021706779645859137980032463698600502206997579100651506126037553191641058898011373031203514736876201842661167219402374861841124100984648647320509056851947281294314425847112505731177458639144282594812944320678997273140539963599420018586420965783424726418776333068766266033195115513595872976785129878936137115043114878035884349768599849066060142379677691675054850621857131340261114684087784754341684818519423368388297501015910640444666654864850588675435483521883240373532565295953530221594746669898742424754202310183023640088315925199266812167628027279722263000589684590778501228920832;
R[419]<=2560'd59872858414274134917887996376613159347614861176441213909556135099436430481702590687526449038116444880857168602675445754823650977185710191719441711553404402968391136716339302024343668506223304461963385430878821578168015523359758813178123531449519505113664432217341863525982853427905755573364572412007874639571709892324902514617078317344902871726710991928025533355131648115832805973682177739590241471279975318046207119841066078760976176326509178467025306400459701288786390391252439505727659446749816244255210795544715598546748868334968300951320127227295344779165720190021648033986554473269265864214967571699443818665870020073905976287357333293620289855206695166533987885058153512891247855742746624;
R[420]<=2560'd16071998050459114315688786864282501165077657772274693713005243883014820764945281141765842320406578973054717942106649910419172432595607506398836762085183809371125231235185131186073771523836770408103280109769513220420841682443278539861706656503252399016171317238555394771061876794942238691253626270886949940039921812526736934471007217960470382986877573542478557285543811259323027326727335923305508052285931047901357255543961161784689190929134100859749474621407949310349906690157032172538404910188909473449771715043378634252603047312207856771993953733351013510853098580839837505675103065245739197407973669941823345341960736154479680204310783439181219596000654247209371638450696646729321875616521062478512128;
R[421]<=2560'd16071998050459114315688786864282501165077657772274693713005243883014820764945280527435683359596305367503631343239905708448794749203169689577467684058839098951914913361799369748843055701269542261278804104765399975435546959816440386777338344233165811184874341801750146700345917759010055656649129325246771368039142483780544386092799182409392217796683793431368952724634955586833975931115347926970468683589336802251564707145267272808305241180631431567800775686370228655490024956754755575528303204675748352344447065908034970476921839269035571805614703209164897351120231130141936320985011515153452468170306706147215028372003493673598470502890700690974085374979561823130969757925403080307889883890624751770533888;
R[422]<=2560'd145542856500637466779511011192686848224711866683983984643117033499555184573191688545554602978920383508211220974875009745231956849071118134330649515759408934888172249457035630528694974670080119758381736391148421248863456243277193659294855630176902692150260362914540907867592790071239794660351664319960920925679377306754240779089574745013999058810117891316738095201216318191203923328427456729311330822961110882948811144588698751820886183648646974651148810710862366772092183506017620728780268470659697683276285502323059575828060015649197178100569414015256294642247247054754343242315738870113950325361149394554462947049101012783092203520;
R[423]<=2560'd542189430255173537666686639498907034953504264642844394716798749643052202035333585570241279680073581186260040910044056309812101596783202764054633192431838058102034393314055866459364330812662496340566600161157211410976973017594748787633044295264091979716605662684778578889747713385118631699469819744619705658602765818427511386817446375952367050616385083690861657450445690552179448278680972863413327485358022923204701620469763478253617098663724949154650005040003111492023009137266025651153293517192529133212338392487860900143338795733335620286402278094091042540178460606527278898940361281366722923808880148528477268120168300544;
R[424]<=2560'd2298095889994821023518975698609509503666522255464822801260920562110446064383806023305340954630224186704253909881889299075023958284747055175681640271379098919349929483382133423160723206024177040682559573563893724631447200751510276164132325723740011858260858783137818445005686564709561775676331911933143619952339309902600784323597363866075604514180919876303522667837808205591680091305423370609248920457009428052676805890020959943720740595674207556747314269498012412629565742859235243473664491881886229020004270563585039592792658822429367381430624914491320523109469081149359993117306015469910483780386207429493981708288;
R[425]<=2560'd135182367475692618321699195834733942352959747211207853694184203089600239935124591976640809728319968141196742232337766456230489186840698351583826057770218625633651201632551660194624638498257128270566283699359307953130802273151298081143946327738142564460038456570466829514017085188941248197821592256217470194764011244020200029437904101202020794782479055444256881305470917693783460741296225006183499039088266234776949326971402910237406628457168064306737796094644518006226285996610891207009226398921163992050486228349947254742222027402655462521759648217817288646922906304424103212577978809276313949659356675291087896576;
R[426]<=2560'd792410683174719618142403921016562069266002468049343401034418902823387987167004328920977190408554508563198793968545959099855777589639191708059158262344484735000249456609466385828133250581140515440190962228310087932612688501859038552843397147551670156386803987248857059541509165621632133849287375055469161315861468051164295180883135375448301335191110883514132997832910059538697916933913708676139302547177374850941012286444521919557900887550520161419887645778451533284046320485224609037337853209297860723744980286671651893803628308441664659199123807527390992501552316600242445959612154726747709449118290008613457285598031211122596043262305367473772230220517151694959706898432;
R[427]<=2560'd13470981613970233508420866657281555177522041956838837817585120754073501529818791348098189281650840292950418274060416403775919222499242430312238916909483172738930411128726891369873047926967142215942691465412841089456815099070077286837564939435662315223778821604021767908735666344470513094597255279340926332162287956470967326953058284800357632132017748832670175981930096414494537640368158348718725131635672448340516000027061360799980250157723420059445878984296923377306806513978095397033923789310451178992851798046820661253201334887294475580440346820639609714982565426978645416973112264439737892487107033728917805441989700371936185814186195968554745192778068677726368329367552;
R[428]<=2560'd269643382844131460043002966000030207080283123902662509776847888948396696354802652541803917760512822515226341965591835322086722575665868969906939372041570233681998804225943775057706310253806585715823463928567469266300837170341847539771855666579081377453006875519145811545731332485700951557919226009537560955372538085968683335378130455113847080547028931827079520196405424605765532799351246840402296810067289688822231475916491933606831174386651650195008512242656555208322260565906573525784575883390792509905831528107290509257037750410610854824409178657047694880416967666337737719340958079577852090058020710618659820029106775028132462032300954075641673100056384026455897660054847359363754761540021836711838921785344;
R[429]<=2560'd269643382844131460043002966000030207080283330209231138754104428175186588095072227297161447849651313570095332160372751562941020078143663646028273248144057947910346470742965251520584908226802695471887817063040393183802577542699764562870689156292541126021848630712100264416777569895846095797756925564761807781503869334414598641358181059093949248569667522172956679396243493357557546215773416179671123774644634935560813151122947972507567662226370815280435513868657345994233139597394808599480626457194239991522482685355018262316518053862752282640637760627469470817640248133475605213382774881129894089935293747777225368266040157230143055142915210064898526749253648270700762083368934449001852512012394929027331498442752;
R[430]<=2560'd287549388736124564811483631710969713018310329665215642316088126448179996087146943673301862095333745446546114612296804948281926091530992900564944573243546318658635876471944444183951485043709821750916568995831055483387766408933386434394080415486861557470507978663924631765324367176372312458320445058312901664185474867648684638304452425271159384890036541267785509722341247488039447474322218525725419669539175846841315716083499177506780529595436226647805335923985760071476443660272563059701312856054638673485049511560884405876644925814159776689339331743663297885680141632251419604216098396624831166214096459774074539032521427761851108198029560809433513573277797160600744767055307280741276798445647045446039890821120;
R[431]<=2560'd845238058904277106894979680903215812043988261786891851059284605293500833442464071419492430486060081575812714298691219121994109708623891866335028618582642643291843496781449798896824425410914251584485542597863047106432436613061362537803329320647200698919890385096038783805497470532319132803385806093893150114794704312209912919587775111322505842547963065275235787987029637439812511582062217748710802224810924311118937732468799283934721387941727835116592576772247427743205964912200698511368351282967505586019850295398921195767637306768880882163025620422143884421159678556443505430573219863563682699095235710232248393277055179026422322339501991038605902190558818692015214034944;
R[432]<=2560'd14811500922130502915847482749949290231794744616576855868049323002173864180226355985930687664885644589159528574400112275443094521205481237006393782470350018009214302243023691257460706076205933516236253553322936977327539905433957053904278728074551055137429672785242192322104810418163353839208303047340138546785994957040314879114051014115621075665099557316093427017774855694612814336488496091598104302945106484341362112366937922781372503703488597144412072502072676696557769155036629735849444226314646502952133842057479156695842249184805122698772473365033651769856163826645097339715742039124891737287097732597826081220722934866862935839148656686590428944124457741359800179724080623795568640;
R[433]<=2560'd13523808992836248317003575416723618493616963940239526826442972261613706096872451237251463753410753074703569888073901347384156198374218970109298669354006957698634119150014301098479482392107707330131062058531815857535057347723364682332251461031408109109895566911913669414083730986086595894489857004242213207263764587634958587537040118118778895075135414319681026172439282564477321626644963694051421842284857924308033545511655874589673303090156914215795430135607460310038501456205168697415422922456917132100142166584701656444396174147999054166191351241774910196875294685533396173237362746360784225398649303564358334988683499989586371047190018926309371833045928130858860542951424;
R[434]<=2560'd845238062052265519812723463545226155851060246264970426652685766350856631054527746102095360824341926389297223771870273459989375984412795246065280717852687321417117059782204304802513656124910527798388225993850804838511065405445058974535924700195572371219631870938385074221679474214818157684388687725605645471890247595171659563629517020226065515155662729123060197530528977397865242234440526752375265343466254359377627929315903825355085143355299254621319395415437942715351399968741829992937676922898474858277208152143191101334627863508036096329676770158939787477690955106937621734955184282450719443740728241077496410262784153061317401818751988249615461924984583040953739116544;
R[435]<=2560'd3148709106235719456584922891962705471654012201640927122861627170309996890353343090866778271942482053757967208956365808865024130678500485192746342902231511644035496747853738914027925953917060645516218783725305022444119990064358149519039996750280710646867070748183887501171850639793294340488552633023766395499171962663142995524275704071478674925124206857776635769922273497008177434898928752015743152729513841535631272548560241970016610228553698918980370016649148998480458457860490901316308269024476615849140066367959431571458671432797266805162278207023172697336584749176812541378790130958077312084079378613765530451322590217109774101554217957403736004462150066110464;
R[436]<=2560'd3148709106235719456584922891962705471654012201640927122861627170309996890346380038953307812758021087509528483335326729113042308413305887686824836021451658213002559886519874514875897706164905821897239749917560317859655554169639291964610525396054101617735068629956822093071797162978414851141052394412750453278041796877966521506690128493344799165693303935790162692483682858025008543458146494586854299608728879685077023190363353589875490830419416839546969369580054326058342505178285642787409547517758562369020149907244955376696743220437941095075349355418903533410511743279908127276055326048468703346527557897921081047538588167780968986888074524197237941097115345223680;
R[437]<=2560'd14811500922116979106857795255782587865282111016134933694843642746086981352182119752018729370255528157829775705314366535878601279590024121230826133401780304939805510706610007970683113629837000680225970245951769534309369604343434247092782571872018579447588497492920033123655326516417826033842877029320750365005660131047470180826467823480933440595832699850393385777781753174541486184063160006616644860085275619007768353205752806056777076021362184792220066777414300926712643237721374995432495790984799119406984335681178524264210634875995120155707787091958501854527796377086488002874747341885533731582121221002649479965764449248513765654321926065494829467072891822614475213511933798513639424;
R[438]<=2560'd3148756965509482246566357553836023677868551730286892365665770119963860527571112951569419897661169166596714319126496440173528437272906176281899476042367689196519579112872419531838897858037146165091865732047714400030088461275394216281887402237449102228469612174424407713251165381133503952060292452309342396530114447718044479107135105338446267002213201134108746112363232395561351856820707742260355796083611090076797039536835089688856499042989260107125922132075421577181115106732494845252656199392534787799688508821876291002056792980336353060101010342210503807365982784782683048748905209699103260468075973393364606767051290220231390642079732022010209364924373143650304;
R[439]<=2560'd196797135081121776396560308361260205244419439620552815370227687006829426090551116870897779926909895076934756412239176000716318188533719925614687090983289874189395896752859828800020735334962979557569452569014352411598495059485856213215877463047607579221789691569813512083248567856854522655384565241157676559331587204779769372499535206894584966421213936008406508014068961536058209375130908855752770290497316866672148643536798187134692195351424510382129723409675051144595402771714717676799728265626643939496432667126151346586751070393567245426513209243362429708818279556737305927132203636133028946015562796282998795845004586735941202246351887316737651545730755592192;
R[440]<=2560'd54454047507783011422259729797097033270194882714617155610913379283177909869002360116005362771992929250036090431105125287666753933946809449647894872753471683791623621027906278272440682525714654385429321432918167307422162324203753898853618032961672820064268470706113069281216850782456711487388430585837422018336114766407637604822872864808259576986182424698010513717822800035155363967234739079916366634541408864227279482077839560903302889346339938160778487158024643387788351536877604146299753770257160822721802708690725878948104067471343308994998378400966867309880560562503820866724291383895643422968973614703715724507502370435880385720144998774541937918228583328873394222413629716692992;
R[441]<=2560'd730263376568940700859625258789615749768712687965711991346677261175811729158954226168239895881274863774638020774561234630385542615154831147760018432740970275360326733515286120856698198619252633784829269122475159130506419178563416225917993890243057486367603571158105228807768895904065573675523887786808417700400229383236545702859655869682524395613164460274019422080079820682596313914915041098487506008998595051847697009534161306452021141827009977360652246848687829960175596834285381509635927511458608802770781426697988680813067082700451379013832071312691587806196223245771540459033119989825407794997750399254307497362163130921092044267143020862713484017664;
R[442]<=2560'd45809260524660112898593220507712568861870074405937356074826032238280469223436234072531722698406858741051918717045216060025340105887264435852193487873932951820849591688736750924252191645112849916267249315786691880602728258604338016909905550478741916461545386250246482640652132968716526189915061786668090522289093898146626212190225397059519936489255415853225660231195241305992741306248078362897260838988721406326803013177723093518747483404548158540616247810047170377718186795235474645237424874796083899946834421203367379039596915258805244955175683574364274217623018126463808377962248015036486468342383709378293265259365178749893819636448969901976101847040;
R[443]<=2560'd45809263085077121890888979581226871864563270901472757691595680351228265749225082063741073629744023580395871775550268981650993336254378003354241978691654443304624138883951824625483812313093294151568514309073135610387369281467670219283971098533696511311913465128346015752536983147859868764564148473406247759143544149090356823164196443128253877524095539617989281492753957121118435000502787897024779315543341714571401309387751478155307331216837112692739382899041050818105395101639834791345594648199340853767392188962853717035357598481537850174037088668130472728356110489930623215564747763119741027740811314548671763988511836881406603104592153827286167060480;
R[444]<=2560'd45809263085077121890888979581226871864563270901472757691595680357754639375096570542457361198040451633845090036594938142707926810475817488830501551293462029389434936286190828425014525948855819981737756187648050237097694952137612797439083029020667539179044726243193455026616662219448007340467466683954252654617252167239135170161074106442516195538302511626281959766971403476094192543250137641771478502237468650925245365028216294830671056011080702485074010642113381340680674032334830981647410911808791908829259617623279603373135779915204249412487198032439138435103691826154960580292540623373606367497999673031049299645613372768311937565867203529513478651904;
R[445]<=2560'd733115970444080134464653929030276989293939918398613455429644867339819748097647530281667495186866876517085167224342681094375006218187326521271771833955869193399902567587186311072706857764636638210200677115278341502068287832819503634309135838262319247390497755952754701145765196066744463730167738091948182616336894037010504117775536921198722727619110460672515519049452856220145745349720930459535464771857616208755486407426535190824639636623303610023546256693212395397652940053152558186293961004946592614993223661021325213932620821958556442500598270697742370156723352927844494094131983785805076177426840654860963926507632451512009468237279912840224330219520;
R[446]<=2560'd733127110818486259943501657891009354012037870473145889994383805000918290657889725360900188829268286001019690770150791938514331628740252630516050527976230451370889760142951602695896763602923750503015238390782061719771302782712388600426974877699841001209901578533081110389226990855996971710983706674099422864269069763860008422181604048562013769533011301930695379882793735293077183219537955887290840749315119557381907022241762487399238044303993249795893747956784919028618771894963525658815798410680357467717562591126369285339649687398244781527616470316138313521224234528341679778623481728455954871150807545912766796732195919883095260577101666507601355997184;
R[447]<=2560'd54454047507783011422259729786143093150095513178042938039359956983721643539158251693961996465407827650893396553715278557315235857398858263772153808847941932164807140347402738301989141812200293693241669450028441499794938129871519697425601545278958371531493126100416129330686152760136580920251565403182738590120386677828373408546424241340860886020284409803429415745894552840678700983038836121803392267491106840247476339952691974012169976599784862661302039530543376826243465613652864757311780759354121689770626169902136195116151974643648707423030833687148529349592661085475097867498540265924646644270874966618621370910101929478495622794787758573179033943628374829849418803432839127760896;
R[448]<=2560'd6613030781228709494345677548871862230391902859855834286189875385946889970147418863843378937639127808320203918191267461212734660798972334263574329132439242458557321985092634264192249172378434196639715274698269277854234574133727049888866744375449994196704090442916061743414279016760767639908978961737481326435522560678761227776614366352108848964613002883370448598529478436466239018254640083276022201769876210222880721911618790379501668600570368676068409539558002257905640313715245227741590638214347747779976947064752649116892277537434578427726868253377283024616785456634033647606824960;
R[449]<=2560'd3742053650892133432367999773538322459225928823527575869347258443714776254479140165467924450143929014376701328044210206508077474988048249115724382795449561804101395202715992313387002230914292414059919513091074291001085655127805431501636336560296045569746324243978906254446466591849730349755870956762936177892782851939643713181740966787046383467430613283629097749174178949040940972825632789533260831929958383570589789904893954262698957215539182337793190391741090833398321104932837941439383124864410410169059865552096602981336053283190008904738843449629376937574265244739303342293716693242787314983121133868443337025544869584683842845704958839918288197694183624029882344176950644163128895865880576;
R[450]<=2560'd63614912065166268350255996150151481806840789999968789778903393543151196326145382812954715652446793244403922576744547165432261570959077952571638153982433111289420534943709725973530190478632002348363667765628640519045622188548733550467879397419270917704869042279905901497514177990680038142438357617337825038059022165288544133831191571040662143605103607622073471930237432906188686528532652635376502133718381446644727642616911834846640083471404715357699185518184895695169730852456060740262213354288703994740980366281772884771041343431643898979817989455582673551300690651390214467256515866789884599870046539273261241666652112102117637283520267890012514113754397755242168196244403003542176238139342848;
R[451]<=2560'd20457887961217337850711660704216106603052382081189284396601488260045146429118212912885467223834120398278215254834494797878096153042887635028461531582375768235145639305911252688342071658403807887864460823865411988760323089076260661199054717223543417949865103470034786887653762198635835677854647570532545651722355004533373752959608405315144793750248255861290040655857452661670504719406408628512230906810771210419725412796816579695424767133605630967580667887303060649470069817518394244695633760844047127831435817281359916125720906586493578435155214729216;
R[452]<=2560'd5237139422742051275910067458563335677476390497642818255658004925335665628343701443101850267757763208003488906016656851207957351656083537981232274796287226688644920531267598182178853338997359545296310920265094654649833710421359191951343567903744436229332548880177747842486083576618505431030836708604923242698658960306178629654578754968424101961188604194627382498277180632776202857356547201573318305034671885219769939003875370099402213834348218326234971600030181838130790800007987849114825472964479550286473906940374225301134698173133062583821548585484288;
R[453]<=2560'd5216761448334513262235020346059532842953857036693831205524260891982235708253796029917131147504958483837639445957739536261910902336491977752584629942583919580782420142466788902460823397436657399954371592590300465083947279102379702362060990670002460583038443839035913057287457313757631196311001126112267844073065954881194546357058028711262818899518847523958911566563201580163467480419324753689252601819321006458995052945814473170221082364693783027833926008435461719299681459485641530102318830755841575872063155342675833891408287281757020986573133984038912;
R[454]<=2560'd5398484928428591658019859315901837254618609460557424960467397595046241867785799819536236261791255857160682828825132898019097135628719052624908726699150013771315308705254311093661850922121851123725498404611126069617840386482507754816797494876919632356427745061425565758646124548671477452321278862327560523404452788008025977509203457669108034616296976370068951527211100740003651069173991535648229865337948932657183670902573147483919328652386308875271194386945472031734122083819108400229912585720301554190645419736908403731720845132237547998731363836189593440446578688;
R[455]<=2560'd1519538322892631660972446247418949219296324005660624011595222751201040299131284998613764783832311835811999056684859548384956917558180437956864974463709618965461634658861980317112507147254549864374039163530415261674945667518581402894270108644200067468890728103521908246228279066125851830914483933740306494475993677541626231874788776218921387681002544624195771852882182800933841321029244363237022221245935281789525239476747159167314675535749548420193024960067143414092081706653914066406732881759537968025847962808305794624779588126810668834771327495557348248582291300001807794700288;
R[456]<=2560'd5660807748171842889009917883595394469475052619920480256643646453270818409482158895416280567894408857367596058491783797983844982474676383739238657903329025183868226914645658194951307391548130659026099072512557787083557891156602318211275084377723144683922830171766050915247007733710267800324575872075878754322866446652638550264105884047004347919772489998410199527645356931176221833249657641478650058701328979042683180822610328327848812407694795436119432985926452630212480064293949232598460562040392617062227834803941387206382992302966499906565623879124525446343456347652096;
R[457]<=2560'd5490282102021674462536968404635136178847218716396725159413405606031980972945914678736740169760034912030830659299187467384220946240814570715391257490816324287608305937025179421088364635214578296428037761966142146143073735204106320559737588779061850394222976611973857961752115422857106061546141221704415068022311392212012582424011107790576877171450008099281930411781277418460306188702997392994166403526587343394494528844531030463504442031938352453641324069947746706459346207782334520956241397098426178335658237397905081340382679588747039531102501425272911298560;
R[458]<=2560'd2250297766757528060363378293585466094909643757097628584211675966172632078907267056294086240674665098970649373303513462755685013357007775537918393306611932825408415628470160305351803125831300962704603533713495202526872855605106208030681511048955926840676736176545671896108157136372877329031250631075239401076619354906914337843634079002429616026912533061368350411797158040366140162477045348324533244592219306643816665325778936019821221051122011380319768027747496477190900088338993274945612594431847987885120756999385317254336771073608852169406984015919770661094668954916388769339961131540354022900891779849203318125141950464;
R[459]<=2560'd38255062034877977026177430990952923613463943876989646440678099775994602510038551423119701779575718676984194365267817533231549432406789619084650439829914154418713400444724739365331524259382491775918665237315064254109312406660655299032966018720680329248427685900396388997026733809617123856947905221947181276808947331306338526751243739140965932059961702094349265754481316214940765147301843203330178256584602295420210816539586041976615346818006031354450972888879652532529996288959933067391119494710394486956753332543854836832638533117484583340186988903897721340107336921758517010309501944496897188683752808854560907752430895104;
R[460]<=2560'd578194155599816621627484493316547994268548466535886801176320088913447313106701098213049063879180391798402051474652513085989015020705677592789148856756327054470737723348809567937812926546815316185587961904667592583608689740667260304054630754335686386736081823942911032109910206852139738960650753394623378324808600484502488015895437664788908203684980568105243887923890418114632410152978585623156162825315256450325623104488023230167779089805249812089557498919393664942994641327640278121381573442343398027983207981344502842639834776033688365284474122768354816888916412097899281211652931155056804375145486278614167519469733150720;
R[461]<=2560'd17892249913945973697835124540432957712749807493348620904754986542039218993891706609560285426472804379965466008021994293174202941615430272135291187402319850069655139320871501257572324637687591284113044777748162693504483476077720032294002383164913104444002110515540030781087076557176158583325438210528444172106844431720395360109638612474623555729459854848788837252018018100061281023378716907909091717425697387304828755326728416684675605852704428203494889965224677210388369505122202034206744475963664444534881851550403341878981721253189082045628407263026993316172811172319494453604631096388010351481352573838490384612892170256384;
R[462]<=2560'd156692734094860193899222757338943175120748314120155527613847053562246184551250611169549460061154468721401509664083974031162840689360289044304193143953849793477964812166946265323158620707921666761939354103983836313814480250733172709496247687761281139165835891455481906688131749916275057612042452466976390699197810546547891694736316711534726912235137481831300730920962225446950878735036357129878551472595263453021061026668532209781692593358490611580222001201185321325021217550427808815144318208560368202029632107220880543637177616657404417235384696070951962281879358936168732777346075626845475257253011596683019676844306677628928;
R[463]<=2560'd60667907776991146471202347000463109132192141788440003476571522293024134674821788543153332786714036411597384955107640624667015965497163518457753120166687084966038891051036030899525518925008266059648539075454935686599784276954881293741098629449712440606109117237868112921716547602933654239733337464411436182741283062860674452579045255278728084468649995446826734620340834657252203304599971784893025529029566865432481841898107217155813049042396272662342574995515405286127559271476642985512589485940586399609544804393683315937101521346965113018688554648404667332415268500360033998370981592069995234784397718881892862317494281257301175934944308155564892071439317553814412331582345941940272365568;
R[464]<=2560'd24630265345133851684592839489774321983011982656112682665468339468736876812293776615626336789837756771381025545554249238817396088481162607203904074540374710073187058030365424918776072078960827719730111103066613019197237055434859360553938933599812973275675194277508905792302237133514130005620068615063513743242625082776242047098868497762964845721084061956342699458428489195231726181927950808839655440687527847444944435084549397079421367059992050711959963668029887855660723824271575163886775884396181173354924770079581644152060909518402816675368971414843847200141886745871426022597767704252359846713797350933562741702378688913474523239589281745969072329504704821151767510049944404519843506435439266284176401187533772715342591808077507142339005182594886308724736;
R[465]<=2560'd1715054636911677635422294878265538158479251037731161574604089646357207061648773964739148946377290719056712207783378194615087604282713267166306510433937976679728933964081744934245786436302452855399267922755402903509021479320002053230906432788496913884452536643081508813220089208832929207185119145772670991066577295069252236224846353071219263697892661391303924579547270048003276510222067136063783205666736062510859104071438372273986590905084263392618387288025493973988087922676971162274458519687246574744613022301430884707806780592745698472137708387031969021062232140515302738256580057475272650285803145943081308726820846868635127252255490298570420416699983602736041145438654898944252877191698187220821285149137534237677319518561341313182589896842816340923420508160;
R[466]<=2560'd6437614734768992877050454372098012541450403863866512650673381132833836909457710653322613378993222334465712912365466799916740955700903491030805658781416604528758135584696801772397016732875570804966201064936314343498618605615823955162552917128122509172483867787234332892294528956917968342440134036047555551875643096825340721698373233350735690569465173368363444510743648483807714358229529591013234325769256955136139937390835380075062394883213752700205571863459328537400660072388661241287979538167202502253891769134154486337948788438490454927118435073347517425556159387237854165943943584257776067359600108290686064107382871065599524528943089971144684396923326144140828153628555737670344479944974455702991219775195882392864345077785461833285621484137111093248;
R[467]<=2560'd6414034110726200009033546941810886386503025053126107906715922020755233929037325479446792272561786227410607590692534063418427631467251867074652040237666576814569932094398112335004343581006768566745830930315030583054887973788485239888976939000657692430289478623605239757295111174100908735433944002302293880570511069577237083529830457103943351556094438316863156455067219421567228713988335319848189767166649863439483498105136083108411887273869651738450293734833846069521029942046778775480265369584901901925897087846259965644765076804737272444422799096115682195261174671014092424259237369285567342119434210466523015486304295415229178656024736616039051176167462601771298431388253131035735674526119389735446371907416429564166359207847394609814372716841097232384;
R[468]<=2560'd6116899231352010588692912491002517341701099968160183252840080180177279449304537884595888951017519723646296354700704913414084395890029279507549927613850179013232576632648908906998869401600065813521492912413895295269913092727682544552863974753057284840451419829278963747589457155721839283898756522407557331196429983396511036164907962668438981329680838126433939947137004054299425546383690506800483309481694913748680000257544476650119304716924293921065040968801108820345228473270722031583437665467040789389720986408229978270343758293839956545331578777228912443949036512109092911518616962456932498232133954354488397388165144419112648965942153369006645857708184891332534114342716178547260628090587074352404137636995961414971441583222632960859507697647616;
R[469]<=2560'd24630290400333921931617441007146556724093598996443819707875036586452786944245089467559389312042984220644044664278154460785157655936202529997837358099552723706667216399826050990129857442895023165563629998371285947587932997544452787518471491450571071646732560609889777508141004543032422877358859967176415205670768369549574745546759910442249861797389816987940576082481623383700931805563689991645705249082432531924346346911923201555974196640867190386597079705271790245433942868552829517181735195372102627984918489897392234868786118493977311989213447243371722434491695121789177305332708722824255612531894163818807150535710299516893950958192410888893053893006988635057529363590466045099033644807953335106811245185514063637901684706954475762059942894789406935220224;
R[470]<=2560'd6725704456905100107436900048333174295956510044095245913092935644490609821169984166730443696721226607314087231341373825808163820981348237059640632169127380006585638223782849229547380632617666341091297725076324192180052336512473551727834603751385132263963903830927989680207445848450350481085788942349654412957584513067072602493314876576519717483175538419370688723570464671163377520069712141440789454535441605642907366891232111629722049754136025920923623039896843156546804519556214811202853774952204499044338488344041904874894309714977962044832070254821684730526042111381258811994215263807617649748931421511793599945805421065194471812682152282803657868640255255048313793542600949505342901734989777517449547047673999563826963452960140237243510624209408143636037632;
R[471]<=2560'd440775767288133425994122028163678371364413113796015048124354045077851382237722743186369036681088688340366260901455331400850778455819776507138528380803825553741459834298741631413872845597456129419568202523364049556906705431596386572475208895603729247323028325507855042048390460261992831662491892015942478012714006083923072668711414492951424761946911657049320727744825805003683990200509123636364314438524875472297113618101999280794051147647392168650640564197002245630790573134205710505464650598173737929150741689414668458869204246458743227704812990451218979426807447021059649361016875786945845043321459351185388692484143766403995220212235739955562980465264384363411338075036348057692920582515313157986089411775875023493207364226509239520813317203414505646824538243072;
R[472]<=2560'd1918256132487621974193347895151314843459405821322660565899360273056784924517511088016561893061021147572716138203353921277904629118532150107389287887027297523088344172692926464883900265426508337945714580423564174061471447844190756904388541075193532632683029700448582628715493699051368240506317064656454454350442590178225433687267033162458867969160774279165254602886044336158483431400162907587820894621706663014942150394744042181029264407019298386670032057593326187897854244832760115836963258610666964704805549506477670881547210008737217161778491380041625789855988605143895785473159356288947371824546164985284153613131548979340230941700457764762602469670905361652887083864260013117466970378721807205720625742396402500058442635535533335106998825172390103619284110996930560;
R[473]<=2560'd59571724885910220160013548916082617318737527699823358414219598071889496175694824584486939478462670779234645508087110321805507538873878766369989439569198156512526757456959807955997459484895445504016006057667148534895339505038231842007500862490508206355685973976085634445805990383526156961070298230349612156211291431170248355649325163574410033298336524897161135897859679336171127365160357877920948925605452243787899907579682019343769457692910941027262803471478153510079070490958451451810618912328753824349501502785432142968313266861175725355887455764108145755137998111381239587760893344452642660621406241964796402411381312418525961459636414924173336451950052097016814377254845012779171347691077791994868095499901032289648187793365596227668689115942431569017638426691764224;
R[474]<=2560'd59459328672721287006973309852862471023149810363886454379565684593635507698543432729841994612555561869509104972700598772578688470190405595195284230533708124695341403555769418183450005993743298969360093301896839802070376769147870507781459049902910988753223466901112219454381416911382111763456480434685321957262736505989535384726812653290136372377438075192795541919774519653629979250746805543873040994112673662315696524567290397553956874809729787974649214418827847638305228768254416986930608770050708587037651744516085352740576151508477603754554096696841090237534664700673097567199276533123929856943991841367598401925372726369652013028968248646479477379818534486963058866040822693118696320339858813779511153211358652903636105275254279221380822597319209722165983723007246336;
R[475]<=2560'd59465940316376669995299468068298596700190956245367989826207244611483704768514375491316762861887787918220560611252636690886127377334695404629887871741498007373453442570544406768228742823682652491534178129580193400804038525294315410856829095487140970205845265790640969865902642598025174019397062724492415442192708673837771232843888907692185775669429371105832481330424332491164642761196124107800337008944026662517757261064222612163151871928421541057527111858039791083115039531569372149768072438027901071395823116123897587973488659506198636344837800228688434860226762104312480244814767239536128041381746386801273348330427323509893363879862072845196676502657182176821335096505305855358655409032504892278465415181374157029762473395175718184050202306964629786841874415273115648;
R[476]<=2560'd59465940316797026500361049184805033395877581029460197483811053876762743697326421862718406040384442648857655488147782153934191911742901737272612351006608976684302730525163421680789441596328505296464883432826534058029218156791449981837642933205120399379822286275220301859034879673872352103513238572524000455497477499511935276792833138718125334840759954189731141886847952980846992181346698992880278118503468223496804008562770620948053335371612175271039007648777210257330798735497010115618128632093309561136045544027922645221930107327099870641827728492792052948782650043506677191703403640924374476578149654431451575868628617306434232727556228830709403211518901921074918869885699893239616168485519042917789647817562270360791842841220691157163188164145100803657692521741418496;
R[477]<=2560'd7052513162176988490277952070353265252879260512207169097889679421607081811548535214358234060440298694150441374056364309242659718578059297926831136661898702340503093247917063057007253787460953830734586994406687748883831798322389646048995762832787905149008883978423527681301208688713540488763977535954422819614350003811266875075459771159949390147757124512468053971620755509570541148566092611319664299004061614510417293054545336017363728907508982136914052850521075159872977182577879409221794942026636470755029472765009959160145883305982750330134597845193913047515706975869333491425618464414039110605706107411380664763400731513416133209147702573469691881352088728595171408655281494885773408625431436940950739850888558530445955584620811078778994880208253671236137501336080;
R[478]<=2560'd27548459183624633824190032542395180272364721256983231403337180728595118654465986728926427866374383047584223445444697526888289541200313659799140353096725545957508657394722554852030326003058108124151706077272870734204812426356344387624135459026824924105593909747830087190433896550555756788255105245231187149641896999948274677982054736148912810132572970107513539197697589332897203298209708085905168132619833985093111767383935817063382088710711140096121082612332345138657777101848701735806258987368881778193097075107710598038169993850003202198206136038344665885082079229972231943731631291929808606286515315373926298629205260088971939697517643294066229259125177843641576234421829754885446669287186126175465119490988995000254827450774799424989706676880669931122418857011;
R[479]<=2560'd59571285724758533885579757649699876520710639178279911664822497227327025832116481664776412656440048766755748121333071609499013298611007842233260442066271742993528641451653458582339006193868318219393197362052252481366887087652043593076861487645186316323342142320278552204881183175945402841703826313078600041816934660313014947711579911029986736156276993243839835392731556029354372089127681575112036292983651807390292637006218260502708856995517606484115189811681524123968782578934146940402755873161584812836870455563936848547240621377041383844580579904085078210227099438544085092599728038695687567486590054190256177932086705189855277451857295521170889896128984040558614248553146847896892100870022554539898284366930246943889666324145842127047839390112636972241283693796135168;
G[0]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496925171969057735033576824097598527785085168107277894831459066049712703896700389723584085603123985382312747032700348759204055392658519515229479066063683907478940621675446335499808634277658221467868366515898746321489526821436448892255234809771423692784338485709772541257076253027811387434301350638550706041630006625795290237392112172169576127108230397325819288199629445391225648884147093433265605986003367626965419536710250218152876774111707016774453848881614230668348562743377910263259548821187040338890302397901142705369758211051793;
G[1]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495885461657362351616942036405055437279889255336241864930055677314763570635458205460184561168312520156065598085578249936891055439719644307377843714653052538577238992161495635718356023918652072140449425214836217326681169233260179695441785720782357967849083623124172994134169194449004694799156564575237554956710998632650193559704098691081187344565085469517502692623892716423545311837400316086299168328558858480524127677460733402436907697755660067445968265274833241942808996787320990971207470182632938529830568454848362249792833255969041;
G[2]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495820479762882398559865912591538877406035824982230441511140989020827003877267741823680994220707377504979258509145243480211848514957438343362174504069686286684287087628569789063096980278065220625429911958738540217069392911932024032125534843934686796045393786140092152894097634177089132858878168719236652613450328411617905812052451970550171320323050384150441000198291779612154739007152919791708171024672790767976023290138649831773079193021441232896799127071525401227622309808810175823632077653727579802877913693746488661453081647583505;
G[3]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256726886656705387690838569640404804394626512985613087085960452164785960795291266319037962900116132588746050923464576825700744542036273482094243137271001010089245241820453418220997674569053607256181953753285570649572828097942504885970199450666676683975310783238291934575770465838185639335359281671756863032553981619559000483819473308010066557841226250002629058919028782902281420294913984258058312856291270601534375372507601463919685131983536837093847640709794298025258153684301057787653311033492737303665729225868530351418688409183162564787376401;
G[4]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256726886656705387690838569640420194963281239716087637041200627760103781157626234004806148409984126522044126952283568265301873440184812202346569955815731691494918970356662483163400759294258229057714293356378539646479793181016196327703169990897127168260792598417911843609369873714859998689164439005213811376889946501104323485125085755934693831842693215633228477532296503569499133214681634548287116594591274422452172970673755502351720666788058483960182828434134651724244427220886870000839484185519616381088687239017345664915448118739697490978738449;
G[5]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495820479762882398806118766760188213488882907009426975330970778124830502226705311902217392435893665946331253446190595833678970912370688344728648091941833772057052841937091872099113891255436085123824248517206272948131656443452209881379967151994189788881622867753003753715737666487200678329162273607104951110109256884055796026167656297860116747897392188645869519721427350813764064918483830722705529918771947583778851179621536172255758268926033782435710003157923575238516382618512471159016192401793462295974159028330529103380258190594321;
G[6]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824495885461657363360268696530396299207188186238172881597180641662343106683607128635195158635697312025023809598136801353534241117579032189092335795411645343863927481433242331619788403346597894500368782879405603530663416042926441487009908669585397200280314324125140578532406810380530514160179210812785471943337327355083250348880507740642580512601583095817449562936549120150996437436242766034758473034544408255381911978823492833444076955216323434117915629489310930414194381740647038770559276759749257626450864458660625343720038146611679505;
G[7]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232174775508864414498583591238394676864329801250749821657960681663053792874854331674239364769347564989278121697808723623247414884307259839149748138519185562796709650272958305193381230690867545617997430837546165766691846433380862908816443447627273175498082666424595776097119707838646635500041869234534408306705228390332475736263432494583630298298538626969906645598807346954182475990105269900851890990688777414388928458460528446606840442134755814723535440110016148220251049841341839590052412566911031089664518527962264259108564621149170708234215457662422001700097288961478191682918284700533108033614217509296880351041546618999898250351191830033404194;
G[8]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824479185114775756264140920112177946826528997419765327024832409990686240335086425151017697486436881360672773801842456451597907402859781510036368043915875205791845801045224586715812989092781906160010313088204609119718955690084657501611537069657454038552830705552216803840850533031384886277818278787849814812453705865727468658060876631490742143539785929006209689167098589919961131946873299293168109032963488613832920560280378433068839632507820262837309113960058357706133329521208480495528382018724083952579453694336253944955742761656586513;
G[9]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496860190074577781962072055128020061979153237400715533274288478437115035947630506740662372593898067522099442182006598829395905702486904276181033664979058753280946664190140600264144499797915722566165997333415784777043111961461108575472954733554261363729712354954164174580819788697740893184708697648521354346113524763382285291670343930633408378578612811824072410798626240074239810779614894274798037888424558757717278815628390727941030307961549382643688230608148435171119536611385154867030468203613840627906109342847369558189729121374481;
G[10]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165752099751766101640786769962842950346001115369995052370117765347295950928206182138885618529781207238163983522805609939357283967308935513766291572919747014356350704958805121167926797383742231445870559655171328841302133082994700264278280462662192838272075849193270154071410341381005210754296977744290275270995796637396952631724874897544220266798713426312157572017468888739914133943713430846458797812481258805823655600713267878194188855223461028719300907644453800617421399636501449375925798581608545448092774243702065804429557745907424891153;
G[11]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165752099816747996121748232540606586457763739814874628963720449047397930673645693713060477132288873458851549425038699749094357512771993754841550221498267294618734162375515463974617730259194936983063380868959448406592228731475827698195346332880565255913785640189924274968730226190772802693202267667176822956123053195499858106394703048475881099351269328303312154934921902463886363392576328864416440824174595450011264996453166789351197115675943192246196866226785461423663427362358862781577610951253047085724100565242815590735491807764372660753;
G[12]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496925171969058743669940763248319605247811647831208998478245048954304944774812336908191093642114928597947762282723841945006852363762401016934149844366208162244397587490307694224896533326661830146614344443050609899904529197636303155082763269419809784598827211875078839026117090063850319572270775276472159067826121516177835579796049282368171278180425764857377030610283024550702824830761753949502475907358273060331460062017099032329546200063987517975813646162735403211290386129021326238513380694599920218899159955533523468744566517146129;
G[13]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727165824496925171969058743669940763248319605247811647038631921939535921258113103399082276035033175254302574097306998481543209594715726453015284369938152363888381485617531031747758616690112506485080849871329884441080199680636875860095409960354609757679866521061560496663917682074739390395854368910010024537115686564855836042824324352632085895347116883435133077556432211716711890696114657549021387506309545433509961236441648819976422513834514797650878953327558938899849194637187537303145740393065013223109490646349410370802757617223278466834961;
G[14]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085614555903232014749445802396013641496594457008539548830288148773554953647919393594519178064120668032893765259160256727148381052448431195533254752820664014040582327444120566723142423263118500510035428475023267948820970722888799175270115820619338529905994308520179963183020310180787108877809683007715897640323485781188181656250109405573347309540194513398033450429042808355744510464193492942052038258109108455177871166449223389255281080447366700160502169911411161773027632272196429401625334243109557002966062167722554201105742867170297308022136687988886684846431670648505216143576380678631505191261147420634866045278103192495851632293100149303123009306526622225;
G[15]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460499385428544099517477423912863812697892456033388195120701513307999921234819540801856518882708811584204518243440689353744255171077952232898711232252945866510976987722063786812391367579142184571658788883753850855331041295810952665052543579831758419299263812291705061779049163698384053016224901615473728968019293265833077973010066710222313317817166305663410455828093631270919359177042570328046642588827601400958375106918334951906898595415995314424010781747408802253234804759498634328072151690975491412942927558223461424215362915807540817255099184328889274571460083260610879591383057955394518880134989964795952854896127601885075384791716204737231284443188875947638191349296670315881327756579099976209;
G[16]<=2560'd57773361470875804093833019566109674433695879417384223129608387403904402167250072637131979281911674448251581307236049970217993113520392092419472139540270357944122757113418820042135829294691517870570749300734767382744626488491777737536128148077755423536549651649782530533872630290384839686995866474746025453236905989775139621028806743450100933830312605902440972457822481872386172213131051713486456915969643903323961612588817025473855540583788159869984360660624870260581637277244282038226747660906391688159889165140051682871927764419536164447759634334870074950522544212552938198520530110500268695368886692961196390277476760469828313834039092403769145736761052901152951483646185812064761543797291106027735165304277436884655729148261132361475230091804974303192798411823915554;
G[17]<=2560'd57773361470875804093833019566109674433695879417384223129608387403904402167250072637131979281911674448251581307236049970217993113561902796670891146474083859820929647618772269115388313439615823221975419955944216016650585033401614194353125674989006753564381396031016308298716779700295703679500700976605838151877239685530420852926696169524400842333304543368084051305730376503645337498878820038491537959712558842238699921721976640734809033265835556195553419076933894481711648579441374738998766782663001023641115086324034735500341617617205367453917696533720749768509951064124072539492224902547398107791096452529077852150340811597580651342272739066681310652059339773569332113931804234353711011642717462285972996180062999105376826696120586868295671097138261404053427406961254946;
G[18]<=2560'd57773361369990237240164763066017403883580256574967142170244182206279687460435770516478933249127167916713661216085625552810549758839157686887192360015491853557651277330748104484302423664279556299905852019446416191810018355786979441072188829115311002917149362909851742472052929785152139006889259540650455088369330148547988560186530171027156553674747488575126707458967617234550212269992491986739733661067668058036416603709194961922489111354052819532385178583556984773629414806620404397006949689063891365721008552914493814068663801978845138365429046420517091187096705546896235074699788892843241781506913491699562380285618047124191606248605591485231664362787006934088737748288173785749740168574303926587142214111969830710153966188224359033858699930807575409006616386700714530;
G[19]<=2560'd59571753941400006215303823886749080183769045374841949891406173018625100446153867436854295960766780898685394711409067000301951138731849584122492530585391867031803119572913471766899532298840111389689226517124398200723414578740156212415759534376212567114273561688044199701202385905430144646443193796663847656849702981783053598854030390287601970870710499637838316274395999258316145507335996046742967312960055186519337541123898484065440457752522993729562037675546633654336725655479461066160046878813526609323658930134355558758866854938911646550543605007033650385402147980498429394172063423791216185821640460708777336745665846910527003330303291637644903474029648072921431773902018377111382081045427556284202092459194576000483111000011683461222653610180979370440799707283460370;
G[20]<=2560'd59571753941400006215303823886750415393128849802575100091670664018299990268994817805160564504158454275751080196444786205875766185985070833675799610507736463523651693118080352080271112120203711693751448024068793232936698057988978925603266284134506627048994196881821938626944893648157220247390839218478907182147065315337570840073941977051302332673817570110471934852685022250359055310692698345379510387771878492474022893039543983900814620684605813915958166129802285117512771533747150937659549436849436468487804547120718716017997180381126065922558081845499207117569298372260297895872591289214753409575537227109984193851137505920070301527399118343818392081528546433359808549950238525857819381598521896172656479675682443807852383826773148217828953759725248097406822403197243666;
G[21]<=2560'd57773388810864421437930531091114993515029669712413163117307995960202087713925947334107454179807402365928693577530566870122788559589242283487533487565738670107163762852042262104702100212243712423793892887281944815269082035043932591322461618076972439855147251437940225701575486993684735127369902047898115163710815434945552165609070348916392793844746966427403106676307998707516516024966495782605320629673856638571953796587219014740757375599196234353820735090333481256813182301743573008411453892970942972963908043186565769404360315222500307985846523148536328016739753329605078958826463789782426168487996694081738877802777038065447674753553213460601633729638676342195192961421322178600164545649364680582665311312750595430294642342629311854948169712054975829408117480736563746;
G[22]<=2560'd84855037739454993595159871597420124053919749070307207440273862488030192032212558413749210696905526655134379140441401731810246931774570251068240566710100896357759619930115459236647146989955767563035482776101039070529497731319759295847732994793395185194520008397464116819651354300578739534910213143935457022733633870639634601442055786309642875524886690755122044680094501693754267159500297314091930905011619451322914261047218020987990115659831389841355587651022773229533376099462041761134654321177672244669739769954215189673762591054469887324133509373330120671715320044156017868387643696575394442452916531770215080461310406798148710783645197151113221814638773449062869817111535808615403643858762978149602260263860409449864442476250453121906632222408032474849032393191465506;
G[23]<=2560'd84861649375964315973845885099264100136387801537513608548830186779299941401213838028006693028521728066952732277283717555851361467363909521179296184455927202482001987750497632315579928703118046611367538394692936803167299286428805606412658034701768743509314817590660924812224508407579536734776619211640236769979676998251562995202363574953005908729647980011515448060601399645642359458400124370790060710406651183845025981317767160321277582181453683371820543257341946458266591025846962527216951817767964113066560941004345788104127111549566591979747407523366798148974751320732712117642494983319304844752574741030797035481266680871101640268099812630170204929232326187672096792478223549668912664308143559077376551928945226172843895610333255526866607338085989022354895218269102626;
G[24]<=2560'd57773800423978826422008855176583123029277642765628285803201997566742748536679599198696973622106724829573889808031343835210624691112881081946153909559303887450973857100125453180148253299953714414097598507500294136557970380575469219513589418965649349858373190334820032812994859638980011515400011790318492188673083021888523781935872932284095880926471488320210078903155786556919851978122509421948854253108485449872715265251877329411323900401549679906635839605653735100236338475586066496342902255509003592073608070773817473146293722316127612917724205510636958216003006840623823674791750896939652148540243122395472308112499432603146343286418397436244511692694870125014424622689543047222304831010334641178633632153930014919363111204780600814695872802207421825094822847347565073;
G[25]<=2560'd86660014513223962792591522700344256656394165043566295334803139317412879706684667599858316908390012711808695590204706273281849749653704577103150234771230295437487456415111005215582377716285036997971729521655269959104895697520761295826603887312639993012247370159909956635151139085638832988557267321700436006179170209875981370833836602055527302266316599222840538486466300351843249809430058180607798096494616475867909772606827100514831964197184459933428889413114589280782888579798570999388814604548822033486631586190444310771638085185353982190497311172510527519998300552400962132437263779713097701544468750720520229458678818554532486736509316397430854306484932683337122853721923093159118019104673313718257537442470293835171829972846065434507551694202925494223314402144297505;
G[26]<=2560'd86660040339904447088341606940214871905057057788614051303714740170003409999004904548831534089820594493104659516864472504236929727330933463854983911684658439985754458796364559798969202574183289589357352392494493857816283282416832763272056726441079477312579557217452365686733395302623232897266941826687497822742593213165737500646486315658185382546184816698369803621128904908089789625610709444128705357996941756739383423747633121650388834094131673002518425449625073611147444280912029021025574829990306943542762510433838041930192634908687019392018106150361972585946698235718653516797411079687220164598646597358068292180948376156492133292569001462412445456219189454061265903245499529969661992607086357749446333194446933520870076840170604112392314206821047321405445801151439394;
G[27]<=2560'd86547644233906531695676106026161156479019208583566578239607352809486450216677615669516001570929543478177497901335076358174579187033260228160700169875188466113270107718212700105706625402079807133056700085445826897380974896620496467689823920064956900282532753057224835840687679776725543177713180534190585069232929923390163631021110464527397841792399040157021861302872076047230047329286133086823417158172256739972565890398770091725267703623355722541056133575462143959473312368451958068811119873578932523811603733505257039285898612448659298887274055764402361329228040492315085723967004304448666125833148496558280410099123211403822766100588887209380813989806941507509354190164845584450446845413159280419685652408381748467698641165369492874647102975551125882403184201282232866;
G[28]<=2560'd84854652053934553614824225744068398425576138286243924469359133910444881964043880193450730255912619995779529260226955235517058170709580779285044604250844259452139016929293360138414377969491272466231761764816328315653418620396174934592391654258862803586949879910372262027180037630616695497354326007694139411600314431491895677259171081897395421124119861430308459571171303817218337685474351649536545589222076796077767732146512921911998992560178609699942637148366948865566650807818831733112213802307554308859450844532503532434914574426150779348266450917564987891725964460805833766363786601695904506686177792805122687994885806342995595625548392149602303626145658448838271187680760123565779414086248391245065221971233434264110910762520356119361403581741477455645674775234355745;
G[29]<=2560'd86547203465285291722476897711523170322215662470489136199964365425258687618796678191890454241767842482254485900696087950633195676139425020183363796822585646957753994772561559322601017896453552951565056846357102701123343251697872808618949524291139285516304125834556986294941525794936939967933019849508836602219909593205812379781483528549500321976714782114344488452127648671166613301273689743610271155665938216156996942764577587117420717520379293383819629297856384922706141369936854336915652988724991918979841989761514408217020792420669820591546328078041871726725600817775990299042072179625444115601893932123158799431370802281554760383850181616604042407416453832512607223817843921184206762501101149985922119732926462649201790461988077059251509393662903090478818928292405793;
G[30]<=2560'd86660040339930616723249281478364409469494149684169156876183907180065310803612652682707429820522544802060219717174049260849377166333637832636740496601870303604881833727904251006499526246213438970770765580881942926698673929281690278951323288428312902768288359071074016326970065395701025897715405018028565826839317216524023778269385986277745167394513463098642504305076319007398379091297048966176490410932937991990799221850327129833932974574324726764998708434868740969447311800007938802840601357828389037315163352329964871613931332569709908165242890586414723097735761623238448198703347442762863190931327028395353976286424340267944254242241942933144481241993466446659963345537124336213731466964727284341293937948144492597175508642401845980199335334128984296173739887932088865;
G[31]<=2560'd57780413681355008640628930113182713118747241993654175804706541179228309369127573683999938698569696370497457919191008525309738713355954437446092296253488048015950072461499178519770094198472828747955556172552195319385416393636038336560417226815752650472389175339736506613057520632806957096675755367695869243251547227224463448019456243774915540885018416822863419255996455082625003472486060762262167339190149400213657869625192085703872641921115340893365940566305596723342529720698633662326534831363338813085334000811401643293780431883150105326523729919078231157666990626819444733238068056218527389562239945067441420883437153229134808970914586304085688681782559023526854160796150200587293939038236849230413914109056006735925216710428968042658839672225050217231019953394688545;
G[32]<=2560'd57886199865530329942500979468504725219262342551789626220586234433884994531359720903957987564301759284542441993091597089985542243633051169241798870794140110060464323935545682820563220851371760417112120254275065071192389442875877162959343946277945033712038650295618237360041749094450278904438694185100328189830107870039547044847311615817406939967606677012519743999345986633472814760966260554017577771477582212964688114449815403042413588596400265773897513874337488853541381155526932798951479789679057496543442746974849694243507004210082550434509737885365905240630491813613044925707157164854190859053948734208347143550475574254940524277625755635700828501877065435356060265949515935868046756277208794649761681666222814751042245035568391938795575992949067514249231137648026146;
G[33]<=2560'd57886198244661828510717820946167075054661744869106085268702554889590085950926884140769977040184220190139012940920188935375827133687972971161180844255580538655677880127167784186788911386627692921236718485460501909456197324405866695636816868275550904130651611465148449336819765636841790623804824991842553473189280410376348175148769800206246586893469748927590092426198579833753131282113218888915999195603334689077477667173091253546277507994270350770720351478216435103743304521535297579876460155617038482675715636854834764778299587159764509387870682236264552633617673952864527558085635061734829892710773319418557891109486627507071156635589183582207479679352539459990922440650724917862492781461391189887234322714568368312192591362479396334981862285614061863909836693067407906;
G[34]<=2560'd86547205173614332816597676854006876673828861112006029106104718338021488086319260357628662440212863533382706568147029747530161331968736551366646351126184278545318883029238817015117816716152439540122902751962647772891802673978839265326692502215233361755172495013520727430124014315080752769276098967533807870505236597722394816520752249939135766611637287785242935328908543901470626179201211130558378170088788281237966081469156827677123939718367790698186918717123622929182531830679162787537947182123278220320253269806216714293920028427937999227561660363970818641119141950695240124687560268842391446783164413865589513517134934515808041262028035705214877863983036584553683309786812124617710672155269784950114771993987457791036933796888248539025192891669312025041445112653160994;
G[35]<=2560'd57773361376689771640823383541146674820641875135557686375809918377490925896274175771886835779009119012445829897850514739139367697677230512565121001098651049848281158363423575448704338953596310138245550700175615095503221166721457764087001592668020377673164499299874225816933830584719210098801882536817742789336583997703670514839420452191368232884927213930549656626714118841855819495705489724435573353995723927971600353586470542664683069599005486081779756057562287286607922298551607642747641336647721244126282049401819907658339136627923403590071666370447904965607845456429671375057304781051754315152755700622566356438297372071129100002612500246357226579540685109458527151937167414079700153454076079320762181876950410262046527407330469767412667707042179615111526910932427298;
G[36]<=2560'd57886198251359823119006638081691267587542112734823965061610623037391202157803115475415536320492323613731423979182718487757005503734268283504487936919078104815512879911770451515375915885934213789432923363804072007271723107151171906513727288474496254330884483879377053165239157537327101064753763369702581193165903340590408446928324079180197919450013856715032160818635122045503640747795161991307662186581212037481291151228927537799176912203291843368146040406744232580418714678888970654688312112627363588453923143766115828822729031959401575910443405909660339793642719760284786049510400893492405064543859779738627237800281116598720888914767381959398841655297947726699818122847513534869788353168845885579406593484043487771918654972327693103028851851909066264206671779610108450;
G[37]<=2560'd57886198251361362884956388865772942505349142361011568304536944642532825608609275863530084300564537482524051045954764722440046020388115257587816074135857998118935803149384679391100187492299487974666972874027731499098130286355031379774450606356847085229600928905367566439929203963276667129702297619643090131997664219909891562888183374723271533173847777381691614987168625654978850143770126262442900454123067883181113784275584675987997273177098527214706310398953347579764506129741476605982000763834511910519819896277018530589043427737994592330564976826171245288845736986015834338315999576084657672524570582069144797650123697203622341891479716776735094324488684274768408590278011902297271992909335513766118439418053524861196237018582435903010529513927821236328914538484343330;
G[38]<=2560'd86660042048680007930424800345681004176341087990407829576227206209746178345307483002399604700197562652106164500963212526023189340038649793980339930972580352679432083332034460513087123591385148125419820973153328485619738159549173698594888409282211571877357583547142898306015112072350205247174317127936755770312411411693586027040434386623466388350397529896710233456477533158749789138680995652610818576500451437259063655345821948860294348868394977506958075541074921727366642595922609965583749203239356406210815096373212591342724953449309696679918901494839009115077701494686084580568767530838380572751595092140650073784987852400515678063033849267804834436483895136116412217472711588333051971371393409306361690400103150870117496165980206234248045291160861965942148633712534050;
G[39]<=2560'd86660042048679905706670498856373919482003898794175655597186442797913916598133336510808291049470179530826091433244407161837483689279714717458983399068705608718463423982668844191285205820308961360787975730947033228784205554511973870570595400115001404958024409040150363471546836510546252112220254743349592469762208251818544966223966506781345018860860372657316735475663700807050157946346010571009956211765691703288836572059946548020617996322140705043368266956776873543059031412491587328380629822282492372629303267348342173169253345297480883465722242117419301415402591205043151548128163893523847739584571124184305104389616741040570007023986978585829369486409042765540664523465812738604160994690648323235147015429313378754547376378805199160782277901230400651992247384439661090;
G[40]<=2560'd86660042048680007930424800350808207770364210028497301754987863923357610205641372752935678039550091572522003041783745934312988038327359585206407063320275194926839170651772835255610135691602168551775290829420238200378779123079554976408936152257332781996038037123362327117539134741957429672217060409240041804235564137101809056731910526844491126094189188948461662103521570928142203358143002428570163069986949953749997869139193198907139767167871204222884272790428141546375064702285455706607297118214720164359224411534404674296895339816798018614397846225868141849272260561843913359327038154053219650426720632769714494197370102395743588084854312171857729955167229401443802955303810997731640855566890389625240489582995154463878181999214972803938474639502074081012871465137218082;
G[41]<=2560'd86660042048680007931892520149873807400491986871039771509184460038271334125267982493978923024194940154785157601869620972194770800722035832975423122078395569578541867574848383078727147606562615679522385202966964639204835346694710913062255413787572672283866051988072156467524611715182674362647441642006513833187208440702160149722989265282912175633806154421244849949726360240496799968087194066513426619308970144848505337070367936072532594147783053654717921663249152773176171907412744127310608627792249177502451229167428495730872454357984598449845549430027421692292552886711230882632306017804662922059916082752788015874164581842542824957708070717125036599105414948250606094621404683868124026831987692944991524704476683897398499820063823090774584083342223360698587011382125090;
G[42]<=2560'd86660042048680007931892497743330318551888086268535203559603953441769403432097744057686600165799285004693908652298606441974580378356132249784747880817894661406182914340337612737321449103395255548634327765664635831759587097516789695604292684211039876843469739824805876449568267560585422605835535729535030097423010863997659361251958923996503899152082566960006768428910889079586332119143005152560948804893238292324046962336948643652418446714296728377833536365639073129899532850513254608675801332265714400247117818624953783022994023433915934818755110935423999759147391730381806265382610545136879302785342101605266695462556862976531700785182944195522406297053197556783027464192301303883549169431263102333241514726988110648354672251150807312009905258073014901885142495056241186;
G[43]<=2560'd86660042054985355860246763780396916595139182190559466635839068717620643410983751612470973283878043979682038317225596061411597801122422374198740999968555018281259349058096889367285539329803776264017294556388629227213048382211949399230713651452609736672323414140581408963617265023746837550025679202405152140389164706442121713283826430504891216959352374160376029740971943662039106710608550413415630605525773289228953698323561448539950494931644464335216647986688347306402714011952472905140060776675150709962334424321591111899227655998383061642129229624306436430986721559692071109299575757639739600840157008186915862496780206541075407246397818893784681180175316913578849787488901905584619042841620919470650133159830882409910802025923429163225524339952125024767402361628008994;
G[44]<=2560'd86660042054985355860246763780396916269160334582353078132005935403743489602691486280209604110762075032424719011073747437388053381021371005483095637757542075924062003385256723917034785986875967151561658751595043770639837459476679911982232481628379789530947174738997808872157510708946636806088920525165957039325218561570934317108747938136780249097782592875767254241488565205067232586220883402529424569300572553643268529189590555465755051011317267163035256224075468125950843040081584207287923207580087792820889801474417518264917943724673615212991298988540099568322964824683497540272962938309202119133293683989582941709871084086885098482064614193897428738618652714274482302680832113905815511393128946997365474103712990967494320292947876922398638606109883492192402488804123170;
G[45]<=2560'd86660042054985355858778685563434785797141114242058606618279755029643986252503841159238337982373373522297453321708239130508181193587222639643175785141262499175365150930215420476322445313099140979056554663258885464376960180253595363327869146774646048293348241851738589776482382411546458591260279200652678111827201917596216500602425825785734506640757584716654700261918021446821983830852542954649983826490495095138826222757346412631606641200969722826912266526057138326855753032592553269327441363632816523213364267098067020947763252537789432485641421847507823980697786264267176201037859119947553721497384684460383506658502280708795646486055367638096250286245814750100233639831026197252572770639983663269917990114237885335568394672320313948658686073541491198935783307410022946;
G[46]<=2560'd86660042054985355858779066382405788623482250413339828470726677404109926983401609525569057367837882879673716659670988501639059061533190796507301330288715979317615683978991923161455227764577183962619778907542542109472554094303208349837277898053186647821512372423648282563326024547826524863117877759415844814019055182358143940423187333920642170143876799721844601413204186161691363458288353772713795744104982268007109471638230998766390143070893203122554730045298802080564234751843798225994759853235839194095432386979750447943741384743658650779508547077193013475970813944475127315017307654525089682180161533648972774299163254859081500767493269254686087768828885241591199416773498659247008239352651124664780893748817581582716583512186618823542017140265328915116482299724702242;
G[47]<=2560'd86660042054985355858779066382405788623482250413339828470726677404109926983401609525569057368668773025623400662470388244366892743885762918170070295927483656670800818907337668544186404805592140459291021099327367686731256291952018066407275993315670813347494785577955399276487194650408226703891566795138771333928359675354783538047558374066115593308217645274858075484253240317136155771767416228797557410093885220710958160720553639777988533137201727653730245843775918844517972731772271242985837118417244787913808585553420709014784645638265834807526002793998618722358228203581774568486172236176320791425354577624918312860363721252349022437596724463935482603154106675173606972682848715322131912701256410406167811418028175130148382228617059462605469627935968313951974811806868002;
G[48]<=2560'd86660041953681068106635190087510969713440941542676464483039772789571657224392012532835602736332189700746550521647143070512378250592769974059210208225936506010129890717310579264561821424693774201934009037606695145169579412924506485936819184245897881768761893399790443063072619005679457830464831728868427028195338488299870666971059537571240997379793854034426032495661859584850481965099782141472667977266300874312394229603973180882537427451472360673258426457664712771275056267509506865999871746669068012206726090742205757068453733365517719733107360775319570590314469875004886307885756955132495717927761215427428718502887981193603519249144464508381707651751396031120029497271158946974718152538989190001623374725226670535215814444508814492992410851889150492436499064615477794;
G[49]<=2560'd86660042054985355858779042580899650700482866746678704041470904833733252705770564303813670944804758412697358339856341522116479376847005978313110320331129082551712200291654589377646395484314385839419833649330714915836425648482795524352252297710274305800723421933711165455647250079204721682755532120936562128005649608726034722942843790817281561864971362223925547390106041092159671008922259389816604286851488889821051840777191447248525470367118465450615288674990520292540887701672221537125054542909406921081405933303903026407698916964516177325423005288070893354234844289146950189296943220095384495813269597692297316840121679319147110179317869518231106459751515772457473682988224202063375939039064015566192602833460870034510836296665604547330546357519043726408002409414664737;
G[50]<=2560'd86660042054985355858779043980968140366770481462086620545595401796867242285987613106704994512471427422609518420367343281228865439089590763145994576484637848798146797928429555580067697568787044605904722067256150036211992223016792815597543373529270477752378208115103125764767289351920362471162881962336062648556786164643667450349270245713163997721014453671779864593900645597745677344744607891290557220722794821489085569056788105393787687549248706951708757226395505280418501984089322261309101517215763782470241646217022226204352806139378669960440612452417474836242259436480489947332242617236069416926492520123053545384099127405148844865968382427437727048914443141877717066782492015465632299338373606007217998207839972801816214101341331188259394178043162720768420624554140194;
G[51]<=2560'd86660042054985355858779066382405788623482250413043352435936699269989113289295720328931914268360236876286703549620207161845743995848687972284182021581571963249461170347198537116720150521568196841670154613461642106724424343503426541990099238091052445956698245557683529622491838211463705697014712530800572071296489420018433822141071026207112230997636269996911769012252172717744846473496606832186446050599195978858900571801623932933941702494693701636250341205809441503305063956861696266668222810482624494016976815333944599894284133570902724027162659038813429950665570787946319376272068806772826657803399228027775516171968011000718870389947345510997219794280156784192631387646782193353033551463137019055180906303330128059904681487917990145720358641865343028013328464934478370;
G[52]<=2560'd86660042054985355860247144599026105824097029988979998940762276780325789130097412983589890060956835943811174128512144286711561552509151793218700130663381006090596347712456249535970544951382425260880999576103080253532286961330802656336551597258989204139046459794367867232059867562542042259195000808293139155549836330691145335769872881982597325860974691542243359892521873305329542028496531215507817167296821851009314637021303705301203311802510459399997698577826067418921123933090242315870125008614593761434473526081935722342557341645076228863805822445748326863370590851443957362959409675012813192663313938274266211410176697464011428840929611838192511579860650586063302923127187381674738472196365774868982457452673503020967358621030659055428043928563942684591420307260187170;
G[53]<=2560'd86660042054985355860247144599026105803723352013448569907098332314825916161197528325533736446466802263249853318558896444694473167967781433179911322579735004264415448757159607884486251350952810936618514875423816401020935806798414247633452655310136172884986605128864547303560169628199684359852190075294361673052454449545562569846867922934291145837093132908418921107393086182713271879202060377248661168042612721595942915594912041817455848479559102792822809333264612690868644068424994363203591589712725146368674504599885808200393699176748664471126639761023891752123537128100812932515685717003398818768846329897148320503360070075386091115658994810879691487893930201329435996319950187571744456848164786539646008310179080421345728263409910618014426229044018717371625854717796898;
G[54]<=2560'd86660042054985355860247143198957616157809415273275606401847801683054913857724015869745738009495520426496013595254019616276918252706559036730517567925473363244271953587105398395330906366393934964797975223198396016120608260661861769916522741701562430487704802565771171974121498748478756099811215555868397146141947629973775578296202785969350407834282082659824478794036290976727007458231432687636371322854234783724576756840168982645647592586325283399145531717890934896224245883118321463189347486181123411894310714608598622387317373797837423011868063478130433130658438155209134363490799289507124301229220315490872305174607888249832083008571358343548194415762936850371307920039557656814731410650870255416906436886636958771533394917216612650844630355500677524331504388270072354;
G[55]<=2560'd86660042054985355860247143198956280949722965719013170516182992918348259992078620245111975407102989111853916578911136083213718743485772775757865926940684976263945545095835835188288633478832728556506922216040835923396536415940403762396032571662521575280428911570127456279089384340186277286753913700687373968115321928218621365620025654220377864661426507486449019759142129249239478096336245356588196548407353030685718024443562275088829022202809914785289904365204312582236277314656335398274506109220768073106488716455041809752306896733531144310276814905618743558243836120827268793661427595130606121998647306549936409736935664975034252464923140002294332016259704076187707574689083790004804657815154570100538770143114324124284153631092209864453133829764091307207712097018454562;
G[56]<=2560'd86660042054985355858779043981309953962880414962069547848095075847775922625427489582415750862091967253328052725540206978325213666061739810634858717468967353304268472712834328044181562989527012538596253710812900954806040517669379490114845623771986123640801384449011394718498708721114687868235859816605125059345700993619764063046495890656224728498081090665336437849144552598671341643630041412567173661725035643574674330802730444146414903626867336233063307290384715540514927540493527168620502825629918147969105637112564149048525634140599476248418606541400736159309141458345063456857152494826856689973428975043227964087802898167014490378516400034064683444741894127522423793142833465796575689313408021018989621762729227017912525848528860760229580771970275881552674274953798178;
G[57]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653889653071580632085654872882052773954860466945031344557388528491751004815415037772754542432001558774931037760633855271045753308239093177283751596238697575492571877863587228649850810627442910149468310501082325262472746958994887076736180610419273367717968381675228900809217769254646675822531975137636038620897956612191230723601761079561482789884126472727012933821701461639816945634011358402017287160713397811586285965706088767883939722716158734901187625345536477908742564081081119999404687937241791681756677956692823387750957045160423229522328366853541774990458755201168200148209490223331170614846925008065789226289753329394830035797908724518890210448878089486856545510497383360217012571350376994;
G[58]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655774719271138450876403253247980525681756927955966313408893360426260923510851124225656679336182992485485582553762903069025764545301208114675219999682369604280730677280663085198483631923891355892708293046662423203514706204260985181959773672542115924493013880045541903868308888110937032782676668021161123182781339203518315111239342409093632303811738022643378105828812942801845280177714538499525275336523047318019422703179843371536885370287948675884308699991415931439016261119539117062677506538690338435646801560327307770818536964588420905074823861949394928438047705722746387671863216717295875754698440463367648245777249910330319181731115072248424154841342736256206543956355384186676383395750178;
G[59]<=2560'd86660042054985355860247143111453335554939794227014796182769643518569226213756921341259859584655847331927551925801083113722239420023735037221501403343888797101784485428091297633820555426628132444240443189637533982397144847074286545063728176258437372280520181472519077892055236811898975030208945229754974394771557861532894593339218546953074265959782279998383053459704937225139156610517274077379498937826253929464335646026284249469511805352044913585632132636556730659051006616145226591426780570264289309424192224557073134779761862353093720036827761563695692023726541237184707798368999946478445971640413873826589891622623607877163896854987379886470855753213378759358483658500020978676937666804110303889982458638106352172301500584091171059591696502376120599261557794747326754;
G[60]<=2560'd86660042054985355860247144511521825221227408942719188721684118615840101486130318455104011422578788422303091856281883711360084916977256211647218502040761647245051742863180649101461518057094087840151819189108974499674057614671235616422250522400472752448260249259811871545899956176160760290117877614210040413383699659879470926122939900051338539712209862023458245405854678800980242689599924078883354409708333679516001107317269852292268317850954089206035577539940725260913867976686933328380837615663909387119286253829702699469042640724440276197900248930779584646031149548226901857160232709144580209513902232730073611422576456572841936087366733901272610561546622627932260379133331353589838330387301273102999180562501618591856542526039496357707062027424395229927093319338435105;
G[61]<=2560'd86660042054985355860247144599026105824097029988979998940762276780325789130097412983589890060129178833448842981754766926594890001379147084396561766514151442423472671271577733176472177794863122290117229327991146330649779988599876270363413514204087290129857463895920198410407913527516136848088444896902525138266280326727798974060509784296848183943798204047143464899439906939430535322610359458495582398461804538122504965104670389639025874127542309375805503055588810948109769636623272370047194653534521086637647811481683316443839443005819800083587861183169439250281450333445303589191044020564224250397150975415711283255824104345418673478663530374775470013642209012515958914020476419772885412931890234560281190493717948886117424940064712916709621142325535805826320419707298337;
G[62]<=2560'd86660042054985355860247144593557088286338093993996778657407142111977074773564704401113994398020312181502375568673229299213298229086782089927547314589499022370200138585108553134264391182968735434152203212672921688901567165354811641616822544281512587480774526369703701706251433092417736083204054321384018794465260161047941010186812917382737087082984730047006516031777250047573064756337075046695917698846612860215428814265313819269540558557398439776460634922058612010320567848013805130933410846600838907792128411476653137423063234254767648774077996288412474606468611190359475636498202924225738676648212226453382000176794280785008176911571084945883687709541639425513238520573787005622755067570683021279389103337245457078656686386079229029317081083556429232540624452386431522;
G[63]<=2560'd86660042054985355860246786176023733696335048798140859661637572745133132077075407094941221655193685997491958710066308711411961925220130909958373031445522292385843115017774306012077355566114773688622847285383683582358559077329159837360381247724659056980258920352488570206225349141535596460106540733395603300599394190034753034850680128499067724535410393039934636073457212601735522974449253511152783567582168443389058870214523663659786863532614635066038869152188286885842290689064308722891679253317057604820768562795974105254950073688806397090219635756580492061551606914753115685502866408397124024130879769520727611290296888003994957005883977697732207336300379910097062204497652351508726415194368912322176652722470555414059290444593867646609145355676250843675969867774829090;
G[64]<=2560'd86660042054985355860247144593557088286338093993996778657407142111977074773564704401113936328769805573782886599260356634602809554320251888855117705326231601099455658690652688217618598901308434824433943915474864242467205044732768881459294144747317318127393209868176211744042545107818486254329886225881362754804420122997466889865379698418997204621840137374200345484093910976585121423400729312662713754018547441152143030815849273285047428102015827044190904933758651140459233590256543605767314173462727484340809640017929458352103275529290362106411955329236895162689862028410220062252259005897122191226141277063379468016527152272099392107451889430174137545550752082926851448367363116329287114974239064637951004550955224348074593717373293924037810464159181395398927198749598242;
G[65]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655774718399874576845311263545621133587374865287058419940707173994009136814956453350768510203102348981932650334168318863929303384803598438714880777773760653438309467308309674333580766875460944163258553664485399703350512389689746009152592891465470579617499246392134692305691882188906687901755226684312602276243870296708998556735964903520686379328169033984560048037094463059281215297534622478298795900231157184848021832456550484421748935713389747084723996705060202625306538106371830740489994778052864551373399262997900463051727027345947204393612565134831068945300460823215836937203120825596631300219200737609154155615517590363798456755702365997121177983711118824673426344802772334068935371661858;
G[66]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531190653655774718454327790191084627349621299974825006574809757877462121585811598112810101427378909437936333388922662171105735217807267199793425598188658135183563724358032057353479316359114754616554325215643178941995856391230901090859599500630364463235959368824600394808655631443543432810959427618684036401442414844223442704537743259568172663689822152367607873679446798919686547135026592474419271324488057680884899658831462461733081526158376459253335403841000626453863934717473404934807137378114636605839740782529376394370848128524048014330580593944144835869571589381734225118077837757559349421951348300910035413251463717639437790513128612360105192064213447571513325311286738451712693242898172633817634;
G[67]<=2560'd86660042054985355836757893132759216999050300176990105433423042907694069227337621562829993585710125964775270602054329570312964848286606141500531370409080004217179229087876458524573909993767173353541741569983690097011452215581692943335157711625082337273452088155362138289609015979491151724013197270317567215016397895589488143744367408171640028233148403530609947223568923703591532337434080808995551208032112472717051380803676170184201384443075252129804075351945885496179914149724178321715988304098213391844187969658063265840143740972682405958357008644602236731043709338815233073262675242050602336722143889890945319882037542546079300604375657035822322658406853107738162463497108344086946922613949873220305811541439403656605271856895022581227425901414826423958301482927923746;
G[68]<=2560'd86660042054985355860247144598684292229260451362764261987656577392647736543370361488313710848856671873072791647228847401301233737022303104481537360942050656559379109093707203561310020078329455616609213664298073261692643884024823015191459955184622890351912106016648553401819722104181655546115603098605602283925052724782344142612161115776715102522772726678600693028614344343062763923568836896432823850079449204882648266403309308892407135748887072114713015499792289361892822207599883377413424244026019710030176048684613618462378857121689125996320360666288608862423331095099705296092543804564100124194321437686435841939382768673574851536518314568569887782433744239917473763412468844755838549484650598041515502392695080274323693426528701197443020246240241189182231408333169186;
G[69]<=2560'd86660042054985355860247144599026105825370384862450713255361959015294025087292967727262403019761437556893730939222285479208882657298300802037575160390820663446459910427025464988327289287183046129933888674557455821371193766728291409567502186905000693240486376757989222554571598683229120888859653263524696001017833907336707490699150744578210589003292255020429401758824390483464760261996791101039665210830411698043690738605065655946827548868455326266465220751831286515792054482699950551567349497745834860048513959155597774589812378136743362735191173696671071195226227253589540277172586531673396101711690290664997436114167944396052162106362849502501002874907669478497240864847453355389428257027314580058540716784625166937389844633065329991770550966658389420930642393390260770;
G[70]<=2560'd86660042054985355860247144506052807683468472947735968438328983947491387129597609872627186651582024600194769475967913546040582144638130874376358646389318118814786852448844864649616750418145221955943826192993427732227178816920656271276905585143533586373115519879198834973942479680809689136819032576647810312732595572241699987593350080061015163659514017086081785146239875106477794600524685253134995910988108331550005681068184799601299096865758881197042238117027682965568176184440972070007071685850278791236878233013284058261027277045670555915937338480331575087435511173575574829886103561003286505600594130697069131580070588727767626265269615924617269111125896874772906631908154138492523244743476934718646027340629865652900225244263688152028139895812604781531321130020905506;
G[71]<=2560'd59578778805611415146675009581581710277691063045551933687756480398422287305889417379810347486441127485821052919679468113542889452684809722395700140936045022572934856316740892564662612527775299204707218185663838635012072754076111058190931232646246903284622465844734391942262056614048354950998749653954621708730071231384805927464554913100265626297716474520693310320586703562023117512497681822088322064496627431618705816210851000079439549733964673296766382384830234107507829212973462685859580341388056333822408667819115709266929113949331942030765735241154336105484549413082790808164475594849201598380667340462756895651089301958848549135503799510269852440112386488122331536158859401750494586734685718641628289919093841766310500080242900024127710319686136400082430937478078754;
G[72]<=2560'd86660042054985355860247144511499126662105429321273068407277388151938834367485704448074122569444172098571526876043165783859971920836969264760530889986184214714476462825495155391096180828470557181509827704450606097509215211503688305040483176269022017505845808269496127703269358050071161707092074104791718970772952653536039658534041538746737519884610030312878945046362214805134711841492026238512161881333319600192118535568830711533085405163924568357858375656538450464542581387128911893507230738836122342122599229603225159031928116892112183813987831334078163660952121246700020305227035488720168916218950633486959406908687460877728095399553261757236528956866684643708270351675359414887359595433733068798101071801564818935401427557464124212599737527976729175141628625738146338;
G[73]<=2560'd86660042054985355860247144506030025673766809899539093146316106265538579527373894217208035140992228093770572926673644688048479952434091876761068352954624370313967179694144722519396115596716221149993677036153553749620405412492028321159047416322212101238817406986707224126155932813939280493474565106163243812093763248383289461620019636871619675083026048451029932647327890463018525846330569091012827951043961281840363813652720803421450634459595725809176904449959904946528405453617565759058238372018608034173761612594819174824643003666622470359816268396963607342574155887874068820379188517184069791924546505855719533630439298370134457181094281013101904021478007737640291588363532012684708463746009272487763618777157431999954573528906051437579347480856254041877843835921506850;
G[74]<=2560'd86660041954099789006487133204903260360956160549643489620338436618377637842576284359863362919106309704243689707478965570827087656974542979942899829084462849611710618939249259608651433216280325477624001316104317596466729371969140954012690077284070616491746351728564471749830002831560147671056706250114477967642600397569096089333639873237374815985680449617611473202653341468188389253981682060228151357854826269269897619172307658620798233705706620873171621459991834543602373480841465702572766633951399857104105277494966054984314146440101192436966681634547904932513426545098027989272415738681311799297143377554507886856890818249006286001241109250814775639853255995094349878596934873475517785221958114450158264812106537624759494253032273056539456887172795468571491207787717154;
G[75]<=2560'd86660041954099789006487133210372283094002980229243248581765007654265653577472194899509236465242444698557438206565622384997964166572406234100477574397674777977505156139830132600223453848556708268115839502061869003420388328807831387577338221680274160140737353483060194004219894535220492435436638099083021936946939639139967824451702131676013475962351090698562849120246157186119729566585232078263124535806048274395725373153488509753826952978246979174053340621456186806072963532835551810894771631448080623550609249689592193110569192389873730482553764511745817030083183665190218365690879571174825385991280416004869216602169328363378343889459927877136698575477417128475210924716016187864188984710543742423461974587831700593124739970235920631999071281594898656945873596513919522;
G[76]<=2560'd86660042054985355860247144599003407264900768742917205928978690163070087408492480637134593336424087829180468219361015914975598451995323508157199382690387690692398844843514928702170390815955241127201596505186844143653741703581129775648233164490994829785826559032053443722600385653813081705720571192837612192008789895713581204777036768429701283390029128714492492860866413535988313649888274937865120070894133677752082007591688015900113548459282696583556119301935464465004416053920016584001304036307935383388149030247634916924973060160457136266216231745761323108368693178494608562968755471783886477741817760726462323763538431370223079186111408194139425030021432821272200460005743589200945611397882829013036913810155655564988139486757628315312202194418455979459998879175549474;
G[77]<=2560'd86660042054985355860247144599004742474340157850242275773905930945813336110118196240539490019284497147557838267018715923327516985332458326214162622923935032900007250338680321292760895710080642733831080771132276743829180253147307432997290084635644489975363748648430396123195922767541394877112594560996448552795364929996576891672177881015439931564850225635004154449269300794129689966712991918235903256491757616054739473066684970639531734216110210497023947756414714550996636483927399207975705990206652969886904718360475734763919556982928349895482367292716115476342446774992956956151252498761107452974814663281784497534204432083595228598354775546782281615644757523107013408384213577019424866752638179442528218812136730985593652630334269396304630857438406952165630624722461218;
G[78]<=2560'd86660042054960725594902010747320149636123739696737298068478322537961717678834482520817700403422358152770703089804200239874430140542010196752272567030863787390542375799084797042880740305436258738701590595005273685970718092719258284346416099842744389568146106365680795020940108979300459124745005745541606269281975675153401601355861428425322813332853822314868282860085603518697367456251787738056850481336079477469278919551948737819618090357466945106174611703508873103241356755282912505867187682504286195515332334044507939923872067346420391291450201267737307196242266351701053576592209146137362958009141113321913274469153424631734344853704883456841716171248282511082540215444006217020418174976790118549107329200324022701764190600284643805639511798376487134797608217221407266;
G[79]<=2560'd86660042054960725594902010747340177776520806112734551072445687533085065021448737070947400136664116789823449632968933407100211141072534280403769520078569537007792782613308474635802174537698970690809478334163570631412643605553283048347016505856194742070928102753525115715195323556349282491460458912876425113469267946730167935278877587537012328036693322053917166377186328222421417452562140040373504779528146445317702735030594897981370553186876005592345917970632889970866951268394574120635906845248615646694132609550556497211472604097622090146301841019284956732129290307426459296785387053797423353574007693950943331632285563368237321343236561559080511485751047627371120384481280497045687940783478938756780680703394917024408763222317734320903198305034840010565975018362249762;
G[80]<=2560'd86660042054985355860247120704888478140837876365123543014150374342850668582094621300469630599648230045742933784209142216389575425264556457922311286053930068582254622325112018075397164352798510515175743577017133975096924825280536745183882775463013210531701767065164325694470222681879094027781227092124253891209974256562213127667449952245758611535158008384943523014702263896852972198345773215598825568241371935340033673140086260660029269570701662991495015670057665468054858190583839025745492539179496075518443982113647629562614224198611078900088975010185705946430345852047500388605612792166307171121399509420106747531104482716050218417932545935284048716286685620621872573041225179656281802941603212553170821511940296270997912335104981143764707985385150670693967840854286882;
G[81]<=2560'd57886199966415999422274459868880719125540374263590124869795440374651327475006935105024159671050131151629198127377876542703104025982922392775671051129536883522583656793447358129814165503768731187588849792514834040544807253935283789448867402026705581432365375058772472597764965932808718781213030096311926565294185957855310110042521569562205157534019507819107854355152510317494284522903983483964605963312489473798774998761307931619933542514693985202534158387607026119398615428324766398489587748219957943248718605013661819049738657691700116659963079334453258255115311280263377575270159758431180536737140130835363759448450906942390758515895892558919289980424573076460337180917149852867993710505728622602071866521405599262333943164274023264992321184253293518166190136775287330;
G[82]<=2560'd86660042054985355860247144598684292229255166442635034168043483571173619710347119691144225030345827783212616222410294779761664479303518996925898282846266761510152391272741003190926623569187827830321629584262815111917596656706924087217393595876587508488968085186850687018244869998586114352220825360249263999775994728817375979812312492335397673203863302790066154748820302833669594020234290070582495200494929173360892773760163848214934974637634110348177502057929162636868254278830623178642620108843250787630827113236425449731118530688061698145372752265186338644811567914707468253620627016699072244012274195258088502328593653161690728502743258132518369470836368284298865727335683902707471302377458690498583886192744776199938910473963751447473945313840479367679935282310947362;
G[83]<=2560'd86660042048680007931892878474455227177971028024371356884811529049464620789125649758454898234272000069661172069987269389899945767361027574550972953530686414156658146882063111746039616309348358824526389848093296029675936468034120445424222211600742719199081588357825713506969184080579763331048295605712708386042479337966354451986290223333162107928880627555641215916709142920994978626416705217902414635832264440558822987219714564201291986753954932486082169720587931507557958295163366806492875072812759787144098478572127948308523884977559396404699160526520479526138165521289185352674936636031862683817235010289653831282257759622960847192343479592912613726360950245590935504593119468479652345238828060076678734350136759719261592194605077595210590771535247821334747701596791330;
G[84]<=2560'd86660042054985355858779066382063975027367342790537400762351507145035035354631882491076581761791269452033454183249344953585965394076337935338929067937815323622118536437564297059738643985622505820504106233814091760776962499864597298059636168145275156380296688159904369128528449753683962911312799230433778806225091259387969225469171675201128841950542531180116230576449826367722593526857172521687380991124864003137484864476578707170847913234971151192728858579471574281800440108831643342639806729108253011705015817802300804819006806509556132826791595285218890642917261770516453191612904071342140210892697080297449383854621207259472932253846052618039414465244459335409020295559531631438526291491079580094505907840769648086836318006592823881355453236395659111836949496283144738;
G[85]<=2560'd86660042054985355860247144599026105825290800106942398952294747558040315764879639160853610891343641288103171800486690726035351073673038897420098791390589178677549463196067503209119942093911134633742650281137952907541928838736039120644646931213431112304087705918212662505290465616993101515620308726321822160039891944288240508538304355195681045858672879005331300378590385772671636360499077146404297835592209696539975963729580103811198511037593977261690843212160678790092497209149901299896578574417450022512314644223478594860607318104626614943274593030863303350193129768254716719146242445724555021203697150864406182823332110787462630238266984160936066412740342336739627906476212971555791033611251789021068735798176701954453565289380761074629664307338427911253556960591749666;
G[86]<=2560'd86660042054985355860247144506052807683468472947735968438328983947491387129597609933533007353684341990834195015035555132862800169749291769193498400956334536367377488232563817334060775311589028319499004636252388382801225987419238993976401404890105498706757207668415650809388003583954191261892980550012471897649945546194087881745460552090656867092022397398117193406979658263660999529979154606521646016363548806246759747276630646428830254854567210377701679472127092615248509550215121741755238221651842306972526149331062532715833584924367662404364017771944166046262895022778674661432141777272682723655851838789731391531005692757746195209800003240536714795470478775228159959576119964382052626711932844204986669243846253798022178028122705615451830431736486204494364140944630306;
G[87]<=2560'd86660042048680007930333045462269438292872062652782987313219768042637666786329122335958460617666226744102445578905364904221461546927122893717108422029525645388751312472799921351044500286877869119547669424756898689829950269766031585682350250802738512990086600498257138856310699958638986089000168219505650452112645792298125168043355099070288093785806974677681179875429651395058070130055538199697219290972676462000385767399321028894749768463796500316714247386234917935903966874879825735126556867490207321468054617049686778077196364220332825960605886426479480461424307056476950210290425255119077691922776496538179629287074916631800112674371952466862493794321215866845955683019940383199952142344488797901438377077613337058870934732589916097121038462490224294365744145232962082;
G[88]<=2560'd84861675209395134570513491296012588649149499105406319276736838570015987485756327961237633280414293741586731088976136143971972148940487030188143946429331268596433194112333477537741339933425127451231940167631068619325605887688332015316319583609062672603847286089448040649878095409164732735514694117834379512161136744289961940515034067303877205568319487864466326362184366844823824809603763216310873172285098423406636309344349882612942032817949443939487405824542659607168917833178514602112722803193492521142690442570845502604556226067924782481702160068820749451593355367918058027239620695017180092248959471178729969370265186115169532639379003653673051828582053830937560743687402763418693303907915927876440158786880604316169809002092108465290557910498115674775230925158621730;
G[89]<=2560'd84861676924448135477847698291933182969270109803559838263045818748479236104726770822156305517351321399152115381979039071787818598716118036135860369432465581798590108041026950802983592206926472677439521630309520808261520071964376876911173288838687824944292629663348023916598181663572056578293027286618106951985009644686038524100352294176314053080020437289159049437202541760441256743419125942677251318766454387953219030481403938808193893231465291978346670562009458062889225045766021703107876705393757635746182560538931793843005228315976760083046245520245688136632736542795252716739877679042209407899160438100649596451131403614287530317799995497836201197236581716823302975687026684611433470991825217419400763670120268007613444667507280889933167337023231189938669135715246626;
G[90]<=2560'd86660042054959186203317939881611136941187102524061743979684747305773603167949495082644218922157711575560708848268936227525968118935853211591921765680522137127820191149260207795389301406102020765633560123579243131498054351599170872984982647133513671634994692496740942454551662383337005529259762188189428878733662351435927880904894491560768552910911077507245816215113903432823048028335002012073412211247661151115357362557463804325973154012584687808645567279304741995775227059555612806569008844297274835442906291339343233052935512409877553532908582661020426893385277100762246654990829730243971258313374494390963976530657440076915392840845353560166659051761954419659216317579997726507014517839770197533900893059799519517117352681975597983690176737590772570711961795542786594;
G[91]<=2560'd86660042054985355860247144593193911341744314216542566567950625121514417320961545265830318831687035717921868537533708417470728628786172960835502560281150536811444322540321021624666280051158458527180083217040739972660683108646960734907174923438148809545509677057276475702326359921351356199716725897151800162569169902370034466580230268157191342897385056504582572198246638448441186085716310377152958640164700717121756407490338294946028988439924829548227277968666131301732078578232716388893368676572081268070892626593236852197383331223659582145924537383369215742952515268592973027742739965130823578369112589455882708724300530157063840593092846101088815575743137382783217277523949194824053843845730150941402027345955312396276242237790622227435788695200035768146667033872966178;
G[92]<=2560'd86660016228280241319705402358421350846742624107826118090937600629889003240141592941162634795809343845528595331948796376943280420059426728206225174983166026905954686969162301194931984869673934189588887336905977389447092857165515241705355888283109705347201233459613142005234012111974625599800771935083018002123941718459699998266559529779508543363828271916113812101992832598629957006715952383584774838566653855239296431294017539641105107417733543686412616418419657852779948152548770559799918658169235178764477808228146216818404018453660976131859432179900400456578002928432350073360801616209158185917082734048162681880639888469794787407731354453407252586086727000973075537746408607452424218360384551034471733566894734598966735313839546562530318185257352449484080428085289506;
G[93]<=2560'd59578365685520599527273209317268622070023453496135301177712986741341635673315141329042546278281588768226098689829256776952615299307373508319916431841088991861144884173920347275376591421642204513020731678329283323221134071872424550292060929125372273267239702001936393372232647442856865232732765958910024114724472843946724781073806920839557672830789699016533482169753115315835209410612555125427000915491568577291642802689898551384399112316736957662725821295865502386187508126826164420645561268783450306164099719291958171799979606633617462295216496813388461092598371906806125364472475770339535660341482661053731183081535575920465665746474223306474539741593848911353187558683653706304025041275219738960818756059694581554894703821979093868508043513628273768991527753050366498;
G[94]<=2560'd86653017184888847290607888860499116793301171011115448878627326734944596382599360131154941098967256317572945405638916113787806658507003343093032328610616243448175383590008784736674063062260771023140080532921183005235204347546320093412526250817370916490706489617900013663756741393982631401145874969955265691100697120391588651330718894869146150013699458939426576023837200578906138315525658080824218783059187077161043787456555229386529967448690631820918935253969924059486428940451687701725801934650259781560239744850315891204149294072157890623000546076020047442194170418033780199771495187730610911877115354789131579341469612130844786735220898547578744788951644320964256280188496879862710150821150183461613478586644227222815101456164501086837114136727300607356577347715342882;
G[95]<=2560'd86659628720512608453045997684268877554522436981137869990667778812834812671990664026512525963115700693400811458189923472768706489557104427707402848609635841029425622463354536924521054296828991062482676161379132402879075677623032776554689312060158055139305563396112543200348763700148975881292317137530077161554189469703575559170716972233934984998697908194612401563791075240431997702475321301617185051026974853497646358475438755762195631832201452267395487868782499796783576469437949165569391200489816803188434802137749133069211919741905418911266779575252159184047164775143732502543585929199976812200921575227889429623038538995561017013085720341203093600090225424262375739852575911017191455972907889320594018087406242507336228512974393853483183390029587583615565381687714338;
G[96]<=2560'd86554255971695601011258355623550115364785881895015729348477658261898988411763988058637255489790982563613273956254331608139476278349510695770746689239347307618022661182628740546318887950301788824771317138845423899527055407587740849250083501484625924489266259783071681167449671385959350429745684401329007963736056393556726724101413122411046683442012798464578771725889699809230426554142833133214217107252521314311918868145202167897835391539087267255167943154327172425148817525478299898584580066472738745151499381542318984991769318752527496618427325684601428323230675844822729984438812183347592621683373668246103882097021567910590170553539430679608862796861308746760936053963077365633309556338659268101057225217495611108216923909852090782490363361767496932859521981183304226;
G[97]<=2560'd86660042054959089991343935452503082992633242714398516883236922238997404852538955170768457869218011904834296788013324429273835373608776368953183717752638611392570234202549305848950797717692103387002492062145905723612861405436213919331624853227279001957876648458355649569849052600300714591545060117703648050020246347024814307544168478890979180428323929429202121562570654383892453506373338984264886044242753929183119484302479588674448721388673533382845160526611651236676778340592308594635662160448558304346470871774448062703799092567747718426319009338879306402555268148507359935035683745707580599046153149406325664180690538714384669431464263015129298979973112329470975255037595338111921181702755480919040356647032898303649266883992788258334668134784009662703216373822267938;
G[98]<=2560'd86660042054985355860247144598662928879503580519033858783424721397849499394200573087902534590125983009847885761199052743295786339410417145675947540670243424242185952893270762379425394223483331080337189350036778009575737659908474964089485145433064572712596553730591948375610023845093177914322936561740607913937958735409093987506730441751977527607300103560388349276401902118840081762375453360306113510550146578114423501712442751418917663555626932137353268358423297720792177136873542088617386465465439153023748140473945575311741387654916899680047246097623242789369383357766387040019028839612770575432249383738009892279308207807088873664450993990458888575161127945598983734601670023527837058119380385053655517705650734292308761150439133658551746105854185752914479152994853410;
G[99]<=2560'd86653017191194201232210530174020461615203946404805797402533605310811939325157651693098787039480532549375788446475899353142381063423834360829199483618737578742541979314957495021829235079925972558337686545952528725938401361992147402712017124918834262108385591353660303719483910705017777204887315741330100688627237945688881412149872996970343528222642707010805156132549640847476471890904934223358144403706119496791581715235355450151847364976407440159304802837961197452866409286860418363892000055663038445041327365655658590325571210534058728856125155725464528191427368468976265769829079406437035290936930508516651530877887575592043384621279585196499857018279015857039914752668370608302453899953697656397868065731280477296501686527073383456831151763245751387784426228556112418;
G[100]<=2560'd86653017191192661840626459308311537912492706353412262357849455382068952953697780132022856653801649120043014571473403339171948002318821178269118549736120031837358567315355481062664417623211795413611096659665244752267972530565984769631503924363184121228946517893202331780989908891838015149519190495491028261356651461485254097920064522046720481928872962622347284658797788827658375021590480610706555264513413934185699097295949741837295619558996490596403578334055340826405636650644245273842169050370932257502893749601966591563287922162088861973297830694097403655533653116513208966966266673664361158342693836676240404968647055194343413622931970947674405034503149247014012015607215324512336630374400578714310473500205013675649019033402591413284572013763519485397683984287277602;
G[101]<=2560'd59578778811915325908667584546007890152358405855393846154784101779059989466134168259530490133310863774475876248812450915130807339204008662063689826795174012548144582730092188068532659159010534020584039903446983714115523233876630797950085894409990532388987045342331138301824437462988099477234635280526431012834845898710065423546597152184126203525578595925025084729733561182611142715531025533638564068108751050132720577449616778808388993527916624910260097370490084071896726556272756119598436685178111939150513142448236610593263727916515285746153840820852407698059891120456175355516044856171229960421387935614101499970216269585457679510100513187480237621743364944926118638611963394320420594470864319049938650290071802680836435134106880147402641740237714439110970084685914658;
G[102]<=2560'd86660042054985355860247144599026105825370384862450713255366273309419531191671743777336545199199408972725121974067476787700932975915065310524634828185683019126850163311716577502326292494484635010015900944924282130622881883621451827640108219965661238684472495541569757446724817199708381302007678694941517379080823111704591075533418962211249851759250050413312004412204739137369688113956110401132480439661814035239509982133098146557014421426285618318058757427798596153002142793967094515071334475726070289968872588220601961592397108144280646509139759661504920612444035061718528461316160634404294258466099383454243151622385750925755239389396975227594161822293703202295043652868560682000645453040482165820066472421188353893980850152776028839101429313862860660045321541483897378;
G[103]<=2560'd86660042048680001542816121418274708133087735184218121714069309759070684200095528121131151229452618358424989144651244781249476201811325365763530691932360645948103441515413521526728724006714559851654784886348550217802339615546860490514727621003143368788581636201118420867407436792199238362886228157986302182827080889075070645751435640161008633004408806350119647167105101498606748311932226981893215389172688014645343007489325076417050892857209974073944895466807307814604156691105462408997701234236737923122557960891269118741313208623225968015517444427758015495407698015006754716656021007762071449482254245082819796025270672055588843838538620828806404688254174734602305173282201385031777930139348055970663055009810853620039501204547464719938955003477396050364228665432220194;
G[104]<=2560'd86660042054959186203317938481542736267124884929639370484879984008043132456172039682362200766207408574768244696095950217132994987792930293934877870418460833334887952689849087911095144844313777692529905864144415173086656085900327319089863740628222005189876886593675861025152301236300660471035028733498511063880233198761014139936520369798488425025931435221539193303349600462825359605337210880813865978179291685474045957611616411357425306730600387998899305227268075185348462181203705843465830126195284058407379190726369827952788953024668117839489272193540056126597941427784943117147830692833458468447883896467653342544537443070753418354343307170059629087988548003225023167070034424771222586410154011229506311120458614732775307837512381298122729102398736791154365380430012962;
G[105]<=2560'd86660042054985355860247144511520490011867604514986038521419627616166279205998182444861697463998358987853822776346843716112966914068847527346711602336585650717021411204835058777422320613287044925775558102739449877344826082577461742403712360128792639411979967174097852838403878490162384444630161525433676190145748292759542130805183788202814811640644751386953822749611260339977587171433683657436848873607521968768212346233653630822299217509479698169389854718687967384990157695105436037482218880949523542517806967156147050792742821483428334333566006508740169820700299407259315342604161447204505678566524499399286052508665064300973543077745718861877109193534529427765238381215709181802816473262897572959013813020954393270940816365081118121950606729131567706613616775853646370;
G[106]<=2560'd86660042054985355860247144593557088287611448867467492972011139694382357828526350881001422170328006352946738808627560341695352712217056082743129523426239495646348954592534136047416940292394810966226944843910833082683719317595857959901873693888897743886138824196926248342336633766899924865600486164442885449447300906959871761282120926102471798935511581371338443943374366339526674239587952813771423364698580963804213893549215754259347611721358770159825216063359056289493405253002437725128695941331026914240696192626889362767578392361557854683832419575809849010247301505483211969821673091405736086086811363951491129084549438962408628828612549361200691474582804402101596615077354176217779556033851432332009150115532801112221949271480306913700282778692679671777184889855681058;
G[107]<=2560'd86660042054985355860149655029953662886182500934189443562636301197143168485863342094738312080577243707953319893851588370792543370896574288963778115362270111613104282780710662141662175277559670548220191001411061928826163549123890050219712215268113219249049338071899793709974529922831131397469497749812697172054011149298335215279219503495837453231779150556466346203330093031023115862152924326385040606839801045191168797604254064189368559285212928647125886778757249984540128882575117932759243638195414328220129489401500599157698550722830622501728379287075279466730727995444278653312720139734792903997778363838953820261893592952803279252068722217568152271082894028593448730176774764925385809594671070282952157685388532386901578693920989386388355835850492758228298886132408866;
G[108]<=2560'd86660042054985259648273140169576149288481194431819015847103641316569059641215220702362129782350109669493742038905000801475775709483047968337069889665645636944751692851290677633497665775433706884580705425282207594267431225282320244883944801926958973506066443549392951552627029226967725579864037963109740410041735477779833157382391125514000711591725611911312906567241983597929653572179751054629738722084263672815253561543185532775740958628031336433681167157154421222213990970218797697194999248996494664514312945704825059369961568444134068394197570948233634203295397124341005163567029753198056193068728164510818635906955956718784123108507576766126019739906220105454558527787161053273248408900649022856057556793379442534924607255616598268536428255186569163133413974964576802;
G[109]<=2560'd86660042048680007931892877167360035653590610219408801888781839470541455566530072215186891493202050526535771182328503469000137235623913785574785169198965657953772138912855960449712120749846141733254927193518388407496012896947179628370234422669510361514178400579162703788940705286130801676298969509223236336847741999000163857317101768886140422389830559597136122457008639837160443934779853530137629836952005045198492666000392972738611740322960762387517230017218372805588431735696918271539267615503864178745721401607153120632386538856886345165992421141223015367955287607552600250679022664702166413688637731381294383336787141054637561676640577697201927562794878536578717713920298167668901896017062109286309047986737412120546095049400008232282265371596365099094710878013104674;
G[110]<=2560'd86660042054985355860247144599026105825449969542042632900029040998767072996059537952825393853687438563572255287907575485204458632165722500920842950802891374851772188166789829351591980014605638761421073032903080545541221407846875526056032049725738737927244409384568671261920670145435585640240253188736583699751528880983018681111693295156334520824849539907372779097521069498167054050948896250245492345191193514781560899231580673466836999595691539932145062192460568996851347982531443843902142459934669598500083793064663776610380829334275325463263551744165133078250964085072759162453009517008301091162117295875426300036911330233099698822087795186186756620453160391018498884376066473869381327403244207714809492948438488864934676175203993466672912197177669432509622892288418338;
G[111]<=2560'd86660042054985355860247144599026105825370715169958785187485252827799513318616949843969036653445638009022658368127969488863849987060137110702632434979307481492750888855974708281754858838279804618251520675084606124895045954479128287542543038216971282259545365902713489298011898136466020442714708925480911854474090388666856504964830000319452754869868837157424790006811865061859698121088961898519431503591286158106619232335949190574690605329483988937210840765463289156612266785879394128233309721677375104951032709453067189446590770894774869595893919269174824783387669179833748744325171608616549982554356617239250560300869160768813901391099880894952423646814236614301286607185781037676231300085429339317575399960139638454523524275198108493958985982151905223976366098492826146;
G[112]<=2560'd86660042054985355860247144599367919767832843946171458095363025144077893243547024673449360351809036885693006612255235701566186274850062756499714903464555666165837152970315673862821952288076905299595613667904778301205242335603976633875723371832484063146016433785842795064582190278057390199433837457521431972145197105389225393360197865308621339260531420861479117582290387894461454079392704008343925065748675050357862400898419413197845770929883998869396431202819396210363087703912996708288475019858759358357047058089411001255276579302581779026123515133313146381135177113074954854881822027706537047037536784672099765615233140140823180083210151529521766057349722520232493200135444763853807248124338142996266980924782601585033173166891709508072445751301374857300283563555562018;
G[113]<=2560'd86660042054985355860247144599026105826643739735921427569970269842902000185521934048317661086999095032192201833219546841405520278883887019582620768009236225959138367883592383347371593894760616255043437717480859755538593623906728298910492955964469527231365793684824784097312859347236756897726447547728272808106066423339547051918635098208980300760674930792778958187749088552027071520913767598509323781076256133884950321038343820122811803400552877513319402679712834864750181794462746365575970846207888555018278017151934135962601242635468845186206442850294446029782053421695447740062537678429051960751064500906909043890120472965540885941065620181624474772108502900803553047892327363501432631159307814561002219543610517633020437984613122989523966273342738807423982462673494562;
G[114]<=2560'd86660042054985355860247144599027524486588532016285764563985693930815780328138483249004206233050550659715898373886167124141832286160382210721927056250738607463729644045743511560742508903048220714172606173248847285115053645080855632482672533320646499540818886538288242355795749940509451185564184306643254580034780634827659370031089608987902660556922222157529951372474179196628126875546238316090085579471417882279012347266908165577908824872482364654497769293718926668378041175873291619863724568460881024041910823267518732284757385798552823279366718023973528140412565421073228744886959552310450725587228736782404686131141091603058648765715883553863883339517082597420459400646491105977567570352064211946972081320874608130445212959366263933772898374987333676049591850032570914;
G[115]<=2560'd86660042054985355860247144599027524486588531940387899657751309501893366630135617390547343470120377761445114141634442734379059990044064539289717787377506791370020954896260205584371090902488264762380955303516197732110070885681407178664832855712215546060350917919679041623129491692972266705213906356968667707927035252977300629708535915536776158851839669203110519966577729673930017807822328379860242206080242104430480983589748363730236270170713604184596920866693026098577230543810151331924740847167974060675886281995349529091501703299143404520530202168657822016840752413460173096150000995212878850719847692500850713708036266777697174051157340668518253028176215393420207255945846475930001425944259374039909758376244823544846271404092035967073777436773764768041958046810907170;
G[116]<=2560'd86660041954099789006578888098933835296901794869035775644270027082613954455392817303224710228263435492372239252497955172355130544379350719027006475636466526568620350637704022331144130887686662274145434226396951093172673534404446270879603451253506579460307505189056805207656279358528748417355080339749167857661818143667432844753424608667333620700346983167693600473285858962800151628337315448495189657188748443913796555553748690556744602543788809302522703315691136075828114234997270948761866883675907824574367915254772794593608661549459276362005186383653679467419594333066437927003847171883774427195759979581140368264587794166670893335128175356958638482308304241775664293961961587381220928670097858300635297755801110751714208566491294812365774512155811706486439226703487522;
G[117]<=2560'd86660042054985355860247144599367919769106529127150244342086001252994799012313212040176904645517326300018668991249838261928952505927735771224395760515003232941548297047653415932373474608124499147973475735143570649032690355234309605787969229606851140159781672913310161434433219760216905545230988565867588860964608018171597659211825151006878270333292826235603051246289946152468047226165932311285825641096830454856317813670492288966748803204430017048331066223807330981288010569487853194440345980425113551846700366199056171099088884822708579879692824125872664749636503936954823881858444725873789922168573998850175725670616346123226272308584248784774969460242609663442670650418144971938727060666847252930268783594398380184908367471094754785516980922697016165737697180771295778;
G[118]<=2560'd86660042155870922713915401099481642334036776174672583319018551416281300785033322120845453309270226465453160066596391513175548324475011625645673796497836810889695522576197054892788741794835222128143187760893181968123035025762556039571244575052163527021991789300858394324569172477241044319547513957882326529721850394738191152904886245715782041882993590149462192002413637428428981514796625538456107021050150024995832448621011471989257583161997538341527297766914539021336016574319003607120220145646797882843869255930184998185200180916036050436928040023216595874049420667582241793246197422422805304752796554591009973692031937532575876078502953144306951235647094479235845393489979814518650175311554506203248932848239565914785919035998302042981440718203176011776309701738897954;
G[119]<=2560'd86660042054985355860247144692364005135182539367195325444837164972273252261691372469817044057153640167439820893706339872661740617280549667106311944414980594193860448350187273514201884819403444570890780633275883322795859333121382760445387664718666558457943456029184633292647643781847512898889272535860729031913406575399085962951373175634456856448312367540881030052220993510222913557356293923621090326233356288919628502380266659795741991037643228882748137006950057873481796904403741300662815952167686996950811515698611546738302997171491802678017953343756565290985327707162190775807992225616356909405387991903514379920476386843087074926648297798580189995610895322411076474298398610925820805994371244181063032357106511764672750501310567478284587630167951433109767227692950050;
G[120]<=2560'd86660042054985355860247144604837025973196573356997563505555995059054939655459262649553745598831829568815277855397816544853095509416692489340062557487657352795028502477719666141954325284289825104303939820350239211206257681497981396223654889801442790898054577111210148902036456581949690801315309597925973795972818018983383339561155985028735182783822906579365585953835428793794644316486848410797909351105048266540062450073280243625015858982726015525328202907228094203150188328101427052380964895199495358952500124174313925564789822835444744391046476300038085081704737390767567132639569571910351441392237238605524455157943599693080798386848947172293316915646525751810722467869000881259724222195758772312373404184501758458775902260990952067292652138367008552056165117116686882;
G[121]<=2560'd113741305298053846421710712008767970354745252404148715328724415064242331614472287194116343533969700289096027230559528469149699554797668871602668277050004692586659637119633323923913104868157245633923963926395585119284553876542601337829353807167593140858965326538523587290223695877601920824970736218146014986893074729774893458663231752165467044494590882104266211146289676383903601937870102914352411642778456664079711765794502648165374758050398902335948105012104363108382681111463441044968080785449707312022361222496758784110446591736045021100967454427516735975940070774558331598679419026020224851561316474340455563919418983211555891526251498301729623951495103907103479966641181020661147884977181142160498176036955168184514459219681548845057620095849993290770917148695077410;
G[122]<=2560'd86660042061290703788601410636115491441695476270755969252378915257856653451976972113415319561529066905838571460457347265081034390201220655212173602862834683160113290360097209085955071294266057458932308982146310517199981441961929512779565312477989876227220098137125495487715490323954349907881287271635805469695503205226302911087158240264608616069376871267984017044465891003704237086725238095924078186527011552052644807351446727613218254227440472572387346737444698387063056542531425887045565206935235251741113363022636705523631022726226541431865455489884075355638866559611977044844974175911792161110749790574640526205765794680537423869633984135615236130660214126718758663205850933437104776995797916059590122989079827415510065044796314882963574513446247468675821236226499106;
G[123]<=2560'd59578778919107780082274201744615140160397745172935098203477919818923773953242782976623279258701979343768690115810812085746252791997164132388125526186779552262369312319257174289758137460348890681451681460955083097770147474257417425356025183691664637633085303598279517098726502698156505088320621480214538595982808944386012260854218781747590395561568311737102566462926326650216614260718458292204319399015355833117400409031196763806723825526636459393128787900536479841698414827049111518095635280593750729754219035279817809417491299681530561482036396026916917833841027027073794130515834337237042504564561311804425862904728167159447458518711203348652062992155598532312010724537809142586060849468819166521053567407645815063447390755822749610553033815010850298792864882670838306;
G[124]<=2560'd86772853203811229389245804881130417010254597758788168857200471096070390314800883340225316918822798947746347097220297314828869191408941793082022345259215277952079414153396286495222524283284728145265147281897431930338871540673741831370017256246362922932422981755389124879145874738843831916972943542586411246631862222196266219432306749666134087286424009862219602628367944637451943512405894761028094244961339666761607817225623271115776182533331900889770928963277835053808222028905479115329040388454943053524944432082425475679390220339404543166149480145323384211072335638783123297155401016651642992317761924518566895376915103867076264689408407953119439153009639821777428016539331711031053604917547479080880539801453526034441946945897426008666626292905790328026746150224798242;
G[125]<=2560'd115433884244440279176937170400711191292356436975518537097881303842390378790409998643517129098388973155256510335016879380647050606856756765720848911674684054150323434897489794670760665391277158602714941753015345634602982401952630386307537774198923942593259242840533039116840001333871331191856196538414014994304869048490457933371719123108295037190284648314329534429483337029594426024667051607903736596789801902350551651942745657911173803641822362601934660092059218976345614678689780866078844526118301851294372802825975431394384510396611235952637159813865738013960573397490894246123287241866579149424621121261208684312362362663160649250500802399865151479999128315337393853047617986496981917891123487082346203092337891113711449687672489593104517604119043682982172216451539490;
G[126]<=2560'd113741305197168279967359731916973413779272986003492927569896550740855482233812019528424827075622775610627851703025298144945068876407012248025808241980366279615944945617629855812170409669093839708884499870834994382676743210436662037520526338255085354363405868788596931428270585739746284556382511524379399509244718871352857235511288433807758515121888255614272860302903658215219253262896657603363159615288181934034132093387283553548770628678457632495345340235650230401495022252418643003224470815184347139077620065321837851943850926849454805815985434837997664452013201714062739625251900050270846503472323544813236649119420296512747207717687977118714725354886407337202825318481530526710719469681929557883124417394910130111087245668954961859549301874279537412200652037196751394;
G[127]<=2560'd86660482723141475309297140233402764849692836794158596186454115562150212685474971031912421787266663386950366732321538638630257769609627608015294412688120031701120034078707920893616087423798130862153958782341505432162885169250074828622206170083854900732324754875389598212084646792231308449813508682673396390748010550854804148082585111119449762875760228650391513726903299737148156639682133456985992087183292323007132370951955452951710585589038591407523822744622947652613961892973314465715796097064015714829547757099240136924315123495707676917362491285392673590704803249183762801688828181762326088986153493229194896840890463418013193946967295886138375931331463820086115688278540616536491498941953042259646507306220794268836403940781381792371709259396364459358889629540557346;
G[128]<=2560'd115433911691621446906621395344017774961608208765451948053988993542650720250031613364401252964871524442026342088693393035769071569242367343578106295586235676889843881374348681781564057982459406761779600439617628914904761416378132256935577688786411232409205294132588705820970248554102715505741044716572170166676624021605965909385058155489092254929566485546898139591242406065247266458449458763966424003700964792845753058184305456126091522180902349113961366758117778784239144470616150499364602789405338374118255948969260192924527777963823239282757345998535075058488483284034201054714739694338948843999334221524307627167772792372906767144330067493914141259296332069663754758245901298865406619233261725011878112607591686573951605150462756202402559805579234939802419734390120994;
G[129]<=2560'd86667092752207329484268638659699181250365130447820249983240489235938442052831601787983170352992237439836281018561242354846613385475545235504291821715352063122794224334257840738706457750233346302420122211054916083966887150171054697675424597500969651227941423855771768723154740040800290464006899810167422050277862484334478863226749798903525149159890752170683523375631149738953204817151606216150861582741416996261565299059815460614861367487794579722218086775824748002791772668651553778609550561757776760076640485407908212854085597976304638770419339010486342981305196226627951500875695427539080828687979308342679784535099462324506166414027631491267596360718405080808516165227731494249102768164153839924835540441475120656765499550547619882384737702346095881907666912326853154;
G[130]<=2560'd86772880651411118042259351832475164532032683832564565061173956304049869666511996078968543581134623465552832493001978093005390270560322586470451359310195249263172250582204868804701001371970468172891981426705690516066218060322139556458531670334158838000433741854986962436935200216767112597972921293183002961395743636452976506026980830718629412992011730618645807106734829039927435705033464632686320292804049929222549097652634924775763582689208856616071612836847145388775024346518124498072990781797024133432066585619675932761487288163380762642222172384276830197285667251854382803112546460433596729429686748048661943945763371192450535851817184164271777988513861430259552463610262736984709733738568740384777589484674837524266300678282802013798352334242254644108420304729154082;
G[131]<=2560'd115546722739980474480329526132057506326277188345202266293755563842614159020927418680845197180062235791576021463593660129469011825514441245747089045666831211795960504335549507766243687520403245963576653544956609720926634598360970211122331501928646137652111217839191671267080543628065778200394950378389071850839575328682537111388413421185695724670482829414605879050867715204622891582489057247351695482059784898475748030614464427667306359894568426382746677688112783654775417653766583321056503391116819219280675168650242571582913234640538358988182090954304055144867991012468518145079815979493146203720798819422948516628292656580594363313728024326604355419072318257622206048932748429706017416535341741934653080673367759515394200981211271722801369122577493037209155624105026082;
G[132]<=2560'd115546722840866041333997782632127078337649813967881559016773917877172545129559538400798818464379668576302661976516942306887767255159740657362400006406752161676358929933714450591660537091731539178817187021354497217260589605031265792445370006549610426756707469627246754091542081044312786293729645214925485686744949978415725257788770678217772773498950120966008653418527439917151797356158777889879121812486266188723249314833929041956330968301653842981966226173116298613113463952802367001954201722720855248471136159923051720904736768362648632308698262234803096274547531889256026888368694665846988146003530557398107652974765966318390520739252724813206918563476554650769668811584980222714646524558156297397302405539673745925195412868312734643717129648379455373060604512713187874;
G[133]<=2560'd117351699614610380288105473133013189704692727879975928932222075548945054987405629429136505774746338813056740161810019409871451359444624269190030622841573473994408515580004065317066159093295121006714438356789683402104803335366031064758180726473368066568444401761163577988965137727960206632933460183916592604449402275538647672487240957292070276152299457615914370501891211066229076429493458994393050821527857657209681790520307122023835358565780137390934776702556808396708358832922520325392585623776998494330264889350711077984951248442161603061622296773178961564548224294917518988824812475400671858893181540012511869083357637302587370108326113180403223092810130390425925080953210741849778358802893380376433240628983187632886434175917923653422861457772203163917654457948713506;
G[134]<=2560'd117352140276485679448040733356479861990426169536341598417618089476803698312274472108315541076051599581071171979968801940535183886808921791274480844008146703941978261152120235079846892882849952995429204175860118508455469948999936388350138819466063198268842250217370630383510282827238019705584060836429994359389096370141332769470159339326782914799993614251068421652879874344714854444338965353174802782566946849361829803626410338958040194302572562832902749697870609171826878614123976630867756911130494439689447998774678105550468204744179247204754364712622413027524340277922181804355880278238283335382771488042702166334777600502811498477797057411676855673234210913043627388294444652409610197423088155122053262794076442771685714984584442347312115024328639214054105621723226658;
G[135]<=2560'd115546724455455467521240720710147800655802196337676080328353206644191505466327218465292872810270508441029784160794638820969080852602877580923045270127255394613301755484311866723554696374622863923442264187057695011698286253892656056665536029939086349010191250566925309910022475789088755076343184091991088911081378924299810069586132289976111124981834114783571751899892802698469284828771524554937245118168217406821491564557615224658983120697708266968305168915525210490429943877826782489908108396319860995890810591972454299079645872055500695623566425706571022481689071865446262062857938829353348834178717790000782353888672653087321119261018405788922419387545188305557605496731993706447018690588204122841681295646005561875357572195776740975523265705178156756596446807279673890;
G[136]<=2560'd142628013430228503557081281218266479248212585769069144996683399245633662009596153772531916030154576050128715012382456842804735875577673674647149933444654388113354839339139602023687371982197939371199692097807650005123145747004004517161280097320387272558661224857750406343579106230107996745111220541296640508292004224008323160059589542606909462286967157117787201018125083934675997892051208732559938985109693359661822947860225571866937791727847720462857313390376491469228979688916558800366996940940041135414543890393789379379966242121555458530947618412308587318639494004996561259067052364607422023200924788975499021425647457784724348425777532187566093398822154305703844025217124042433252892525901662212779663543573936083099188802566226906654570203425719446124392000279159330;
G[137]<=2560'd142635038193554435080293935748684852685847368530203091056651966548940930371522730987522414312495251543955545980189530084710889258158098186243101934465013747983003364790447873387171773742648055933569980590461910492750556206941039327256712154666548845145759980239390569297427810037669098969129737377283362117480836753025514747428480371310242110307824603619230550145513333629118307423111640475319872035848943357384870893575627435436996299676683331238898043009918149744751003849227640833649163710448087805604974936095031511705213285632113165169763809048567542174404129447983755415975363259421935564022864018240503855095642401847085030314201446357075797900724272206727264968236092442285892589058590597386995366132330093160190085026290389888811059833445338308552656129227891234;
G[138]<=2560'd115553775051371517763048858957117660329690701752383389290083229214383843940670454416209368991877340973677102966579354923785116915690634065938696359541695609614053679807310959049691159235641335581081516482014820772295013425867742164125207122599747794282909184287520215583740993401366738901779501873703511149006307482413402106486008199178220130565032900379045038303019257279005814742000938934449341493750956569507301859779978346245520678026998739959749471741813863161264782904889133880132317154404787779167225716681502040734360580893992226465847674301206701209168537805800085148894748476662525924092983677301665216596238911694991845835915416651995443142724016700790055277810425065300988725616754988868343812156051437783329559285346994116855742517059496953850404729444770338;
G[139]<=2560'd142628013430254769472969110277928960657550910781411454645039951286106835109283106402469208982902919445754651827411248917198645566871629913884413988758740147722341170277961446331826121508737146806256666969088445203328897580932315784610115090570871824948192283375904537155509869995879153717881545989864945220983051313025586932921515338106175431146823539198494939542561743896561461289872648478478668557234321798261431005339514515641121863736922557685077166312179289876883858178663698574484247514787791748971183610736670009785049317862917820694878678125647977169299206250904107495977412376361554884174283801445368347036386253221614234959387141138220818111402541967389739678988914251763595084670168928855069132786403424727479790915921023487145171388779644260979670825169986082;
G[140]<=2560'd142627987603943738780099954543001557318226344960567346187235201862915381733807021941129528526297681605008410310971896306709923603008144289579932726074624877094322157815495792637110223994870840106107717000684795023636685299938423635826476073953993240725659643662708844197250824230861065775916338202709556162270971450966628582725558755653684853976322460246565384245835479017993025945287579423660793460056141766315847264154235417713825088079776740716189768167485310783076603786798438895972345934197024174768606278065854435195540952023472369719500081956490525275051722801899978451524056539760352323009975839387132729393564500236721527030227165175374804780111977621792256588868585050412050997080671858416190375072061896989049803551771976912763055476231702277591011036907053602;
G[141]<=2560'd115659148109124404037260598551147118601660598798483816134459947692508200326127097906668682319332541041387484196040097036121904001914479629116902993191775129330855201056774544065991921708423220504325278042099440735385595664592917688580456513388967881893713270907456891585637433577300365244146840720679577774504185407995048945599106167271307022024311863292763891084087795541677893010430751618665319508549552857105357902449992028539209428827396575003971729081626415891459451989985781575081270324215447883680474784142604034815695903331100628763360040474474597064828522832032598767019332075960156749551622151270457479142553031667607736260604084098413001857410811319419279776999155234226714278057952815800907823159049271852117699860290262864668334677585660431231110525550207522;
G[142]<=2560'd142740411245001979815233565212556027300465553640055745462782506843734964415186668376160815387863343418996413166431124869196622947314954016579837333787927166508124849341924668407599581220724197724023885593880850453100037898326815409020893954430923208104974045849916021825548143337023452015414703737642266451859670066509774153437402010568519732997659313285250746247174718040331185894760221857675531183179175502279158795175781148356802050683265159799988300125006053538116642348949330715867594291780169046815739132599489056171153243865915250247337883716998698114173847200663739410836294503894916581211045945091008790415431952997657112608333402257216246718333230017271743426190831908513758712201625203197364911572643296273831965553756169996610573221166072427095322518718915106;
G[143]<=2560'd142627987597638295391428446438176309383278691266693932275307565595716775136285768568741656110877034396084807908772510960130722768598234674215845331095969161552454130315744264760991676535610767522951783300212116686524003308133854499104828556563596912031169447347891561831504608052647423658701319451788346577918566359423336681542342034811663295019312863543876568834878374961397125066250512290896270307435573271362574724475747347813315368087864605989176192644892484177495857529157266394812677937399756628172094548028128388618840513943535913515530164252978228951480285133378589137627423250364552286622276006948445145839834298748959730445752932177105625909258912474927993237231921030251543341029987137603724660585331185986211462511189959966852396338048909061508025225538839074;
G[144]<=2560'd115546722847567115525661377850616914447663394563205472629566092856299003202915213009757342730339919271177687263183000497937250624568849295917183811229700509152715928629853557839167999028869986508737944555430973443121632877605046029980268921999267336237824541655979308609370347905517048157395015933999250207324863165408496718794754605248066229821203350160693794617157702057052602386195312301300928101708307801435910159336337561750032274812433220864413900293202934289840531027115250766702237631645906479367556583140316263875701824548671152854896747839279929259148648195153754777977395407714506278144582173596293752627354067025942025169123632066457295638342645085187549398308883636717166896366559512895849896271987832022931640371416237395358607173718835255609002577776227106;
G[145]<=2560'd144432964370988645936159619263482075605760031238280361861418489931734852553236449532135629081054743224715288152824884696475471025700104903823109319768893938684659427217211739444673980624638028490846764708572083568051553465974529923877002921719506562168009036555845340473344530211886005933180960297465594637089537575038594914653794479802340639834699253501476544695349613552527700085163875107753768048139083766380086130712356710640207537361960538249761135780687649357426737420161181660823928405107859413305531022296726611956163059176250763426322526554544745991920033014969886585757788959009809774584937996151143775843125885229017446224847505452002108410435993909804378218237498675472396237755514439162655853782068390420398331391513166507349515584113804524386569125288358690;
G[146]<=2560'd142627985888889102667148982273700462262924626197768430604900726135317488750968787611644443538881067636467688672046236397284922794569128138138528833043461479873888628375716529170742651963184267613939868209741942167674524110576038800352168942556479446777977832806498623004115814094054675359093416855151052817523869107272045804992893528486569841664767923154942481599879629827721336490908424463408319704465532803489722872638113711774995787499672642974628554464607847172543513423838978047665723126669143413621464474192912826376635617836234971399975416222838142676167328833867432106558111672636290126818425003693412015378026302880040071808069875785541202643457722696644175901805301228701704068075153678579535285442486586966397814238011475839134239358413230031924896210438201890;
G[147]<=2560'd115546722740400831010446310305944279254712553084346319214516267948232084959092997415696405733798435090907681704829284539214124160690450380250840407037892905608644569992501082650269571136101706010243523546897573036014513036226951616744795705854807621837236088159902874976416218794284556544107089764666053265445900033516409903615592146712406084248387962754011667702141118550566038865332562031838417636669667468621849160744647065566320340982122654148271971732787716540158447355968891674314768810845116813949774771898333999151395537925500675396523785086284363405100309478898929151095334030453332628208640242351749467028022704907771259814196349714782032463224240767961848367849327121428755488758523832075800727896884949386101282311395437793587903265790213664903257482593509923;
G[148]<=2560'd142627985882165040180857182943417696795404570648039823193039361563476295469117443158015965380570117786922091451964078313216705624027017057434102556528493999935530264173928891627038446436224898131306422280989380617028638091787270609610660868701040669620638628288627723365047875445084830562662658324496110665229551476398507595427626740266675649947849538742934195359690124450666715123000031210060170582902610821187361064292325189243423670055085585305583640601446876236798340845553996462346072614826299817860765579212854302806396950096333700996737733549066875057239999655661214488400999294561032346215634513780840923726015477368160736197853618780935557504107397647347094246316696374631720143879162643325545170954333751869279998476821955834628592354598376361783104145626178083;
G[149]<=2560'd142627985882165040179389104726797379573142758223675460181216702640107990090019787053360370948824196462846226945482515589157747772761876442398644189793869841064509865668507169576714796987654634815609092504922428178341527166850025139266334746159830405982810652065557306506486849569543116606659385081364252824116836575450455057324989401497587360339793803750829022513325685717399757769088664700258743955858851306862242368317885751106804410205992483058064136615534973961291152764329925777800729852496260068430145295529293674263848953573122177344916299587301356879482706167439967280362374443968444971336063227810251141094300763334685075111301255920350819152287440183063197862984884068186974973199726292693997547765604416353228485545524959945116455643894430927138026128539853347;
G[150]<=2560'd115546722739980474480427398013142828912679700492409715812931261214948687077476643410764615230881982208593579657478746189027867219490500397220981367124154655011105765173675197860632932595275939703306852949408934772258347804142784675424528495396861015625418462501559871215969389752361720199645796945084263969184692082567330985343380920153382471235904209730191341545355672631258588375167942385528937866358323842615882222426878489203382988312368936524725006711934646866232444380187442498176807141950215055327608829563488314564328834332596950792853650551175499408734029805898650172956784794318634859592676893263040084603138113283102277627351431176584255104655705176076682816785399684783815585760170384354682521744726073193993643652165869551423253819797807134295414275965133346;
G[151]<=2560'd115546722739980474480427397925638548308531439652549040366519478438834654444868392246416125294134944568058844212684724674525317405057630843853801692572657109569163962786637903340877505940433495603772752233046499028124746237022261328771305857933499832301001238386157593578917598001795739769838315884829403466346818846425781504141914206877417906853881083817949483590952866004639116819241422616032322576302203264190127196374889118006248413310871791582932685077064651798464149525172016815730934698663578493576336430119429469731413567799433803450780773902760145439566669468145179987284415014164798252440904001188634582414093542886428763769984928784503072535871193430703404078558466630145146978900113389338925347033391825897796556240458398237430907868017722398331885312612119074;
G[152]<=2560'd115539697882470037139474402743857410363892584359472314316925722115474212464212956018675945793864505184351152348820092921116865287662510504869064898697120625595469656923628676008856603383082780377639670828081901515972189579566054128536088358363732501728933553953215039843749033008262015764805676174939070891321687478961597517097828402155446146088311242145095299689564326776687624644506047406997520117992636652354334902977413952629059979213002726618982912026570124105164809431916959867590408794843917778161495702955918809664183115074078097835686477871863722972918601415269362884031189673331065147540018674678903092098672346306772893202798895846612751362590150196394259281176787621678711320926572102828496394178138392589933612947304314012218109097421056334970022856835080755;
G[153]<=2560'd88465459496493269409467143777781201790675810000144956849697205763661158676198350590498215134406858912178694433706536602277619284045209577850705170245573010748411411819408981189670590744238284451838403179418350355793914558559133070215999067848110197504582427484396748830210894048467927317147832412439146969024218925514340501143454363608163866742778123323894566649134312662156282375281662767631091228489661784914567510218391531497885474741912760117939676866516453045498422053895062256841539183754861433566447476599375017183023646059021009606517872223311701148622887858905780525441189315543030972003824236147796504075461044923713711607955600950384493215044258550372112404355435994301884377379794659389459086770974546165942728392398779883964812996339560881420574310098215458;
G[154]<=2560'd88465457882742914260173878620787944279274701902757956531911908073015477766881407593834260047377701477821415921048801958768908135575123796054242911198818241250330346178840822909446718181221875621464785538165299937549956601258266958763210729809379616243938118868697267008735755336865881808074073721347337606442723863572091811883084903969642469118352895644550741226358756580381908778422454127406091572891722436209524731834072768694301205017085338589646792536429370659114956096785313702537505295201808617069413300407167471432804864589996627703331344973342438671140856135585829548690448301507954606609355634531610389118638558201339197031109087665736616493450507344588416942983524094301251021429765874479596665546731966310642984512358761039120698882321765735814291691475771938;
G[155]<=2560'd115539697869883971922470567459517591622676940120312734509133384505303627294176414755425821157340427063879939193515370356166551383295220986624702991731492700197619425122582726063177158314817716302464870412103125648503486767647575119229660193295016000641380688172116868280218437990264069542586246787609045845021668688017893638813378065873996236010101078034776825009755620475925388050917646227716402796240547937646793043049918940163229884474564808333471484558323565697921014150669020618091497688638781037773655972964540009608080690841032329929254327289329937789599979896944438366323955250194753532803051705543321007021028497211562372113990769591494449838052431028313653010529902736563180494322300492170493957332579094521856703477215074810220636914634853327814093001294230323;
G[156]<=2560'd115539672042784773137874761808964209036897237077708390621441006648531858062773345472071859475079106971214627266123801224326743296295339291291993094586476767844785918665213984925945966520354105332350977146993336794645844783755569770688320396051070659586013743544663356992339406605149787585463246065115038318126670173755430830175338373939359511286686641696280837984733319755298612529969974724608347439833555413493721898684441496056195405974396430279594730568032412020654950334064337990013877528281127212258871283428415720867764577075655341858255751676906564740745308974909852159415926802775548040493909609747247368859910966262199912537380495969503598637974848607044403389649047650442953573698098846350383948866898587761089036944021085820662792145917966310214245322162647859;
G[157]<=2560'd115539697768998404670953114254977546069019197573880392485487884831846386064133347215039807707789198675842711996192754104001108794157534162564245418387072206921733292221617240926421756753730069659295266630148174755317343961684345522030513389897437259754880838334595638910510174629379022025263015950124804793360346302156659072440245356288247567105629656729184310780924002951762903981330638116181396542365640309249632700054634255685573345302992556099541101647503254399741605553600221031436521725396113195454135840641158937098821748599953141798638674108938596578615562578105679587300972653025799816708110994397221461540823517516487535429498268722424141120135166999705394678146008533848662274050723469364302973916057176603508244094815693453916315058282048083443282906849686322;
G[158]<=2560'd88458433018927122954226456252437156804967733885708061617607989569679458651499469861605752207716654612074528032077696707197882444283678031036094603340129412790421900238963360569081849792821571325863426234297496563973563981427236315199592275250058431506457877812537897719733478456005415315413820541948004080522106663275875725637469271777814573321589956321024457520553402812649631793768361487592483608608135745737354824244251972512148882928057293039038625744021407929847031298646352185568240751981990349338825421615511632072875175539927149867226388152509025881940827335099449134912210494900465426987765745353599159779230295354886684922299496224413896145561168688946439396277738267282440775311309592962433274126020015907839751022903194907174510095203814047568884963980030498;
G[159]<=2560'd115539697869463718019927466226268559405427677260419490029380233834677904170548738085168391858513504400504040853268418373669706543551198986492072276045440197063363383653965425764653000479605622325102823743053156778149036854596443648423796466399786027285746165372874146028458999646590726453877475409909306692482632572888239882555005580266277695159404230026754958553655129446851483944925713149136610148681846446272466703465022614340516499602694219430850324481009568740581583192384238353461372459863669139694241022384289829524100767072262536204755100170581636038304964836461768339684018443564538361502809054970613872717921889953361047214993166759133389792620106584986163712380068075029980923349768929538887764924644950566447878363960383276736891880515381558844058702030517043;
G[160]<=2560'd115546283679267829273206224454734348026439054486359117310285370833797594765700121225993030452593724296146801407664025558103210205963343817232383049428970087595597361889163279902268996067026852040018527893173232656797795331983377699383498924641282970354858092792257747960633416068773964851356713405629376627719760964865199035726622980597758480065452714818391666417643552171803946526500062553281830910666939024893929062977819133648141728574321882353646761652449391114235023829209218703212873108006931415201111086978163916317480178986740358452695354058681469066300286714289245665467041960871708640255145007595877829730461304337329087330671046212691518098521314612008291045665616110729189445259046271563712032974150199510286017325474018211055298682773416693842692681917211187;
G[161]<=2560'd88465432049312101679788652114917014341211474172827402852381276595888026718132566037135344582987074675928783412487339144758347654888120538258203969008373183970397042496673783562652515245597219644803400738725280769884338573630169574274259990755377423263401075534618645338664002558506442109226393568687206799260137193788587305110784980714011253486696788663257683349188550115547245078869953800105893193211240152022903871094643259295788783348251742356197236070759982756623698452348775320567771957345047112426445992548447422547393259246626593332919864300363640645372054581505677631631076737931712404525068077387559876887460960686646855081380339784509805873520852787898065937231317062104188211983626242243470707335019051304454514563087255581804848432080125080413283517159645731;
G[162]<=2560'd86772853103319753193665341698920771143646097995210854081609920496850576303964698753463797321347130400089286477798859057879915915162974693866399961612166210431982382448492300423442847953219572936991714719948408326360539523856216184799749291885592308792804113988815759235105897077112628718189120581785739439148718328341847513209400000605199651920327162031439244989446303681184104089055260087782871875382381498069359541734411066662459329884362274504732792322818931281350288673865444377269110275435338500991800257980741021549457594839540096141100953343704338138038397113689869220557470490195102139378969606685740363606953233279342784624714670640256648738598700208738834001310556400350896357780790614213034595864117741991451102661434780084168112548868250170485147647578677794;
G[163]<=2560'd113747916941287236877044712028095155134553165255421917791512490193721903066041546275285772485943073460696619647771077557934195970507491770429715897732674644762524387898043628507376892768358503450971389421505017670000233708131615821690373672595191057460405698517947139948397608930713741693315778035692397922109529300971681705946765585909495568913141132581061811111669696369275711053376674408849566453433878008173626230264461486500483257046350993143529690519619416203529493559529712323745060721006723432103647922188737891162688795966830080741293515895212042421395746759008513654433866004587520284994917093999861780997073167706166446695674809762473924317839292261620094378548308708634963211280785344878593429696538564691797973447401880796824393045721253792965124183197688354;
G[164]<=2560'd113741305298474202549390532644703535508520675597197388581992123755693495439564091757325968027575911698946383024094649605455130669485614141882945250210553314870279233633153747823780717001515428513380065333603171527612596859726313335130972442958390891452349946069407632087295670558744987043495979832276053479318158718223192776421865407762691696184740832704136460583781312796190390487446963598438353785010717848686356141922782284802871131539976675178786517770357566880832115162142264593120210003246373757780104893328321864752431322814651935815247759398740924919165238255884172974392161519235268869238882662290866541386105322476024646798814523173208804315723710379404446231225315472063284324414798755085852833538051559555970842152277361516594611081950398013999613642994299426;
G[165]<=2560'd113748330061379790699678668912592370520551954942963963620568066779549324889995961998248955937423387200042396312630755284089459113811570441060832596364577960326885132197130017628217530475162913104889277541002532228328121632323488618047213115236083788471931104161785070213054106178472743104801586043680117539382362958103165177729701831242341757435272749522899168807886354055416579528832792688588671739041372970974240535005917589287680949583479710052763905042877880414908386503771898177335281550842042724163706349429453501771166585337744160017168526827641335244563574022064446707146786534709470958585937745393043683769044026006865859213319567332977364912694174684039683703826458660319972687801630550224581232857053654606888681549535208674112432131169622981774049768588325410;
G[166]<=2560'd86667092745900442164330280849212761457465197622871059630889194229704232285412190961604724441971690923994687949458768164078916018886077163712851268702903371622646789253796428714126738898117669970712936242414798511338233374598068315063022859289347180865940676955929806736923737856284810350768529399193076583757061590757728898528927385893216253608698094122890742699748587805528038018264876503884874724493594533045902166618623670926180216743112922270279415908098895041647030424172665846880073535708391873493432104952231372103290105168489920419058997781007910624370086650801251818808705068493969156322522581379642684666641457775382154850822624160647886984073252054347790364932351024137498706080687646853349394110658392932304085211621520340734105787624278855708183175077442338;
G[167]<=2560'd113748355988944199832880788635764573141166607235125770080410534780230645040835505330814449972561918941582820266066878229412090900881147825006819366956368761870053939028807600363596639464353225844757550611788795322843301080722584576619475659769649687771556529064121448355108421994755486094223338250711500855730092419235661857784664603017594200373317135301793200926557097322976337695539058060256965818035123346521510059816006398427927133691356999853974118328642521563655898020487401423128705784857919716115339114709060507994257954189400322690001234143798748145219346167082065750193588021744418132386677254567873276907852159715376979894396481266391657462757938076501248395954519952018992879992790112913102298594678414488014714792104055625319595477778158185190324494305211186;
G[168]<=2560'd88458408906882464469919517012277125873628432622376187574896468955683033195471860297036492009812829570618546726448327320228057763830192741746015142293620198615496523232830917612800937229130642373642157633146562893280618143802598775675673261854348809180887662247708053324898793273919658344913119604954194111640443321312894094452738432236813205010389179614298399796415634554786170174702926617030051048893430059717936936756044748773618151245736931016051124960357571533046960575153645361955213131838286220408762136828279121891980614374328170730915052895351475950806533644377530134342724323124443048994088657738308765824479812372340975550430354462598314173594254773469329910906752684662143043960295407056631002531107296627864480079335427769605953164309855279624467057896272418;
G[169]<=2560'd88465457876017210180558739298088390231195385908864625869265837285188960442730854717686879496023312052215202777526170588552031977144647656065273295976445286819052572413049974723831636134182625945664319370632625531182853790786823272936194890062525271741060393799737025417054513546256233577350276603443814331112038483906093984118947246305543381449311453037901861856098847948560146107693226311911963006680803910701978752556002618560450597435594312431258762843717607939153687776414589444238729810255298865701772650432833000734426813196907396135113390662383220743683212876538376706271545420281791518803002303791682367293247729404250794600150345539408642268815991215057614422847751405106218930605399963152857161881355573237934348899116158230412050752724911676138102494239863603;
G[170]<=2560'd88359671691894227793319936367956630219424522166507737352194292646464006921697194167561539910344179867867370658219073850587389302724263575503997067125210522646966996189472083877146969912374797957975606862822731290482855422109355003339381061219331073972614197163469028950744046897654948515442103629801326695773984946399833149966051980437394026558375310117759861673613846405299976623308887208310031405470245211980611894509377837838309305597076092904172703809595931638102973117681852250469694215851597518623051395065387474005739885366598507464749310670262080692562500694934899139217398859947235910857420556860570813971396370516765971044578715172437022423612553760070499650809654408358098648353925527790428086895104370139051382103962853173125234271756029255529681255703650867;
G[171]<=2560'd113741718431175714024118447237919878448438926654456852798750482116454039604494956403869678844454602291509214156950041730387188853092110253544493856996440869991953613933971262432670862130162610267696590963394408729072610742216307834571769395183441869664673819550161727467831050402302423164140458998282127764366391496699270505898953418072636753765712908324393783260521181389626157539321193720250349757999846000265554856618696068187277881772903924859955351896864639431743555266289535607435701756243016392842100668203995230359642914654161814633204706260106494455308250062206356639958327795132596712315357110360342639167230315771393800581154160719217547312060043895607439012934697668468983407577032718575551023883399563761666053732652665287924972585230516369031608530017395234;
G[172]<=2560'd113741718531667196630705111224937734169333510256369231716623844622243274539376466100086609835864524286225438783119839123498442097596378014295408438960405443477241030538221731699727232371904400235493296131833446482225746528365909444719147279778057911738785247273207923693069449513720856090888296691735617051727854575254416158316575618170017652103780462856155754405360342652320163072122224680135636699041435440028316707046764117748726257181371038320734527661264308591892171286097131570361826574428637815920465920162815081932694704131891988430930842744562672903125011282686589807529211708686767383907563291040888067363895507374886165269582012253539852956722488871003455398061446850914517731261129980908675456970404035541544890195186373393935741279433090363240029938892616482;
G[173]<=2560'd86660481209857870253996095267493893809253665099487406148372942674193345378274131737568658881282684997841936494483420797161729900682270769819997937463165035682258619730506105324464585358802935598649240482443501448948575706008554897488150503439178628617623340372880420141241894076846450180979548449615392639795598738566074140463829573548162394452227940317963649126098685337222890620914285162773977079732629696966815921761225301516524820572443862069708470184450493632193302786010442122908978726497873338136005803573882872535467024464070992001598421619535758986894906735811567233114508301828478395339157828731164607552772492464938197332934580835761955788048989553450978264218545665712953740053983859674798105925189884166598918413950991496345762472038043153541234364924506931;
G[174]<=2560'd88465457983208130975830019325293843907760885196073998519347835790111974868927871214788320175929075743223376392095244945858858245365206860640069725382287311158839855558533735732400434507302440955275153402358439236029495370770695715885004502119826227345085631016711623370338334159733960414857231941680020847100695704388082052053122388600313195783960155846796446748342656960297749531707891780748595254758414790931057074163332984541713307779066090349255793866407385986583911431110002943188331333972761299264731644797779238707502821363864058097965670420947000410207821515250834219868712916235147887339030101962329402390860894062251477167478561089879467908368312089962085661534873544067178847667126969428682036362410368848483651535219389945903492917995578202449640760498402099;
G[175]<=2560'd88458433119418611951351097976452979021159067532142428305848460098302049925250171772866193195159698843035603345553378223080467119797086677617741976507946191378772464929980870905126371891476932428962437977182210104798996674291142985361395315932343746254162095335836012670494931254965561577446252703122208562871977208388427240184805216967151511552394320809102053046393106549318717239883844147101509886604884357652300856366090017480146183437586238258974771878737709738724531674085998339491150777459926438393750878632237369240259280069404212828825828500637579118863196222184552008621594532859425285997097900093675927761874467632758474196378120842397587650404961302965422057259113757278326315838923653659850548471239386492788719375961680534770992213772452165304095885237629747;
G[176]<=2560'd86765855787593793732341937595432799895471165791851582760673985455518053998346506734352370048600054707413123603367969821685458557509741694481517599240136451985684252910788339976059482952343591057860970365095175271569101997052865081465667553432739611906001577146734140000661494832324869128715029942879446374870510265464573148820015466734473675122066915816030215000092070435864966498875652595383585000799220011964641944427681300049828082397510872609544029343690945031241807584218512467886577585841535091869491925457791656659524441332760905014858735394028400491838328010346215991238089805591212969382060559633930097107388193949186039356367712674535206312604978863056287423074935831067957573968413113188767711694898808762711185968575607174456307534351568401778612345739883043;
G[177]<=2560'd115539697876163150195363348572102292445163693093528473837794199984876596896203438895259779062167117546436769739480899986052176435955322691293544009974107743411364920178330248122727086135447495451101514475578049492318875148861138513888509132910837138363285027513196180154953388188880966136050441313564815192432321953364039373473152612046897284454258305520028558686589177954967362847391796411861826729247294083043204159563688533238236395052272563982193794357930010472755166386444141530569682210808925710639952726823892511505773944580928123675045058462954992935312501967232000850041931622330159842236451375990378870148567895989492549092369222929444001064091210686442170706796864653502262086413596031619193692833862368696357900272560102484773811194533667552182423085661762355;
G[178]<=2560'd115539697876189319852292911707030498766353879114962661027504560591298123073018209909085345367518415736585000112592540752818348124075895159690349849612093991036287698783781754126311405513867524986337060711184701149105178509757730878466377220520029288275811926329805882081503186391988118800468193567514089813193850786272798489440895496191777539611847450749635306530436637423349707095472308918474352851937099686453429178002386584395588642226376286454615916709556875134223360073450217767600608681789570686949609064438590744903405276338908855661987914516137219256161494725140432411198426724421650982638937129413159838613731515490515170917182537399787842729685963857918723106071905287437344660467514046565524093620524028010135899870570272205135215542708629407412361329972032307;
G[179]<=2560'd115546722739980474480329526131692994171050579650228068003792669953512859360647854133443976516690688130449049772577394838368026047297002651020550523057800187393930491412602776748657941817857983804892100159188344744045978246469984719141374956385660386606574871078526010561538361395085631710410782256718435215414937164118810778850019367723207026726550543640084678360800567617815314899835064681853501816692553682863595739875583700655643859811255763384261892896560075864915397285192031917554354988619272538973997512064548247797180876237108714588656763452420943987426940567404714882233977524899766509586397827446407919308668663765788622302267533639285925808988886909494424932590802371297834826782551066277879148802796646250023762094250363481992674920867917983074652297532482354;
G[180]<=2560'd88465459597797550774002293444839149696732267880398671379200405461091050511869719583291883958031562922549145292503827862461323345206183830083815318396943102397702722640022010953254491366123021078797060194108539484307143163208235353737582529195267971589855778321776452679168572104579944598917672687453018641021442514176469218302168366747419144274056282333920846391359171726823330709148686751044884875192477418204378514129645495853571715985505352375835074584795361990411665334593406209108133830166081460585111451373616330134789414571715869738377131074551948655914113940648994458669896870322766789700875758965029056980125921482169190665100085235588480059775600904026458900921071861498016822022809738303631632262561819213933556765253293404493506698121099330269350327443731251;
G[181]<=2560'd88465459496911983920334036944746879146611670995229149159429173901286300536847225658974396393109649579354769510057292508520030542768807361216477345977366117370483408115341720226433018165226065769348279496058782867405180250475172939692560074894626897094105440616467095725308060253347937064529105776339549297382714155953829828344874569951955346970489177058582192816132546987770776166346213449032478418768724338583277223116602397226147210514608375662940774543576724146177934525141754335238054068901107386090671980106599955738098401837835709611470241469822940233118922141666167620403208360466267412127637629839387339334542212043203284510449689344183043337698104699828695002028285012303590502738537447336427357132610264373500413241924749152427738269965311945704991366629765939;
G[182]<=2560'd88465459597797550774002293444839149696732267880398671379200405461107122508902340104564912451291749485311799240600923575268931774954478599897199888741823811871830568391140822359710144227806943045336776975414239278638245785139502132017680502523599644118046343488715740157686356337020066763924313144456195238732174541698023353147208210300747500325810666376246135323881583591958851738001063095470800768424171316970699362619825063347115528112846761787337314617938526043666361066694163971797962936807986146875747500440186363429576413224289180212991005658769404761603790397673243359909293983826248833946082303161567955160263768448232087771497794790387355343839064787505494268473402721229024665502361127838918096879267272270382854710664228390124786315686044327212785799777169954;
G[183]<=2560'd86766269014901796062988102815302622931738129319293792376741570527223260854957432704307774942480961776248773698756105412408930811630633088113496035940405718162449796195660525960889161098834479158784892310556495722483684860226598778089843227530742633707031600490753028831544886419477253286309077946109184686551400529785089924165759759908697062750276205614589035508918752575834406010219124366409801785792827876402941633315130426116265071557691683648648109672298338601424648321407637773979665509807803426552532307386159752455732021317350079608101515000090956183532963083654678350760744700368914607698025325886916722271118398173354931462209870784245438532692225037664255641934585229309925181540710176879871425622959543693991655067043006878755321663981165637410566661851001651;
G[184]<=2560'd86772880651411118042356841401889421067330502551072460638105906568899001148166278729042257118068485318320449105993017040506955884327223349481780464346649753599749068531889088174423954538040950838867635524942663342595297650766485566229293909044842178200992648650096723927527445807262767606063344459522704332529052643813990025257640292870347066467071138129434824754534942580181786377870319176557351932436050788346823460299262852928595685581878225133816999684768890258005541285730653390559336380548228134688803074049146933067808492525239666093486561908129424555992734198722191106546764305746728729754849798901198938925026331440132938048007018583883564220540049339091386325834982781676951363001044618315796941102056181792106607031809539565497847468658237178581850240266220339;
G[185]<=2560'd115546722739980474480329526132034807767160513149934207133187637855753614292305601502666089666414132916136866416189279274022929393148464687509833318100827192192365813389044246900089360043787883963580114538231644845762338971875789638396636867339156887053078916593575895935802960009113003627298763576214826817597727872145686181607568771114341289575975780884669640822817581753059350783394193305136261399195294960225490742276204801568286114052826555482710673751236233938231484170472963608098822150825247812273548528761143683170410674011732666452243824768634601124714055404888061800860825234472423533855066723074454354808728333517589450549075577633787636706246444665461316782150403040655576190256419666024063074353475569078830607032658508820572245188258834686435021962326782771;
G[186]<=2560'd115546722840866041333997782632127078317276135992351360474396274200383729588400457315570602681704540971193679761565243027243273784211233103331039031891978519302543700083237420485492057635519154044632836153920236473442224093250425424094100376689456854364513219429052182104720216811886017317699531879666435167452559253650385596939909179194370280312117150810214852604662033316581975115812200441863740579723478149223641882708552666527887518888254538193194887938367708850103328159234411372508001845909707316637207610282782612746211340970472366455915002805249690989283364699645513176546602251336873180249789876231645886858867705636187095476622015233314878503607994470412550856732292934063376227046354079399991062457262877620476163141253364093792432384198804486666902737876366131;
G[187]<=2560'd115546722840866041333997782632127078317276135992351360474396274200383729588400457315570599278326571734755465870332131438942111932682976999580848846725591933742976567668843760121806945725791677139426208527215977492027762114716137966885302961804897975190370280601953833566334971409625187346301402358647392808407328396786754363979403043192162916029990357179804188551025286321611187625779893060708640375374046891873118132823479395135733729873417834243035102770587619050954723383647237963276446799209816723281926007984185524782056963201882477647804184301532924033801274078896432525003617886347558199372162215875322814711917943034624400313848348888960246944659059242490196886988381270510515377193607270098041541741916127985189321039906316704864613261477306416649809406270321459;
G[188]<=2560'd142627985882189567843586321954178700299176010856881572124877031960185325511096849405328942890238859072233089536682144250107340336573228308023644419802292336032324922187910040122774765517593495830634826710567521215126068092581455617748364897011072331464523437034947847191134018859203079869610957298989601277399822976045915816532582923374232888565646532837011063447985590587132457702792969334458889791980303486237149143952599720280029958726792860302806193399314961529883822824153388011255740850046568352503892107915430563572548592822156491454374990856821407353116567844935812609666553959815865856121471110548434652235377998882485515416705498428152921843779602329592592080264407347526460974464535217517782707211767797009054971417630554294248553014802228226687197528292799283;
G[189]<=2560'd115553775044671982963061113299530222941617574771310099128747948182707420331616372522817451912088240514547353524591591980517050536660083790938723388227941513387572525268920202607112963039647318406873898300994415080987240245338926413792941142159159547136954839060701714014090574346722732661481120738463730140570658305523945838064186622966017488059967828363939191366554654509702990494404456782381560699531616682253123738478770918704244921948397725655373997581726675046255390585951636675462691341570231211784907366477995295937373141018851935990011119307347173990805159956797443188634847637248509169779168432779018207146140744466531661264910462614037832573596298762940185240248244107593642166824714046143642600873530271064178417163545321226759553914979946649014168379454599987;
G[190]<=2560'd142635038287740473524525061522409471612043050702934850963051922554183032967348669678980549907746197070834691837840203511111896624466247531147307144841913840709772688190797406417301255240300976425453297816460532960947061456840574338686819636060723996524694500782389769499107053427729478517086752614232106047033686357156041740812871538069217817188619877735515237234374988382065427207396202730808830611450270113456341200914426690636658039556680113580497837584748870147493409240230962909678388729928683811036960529262999491030209252499991295811122805483499522437241817621824020647010596757843175493118065577356710547367617691088924591930208668022890834705449967486584810512416789947276064255528170303113344322531893139752844349778461167330626477643533557788365282941527601971;
G[191]<=2560'd144432962649234474625377460308921317708496549953101969166517134816247468544710315962633728031541483550503299381942149786083053474237331274265274934588404887233631041964169225706900189513968845768018697084879535565971396367979193599865676351936006867102027986460195727867757415257169250592153110631924457310454833032579482842385534984607890840807059425613024522740228463719014349742289908780874560776102023450533570212346305641445900212590856974654291217386843562682559056544611817244887516355125806475547523865889838591774728337228799982249645978375176104775761203319010472918105780304864703047139055522012987415851484378535411147375698506600064700798818275040602866212130384412199357265907396668037193110351998651377131488680506449002967753500604088663403079721165206323;
G[192]<=2560'd144432962649208407568030223599843305219609471852869789701258734507446022350914349852882883535220260407670185941399337446998209564179171703339301043391637316152766258160131263835161589001990966049868608165449363226146012703459801059019547162287486053262443509582598132340273257219277309958929561643392823949212683114823834385356984711402262772454374654276857762214449917550708131153032418802067326218604124721720623806024620565636198393538863398335486961034481290044192503522521912833321748300068203860119982990245238285049520541090716120356031172397459129245506411887030745355854443632558276940091024049328188342955298949938661588593871319123487535886082388643798636316231017141295466653593619819038405861542255333082341250611808808771634079263337319235740292482075931171;
G[193]<=2560'd144432962649628661495444634313124354774782849269215509234031332805946638802264592922408005005779631020208022236421400265342719690216768677606150904421430323238249091635025809658182517728575351811081618215943806290817656487483551049264077442896103077859408577514261709112791162063896578512433189040831708984401622496935128899829720516483168470275902949581448980389472289011092018231066849019525325686820639833333864395335404898638738822354798288969394839227711510570104521542473390800853387145584274428890566848238630984293013917851093854194812507476478281518148638420905632514503424871527638465807291481026503844615503124647965711870688562732045100936836727739061533661717350061394794819004881987712606890325205492980336356831983815523111038084593771440350735157389636131;
G[194]<=2560'd144432964364683298007804972413597119466146602139035604920591219613605372430694373675366810812520829812094869611288494624258787002515987624034747515079490117126223178115717853076380159704041923617339601408995232170979954932718866719363385949968403195072418785993697407422894367841991537900318575327449710384480807815388119192854688836845847881218907065538936161696520679201220520670958176736471152430568764549621216502482624435644060633617882015075396152633561705873341794910418825730094211515478999728034543581016341937730249054303934028089828572776306576077839112841327189065436227473881483973740347552493753982483820545923271967837805283699641745869762074916493178354929868571510077383847871630849800610978882198747714410542830608247336876283411340580686299109193364003;
G[195]<=2560'd144432964263403550696640592258539055204017168665215443926926485816475408688593199978852126381060545426929314564416123044423414454338071945975017491865882830351561214664073581250526366776940096625277291499624955474638974063320982625621184121886531264690376252208208022415059008082816486294676078055252237120874608693826327910410407333846502559074142509481271000162218820238855987850256284761082429836588894960668893169543078561484527435373231524125587822514351473765549561391885283193386908317763865908783501501721478629785782883665302280716241418917739702217731447642568765945378075547030100845260885462319398084935466643954157811919910891964068930803205342770336041033811836983816510998737055807832305189918106453710369955427130318578876924772763213729380372988829053491;
G[196]<=2560'd144432964270103079082491362763389805055644408395864439312047140339444566582139733912534493870877803184672234623227304565834891849749299202750321584271975915183389955904387943000623900828148145868343884224306151577078601127801816762092622921351102245196902846246575572997167561208691995996840792545430146231269208710570992063664233807383141815625354574720169335527040885861677358559573285911225947348032191556690570965020364334417350291351609847137800738382681564137104827163262260305157157727930790426855381120031825942827882670738864615985431534157678418005090106316682646886933525342784940622654677601144742192172105611283973747210083072617675905353458487696205698648702793702940013199712157030618006456950136769296519246193704990718296112421977449537083762258824344099;
G[197]<=2560'd144432964270103079082491362763389805403355179173207637160674238787085223731020878878914324099920060225306700766273212009999202801138194772231276595914226826454697539967571848898171785791729942634454730126819312894889910050223848219927231833633029929796146836673442369972845699247547793938129583284928810985257612131408808532689470530915814694555154149087024823284312901262819424481815587178721950692880380889008114868263946502924672269911761499371752314999878548656695990733673530953935419670469979746208962974155139405043738389965077859338993716821579590870953098950896953532323638623413657185864426958803241366279882650944339552240355271497982665278716361063611648697505804451032515217917431414844015247900897066711753898620338441019894387659283473514299689141997351459;
G[198]<=2560'd144433403424975593101977833868269629983028359553247146887144108186321917675183230277447311366100512616356737011469953456808170085214896096673224337833621271698869899461174035280606759573145294129517215324550726087187904439034554152333697585092906040142063108991926719911850611357873388569374990354546526542079288173840938754439515902995059771792705948543666084190184872656626545011806198061888587254826465741910931505167564508386511506070025829797230167519837443954952937409744422225889406885142626786032137251008950019854329302818034069714717912379651575851821453049247598043514797616165480602847774972998258539490219608207043635160521967974895607192166148236655013701839962512091399957387246260248667464376521153119966185071335160027163657744447539157670371411348370210;
G[199]<=2560'd144433405039144662784159189335671034015088476217713133368761947408388184150454168636927079218965007176632751981845655124040491923101669138001717370436385217690451492757447195739329773993332788690179924038630565915242332152801923252945576586431523506787989565973309530549652725484473126293661336561000997484691414681111935363022319920407469648592806008743631369506828629891757598557181612558269974248456926545204742129409111925371991424618788848238772117767835490583640185165542465542166532452285091145736531181117845436721785754811500477862017232468435687476198849737030789468859528288460448955538031117813267425504374863599782365624393602530777447456900142149867669280374094393255204562390693209382706127194338089294789871723218271907739313170678569210367422453570024226;
G[200]<=2560'd144433430973434776750100551007864271741391955345058377099736429711189101240308987318441284501530128138165317594515671746563749717970900693523008309304400179680015742873477607408711491993190754462412096865985828718870788776272447135911444710423332677089887166803263135887102922468522548475487107355628581454260558779081127613907528281944833492797014074502705464805106542561100021958368689239559037248822583145522171652596229316982241610440574259192224756509782656895193878552524795590013954522637163474836668439743317847882649848509501949751044205525592819646686136175188302781966864383361597334589369760940056447360885990553800111079445869933028043511700971437148098388867873582411782564583275409077698057996954764697239227499816963010443061694265232103979806977594438450;
G[201]<=2560'd144546242021401355282619094036979267890098643054302107817891399230049457496491041898318257821533346632320834780737946864112276557630202387332857999030122865375691399154107839070888189981043962166461608095674462648584318680409168984822544028317184389441640887131280966536095983671627947548127459796452329497600796208939399768161575360953725035521923089322641138169690827669906244849678707952423901474055650201392535789451043221178118388759924997247637646703612103696141635854796139069981749922799320406085940835612643430280170209625156280285761362155528532946623475974314445877371301830150896890718503914588284307165691598074789837541542083218512106561627811233594341894184625783249618202659019361890420708087729668563168525807332144465849894383573273279679993101063234355;
G[202]<=2560'd173320084109996983626232996962593971088694688969614854039871639958353695541733800769877442266251813059108430002327149761423542021619093080507489059446200598382524872487870151356861700093126007770801449586875942784372063532972161756302155723528293388695811468885259456010950119757662088863641581716626351572297747679187985876163139254716705516889880145181144445439455825578864155623047945827329283607676129034676919638103947903937638566998932083894811106361238773281851452146885025165826683889199045297164716165332196839053084696338644606805367809835933496532400384018734326872055871573770761999959264933629465000815987592614383706121911621726511640566810854426692128816860157351766999222721911301225549541488868322447933467741488519695969037005743673452937193257329435187;
G[203]<=2560'd173320084116696416177405506298035575469406405440692603559434358843489523483537070494037421639040216194996198592573410104803849074728940439600282713142339987430416543963278355227907520687927193672460845473719919299652357235476533938008039191999156690397890237443864501698746001477058381962973337665958038684321096725606894848307104265768606829600213519428623602053020619019167965330692745094755981662127218632946139769214403785525629416646117670967498872949057148939091939180032867605909197304325306541339844108660989478792124034345537068998241140130598299240296626455983512415754919511796168591423629082164991603778681467970058263933383208896136088356126025077674422591880751283670511783956835701575649151337807437343126083943378728734884804259588757401554809346168402738;
G[204]<=2560'd173320084116696416177405506298058274028523080712472320860405957010862960683248801888344445420172641491905769557375188681495344590999793104431559299363203503781273112398197467212675279585881804109008690072721416683926997974502348654708352291267104169782409116258865233125331097245367444658601431127002386479471036460049193973381494246676656050022414031913637635023298926978834102083210334930420152146389606278828930083333421293981153150723576319345655845942013122423536574448162304699550631840008045161928680002330297424541638628802846203913293045012190326331419347674289594581486906047025424146767691245406139243332589052656042016853282169490360900423127388911204460721478342119796337269428898992103884262374053244124551829538186708035934654203254533186708700690182779698;
G[205]<=2560'd202093926205265772615378191028203749720578488513256486658669992676615569982820616559272328723622733438024479690556296062743752020717895372786729876262201011305066618120568358563286159433915019459743910103955404506786235653940123726632058413152237627787797370502796598530485931417084593585234581831050215008667772076645558429209095118083122547518298349132190352405620065602619578025808119327153422530088086139287685978610748971267838288290563243170609396987437234316278318035736012598334822555499490835941578306447045973906233799763128485518325269608988177982419879507102197111578460374911398198706073944614335742957964248579630211018280901086032974879900751527498727688787852116200521865066897353836535919622257949022331489606728355077018998767415231170225696122913104691;
G[206]<=2560'd202206764794965836355293124224501824937577540447413110445698446391508729173465436243961296818536339289243276370351515517530341573929903410909136417662503692925687750980209920751943847379026077858930456183073123049972839782672344589377244560682045138011129586004150545100391803666408637414170212593215893090808820431295763261071249344001587130149642170709157462733212520645580365194735888368058250005585039032393685226246747322098111369245858102927292592951648472082899266932571277198101239515706997322342212238055534794558120321049438788748796322118797882552631113807407874620311788498226663324141743242451731244662741175914735917484464494170692496800078355680367975038411206186554799728486118626745617213489627057417142129290927768621303121641264288067408995952243188274;
G[207]<=2560'd202206764794965830741454159581067268657153938321535133832722831691539636963707802406167276498144084768787214470417530950934313155258707618137462266974304619749649788627885365528909955846028075070100603964667821850935003899994356471397865522298993168343988765210219948025926312269701320698674139113549741987010425473976886659548937773002491509541168255974097387548620981422498326472423072010523854482810381591728565024605058961730044707957888364281695482880061766162331437290720371786880570471866393412360149543401782216408345837835777977721587257513457317829889600171090945300937602712508816140317368205376161584307968684988568567202927878487333157157976676405371099900783996562827556834535137609140595175559247719320749395552326091418689176474153690150346343123160085299;
G[208]<=2560'd202206764794965836731121528498295483810995286654075820427085133798925475948209467869620386522345807035507224608471681006365953747927821083333911613660621576924717427939097054779208598241036933712999755188557402245893555708639223050420202521738893873715061784157891022493717611621786860275529709980111994290651577347807872833800117111965554722800135672512325427143069889204269697771766246622429977232107215759564471039422545009512653163316991522658207799910711372284699753747393262249844762354676220962021113696264083944983409454961956727092103054955358684792472106809805034564628246580851553013552847539271484232713207419319827113520833757836138678224819784175842450637198825036854121684940006591681842477378982370514482849960322071237459309095525666047797501655545754419;
G[209]<=2560'd202206764794965836731121170086231146779124855504652175898103063331829876715060597335271966355115306760799084866192070957646668382116406207703518055511500184377973743935385459688912614974297876212492975725879517345946991730813693846826951375461112538082111232771235496541101013646263629322318364485237483992559149023877114513296003726759263126766166452561996628741574146784941044735025370963197805453292889182743195531084573103749103915104129183843920292636828813738460365753050106821842266044603308607590808955103213881121339939165767815051840916734981867220958857857525666170366593104581635925229232655417216273450258064750184302981453643780560139415666231647911827334826253977477093417924174304477555266872222613980286915149211341422686362660723807829561130944694530867;
G[210]<=2560'd202206764794965830340577053043096491800135556380731119920578647859914712939127630186808687551264149538066717641746154369418958919648065685995645921187661765078832764982993247537250419530323527764591967215091863949432262650575634323489171619533482371801898601397559152935508026140164881972894652390007569217929892510078093528070426648106030461851235481700317476593633385295720666961256745777887502738879821028855441367982291034245867039213842450984684949100214048122216834862831010992324232786688196650398878976901771652719506122244821755951594583055878292891507034812705192452378031060102741746422615926044877397347169301882901817837763840627285883985217822277874221306987779827657970213386056573077992073293419169916641586215394818175845411536080826534935620850799555379;
G[211]<=2560'd202206764801271178268937053754885931823587658333574027175746566597140267835002477551883076465502708248231130496332291426540685497803200231371136870510288687143285185754788676093033686700356701779547107756368304848031775484066789039057705012109321540896265545223865492458705988547798568529266726143405251872218112916160213144496650530465112424629067884741259974628003745064704677712422003711210598944028214782247000676543669763262954841100418290661388532785193483288940275133884218386754299884668346370166754838428842822835750091972587744076154704944248341535265157195654987337652211666370035471241009178722460024180101761010300620930518620370885811986847880928811878969060671736112417246912167100410539250692834140803553123044457867480578133300431471385888493075631911731;
G[212]<=2560'd202206764801271178292420570540277333961459855948630839145369911508569545274271495622802072242910382729748612563251200602556313749799408538574132097795185561552321582691310605329101393925622571643703864775541578752744978660392990358638454232244503206845378264006488619837030110503949063806840752584377261048555469602849680478502126192530263032209891055497688748108346450152156527907239776880496182954332408139065238566301007337154544868811239275311392600396864723555124987224355108252644597133059203403764701059273201099224304710142981995169892386011647654744604192380418271190962346695484612126075820560466506681548448035605130010217797580580724896394523156871349004436207740744097876378739446183698779726859013193431926518527785798394647771064001912408695950637758886707;
G[213]<=2560'd202206764794965830365534001907012695023734562517921581926628643658586443086082075549327923867822139449773826546341551801340289622045329269771943087845384217641732088880233981848579937998946204121700664805998864423732468232867161412280121065717600640575249258416198919099443314226927978174504865541044159902009126053284003209010075712231026030297598027413648261974282990074771672588243553354625025097367352240223534315439204268632218565219470561952512092970725574660669192476474644021896259119019030381603735946894886635449917528248844856906147999565936682312708294861247870054005792372809574814420556742725085202959541265502370590097872633738905352673081344782450688354964463300113551896235976849793310534877467430660126598494128878947924370046557982701926088323210883891;
G[214]<=2560'd202206764794965830364157677178864076640621615175008045508491129682400206748389683972171994716730596332151534660341228055355785530583346802979167896910215394636252878589728820638342418985028972484349846431207494033942980324363608714426147954756755481391526403844483684898601692274708246660122347650411904869071077894116691436818516209344706924112442104195709434155568817760925530573810491858540750793708202950032824378206479476812652220214152737867797671006593110521033633174465022348373154921177321224884663072823135866738329056831402592379095990127726810661523460946944814269320198775867548041018831490682800862037962529881769730076750187383619855652383362288501598180329702195482280423299283980723499408599439414191089884463946822861116877465450266135384273476799116083;
G[215]<=2560'd202206764794965830340674520211074524302039061178409244843918267594069178829731915380527842419118826869046329103416603794619792773499705284387344813796402390398616556244004549108255294750088926469768640149545095329035949023961999781250607963582309666220094235944964086089853872866574185537664733096575391869945781895187369451357872039077124053389207372579984905672772795682201503391521509709275992657716278284859241307623886775279046932289370331418822258067865047406945288448771212626599131693482247072929201958155129154717088662993503641150899910279378554083823698666130257078862234040325757599191443473304508726305978116274465496367596890137972199759381476091194250822853302558817140085230557945802670472525999842184969967122445210314594305049168042951139505852938138419;
G[216]<=2560'd202206764794965830317093536257706513907397295767942445827164743783456118655166687420624624783904546229927417655769507644668036147464284913708153980886719809455614489240889489076794021831693234521350418934641294066058186744294057218917004178791370486584363225752976100190876297245217634533172899995617198227416281290369372572993663307631950964992267455794827802725312435509182072450964589586162332309188995373765111023795220513628482339455586333200467251469322281445508644077822630950316827379039650716127188766222428869203214234680155116618093015046187012488860908745967049345900265988978012278518067672013062438150192229586102161044586155546826230708682974273457986952282390242802053286006857932545113629662445923430925182527687549723489587062296202672521035526921401139;
G[217]<=2560'd202312990033101929550557182203175902649691532299164984245836705556977977297548108546923042139824876231092072435117313542242914430154799967823713624336211129961829101556502955491349082394121919083945152085857002082535747292498552677513249240037002672602184895819052458295054774708959617626047694329873950019668850765399466638489145930234462892470158949382415774422431987884691895404245923347686160965774608504074327831580399435673635962779499376867828901949766023689234137889112889398064140012463094567066870990342468447488145704259053743387853746472131674043994504054928855316525359455539523376934560168166567021257070571930283018840678211096189307437502003178521784407389352137846303465200019911192010489039721850624477255383385202363319416769206153211869622316641170227;
G[218]<=2560'd204012182337357668749361991948494569039066604514340880168345875656984278955634877261575288649989561799197200820151296229695321801124553619774396007166494240966246889880242024493276090709790910336632473419224892296927321678528059601823777948997887423831286838686005595143553597124990904491558055728808373071776411485167582949813787949860198389880437185466547064940291060351945567193000535977943828728398236652404325757056278089354772413197242231118708978537989748664817118719771415530728541582196620763855052506982148795241977644889481609461531065960043049571043995800318235658393939243517921106109550825369570886019915675485970026064015826503539581861977541323644027835951476146748891352157662383153206183914269957440783609058367668832583698894474169353316235704259453731;
G[219]<=2560'd231093445479936312306243636679167430106287549127325582929068861819036558278314234707966685888424268242247943669655348455543184264906197556893203746389123718775223424177422172782746245515558558739611676916712892132870327377804847310625763211686182652521327835818694066799969875476514688742072139223565073171804847270207368249229141013811954409667807019357476724763366155651116124474090872837723196255588879855816385781254438786905179539542314338229078511170079796599305248825794987991323836005376649115355726970976205114244494794265797116375538431665431923163036960292194476819079954374194394310420038986364764088333801756491998647989426204470806794222049401629926018728254161257653536800713866241031965189436925116794502818745754158498822620403018671454212778384793215795;
G[220]<=2560'd231093445479960948960756924151011255388141323982689443570989006646355925435891960358549974341868608975610202671620564965768235841089168947316334854598995250295464223297954447972598041652726396783068120855007298353100904935302800895774397398040726178346199636474566274569945654146470572562938802632313552515484993305461088910887764541658304363366013285540528697461788248565184226021561339758096493886134750714400799155374711531719095607616782784424984435877522160451673796825145688204637008537203833971196670947503970279327671213528237743802916923018678055223574975680167212448981222365439568018176467020207677779991974046157192029814424617817270890173310630339895386980065334201402447998224269935096792351076979965001223020466028480329498260175665984495460905842612904755;
G[221]<=2560'd231093445587151870156813175184029428501041557337944740732061488398161467380373290109678832064210544324561612810081239744983762204554049967662548296803499871522136858648922517478683135075426326244536839017008234596739099986305994743078828925120034327924190502290461448723130128810783993663604662118816048346963607139745787285242475946364490261843957777748210749438894400140109993226579906469903491032842762071270293428921200813122647201013650644148252140949792117001673188474220501339100324664406193383453180427080927020875418375855901412016594640849506002716246691250715556798401795388962282806938514549158133092753605244458601462534430880554648117303454104616082960887291987285794670723473725394155037031819741147327423939380219563629609939817686290777812780767991046451;
G[222]<=2560'd231093445587570681280531586918825340306593988528419704784768997263065403931639606862211876270525464747524252044375065721036008482906468345668841325659159801197121618288234368495263958699821413299572623582247219875595204177780212433301631178541098828597665943122247699303666860504708047956276651176616193220223455641702895082922511628921869777698691232967424082283165781013756755076619125099880312235332506230544167302105694846827603058465679160254797637540868934988861470545094548880699701942987044557998830601514775826529747910066171673142869440250289565326770826510246912605298623199515410828010255953231205579435369698382983764813506251639622001104633746264389950265198523712076419906717924877042999280121673210192728091658561819748223432796233900245240661888867709219;
G[223]<=2560'd231100470445082663626908380740093018126628676414713026849080181064951255178562785030694672132727385546201337555271768624804602671351754030328097220938559615510617750612282544536217209807523932635211451102216532226754214623710751125121418612889261203174691495921594145797514465900181619389870515632878919719824515154962893565648723671557117807720659188482625536116214343806680216739846371333927725657435819445583719300390330475755229961811976488902146926537040393203751622232722862059389286944309060280220373686256134595358616587287359422053221647784860879494648945526777561110131804081506983324924706667815391631707685515405783459496813116569211669499878391842847715212444416378997678246162264896335776496030968664694304966481290394553634010851499061586191246498944139556;
G[224]<=2560'd232898863022799410144200635368198198811759139355873013441988371542157580166218363001918169690069248898224786444046028151911616899530489626504543470540346114004085696478995828880844917068186386303887671333794186065504048314204882564572593741303655532119086285213402718998481878351875129472002851552066827816459654578870696236571417778265957112927796626873997574628275414141733730603090651618615420341392212632008187335773539787604102831362756618364052782614281146142347566884240576018536448569450334929737400083926687103595023773874572335879457352589225991792237567117270323014507015174344060541349781332314432379326138281437893197613469269482036769011334564504595639227779642802790268391499174313102015072613299546369904036370067208560533777567833839032256479112071361029;
G[225]<=2560'd259980126165376424109298386359235090914110092126904546495232452310328828763000854042727113322735931726442456185064550299068115002952669314275659912264306301772982272192135378324321120595191480046108868247526283095295593464446828329742485868887292778606833507645837857994990448730806628353277473887827599353857188294893623345995697186780862481737166317853747031738038974988701377587297220589328661899761174693554632779197180579805127374382362888356302465740154658021544686066380855884699922071794609363629232078587606646677694615568822522580914241578668628271072715924421379051023615809392378646614619431967819417787074807984820610174005246576074087841929131375369883279543779007822563266996280009949070154819946467159174618260008198320547710046371661920076328493640725268;
G[226]<=2560'd259980126272567338891418779278284760543027027996828807674973010333374187163879525568396516595226676647704190560142489623998578199528026331028235476828641380597114914264184076973345334906480679058387641057933030896364778134617322600267830786144062024101995864399201869579526442666600154378604162558323507835416385470113091791743842035291528178488803605121355599631220499782316502003358696203920768452720378339247197298623058570589216542171664648455293825995049547421290091891141550133345342449460306116944782944869174781322539019026450771474132605662634716653967660445713249641872909048790466263041243209682342256771749147968548192735246085710701166687917846612813498154726290780940240925320382968827046004063448426436952681424220598930973909459581121150382623446578438929;
G[227]<=2560'd287068414278541417250739956073008756696603323301776897854239173860162483966506780529741496396725935175248086354582421636445691994274515244852102062247480798677282212347607045500009409807372043007595194944495523741005033086531654766302694352896105351086212854166989475532257433148094590528421767828246216075474049262351996872323487423925120006753512089419502076888503107602648316943696147037397379717025729491417796828661772475962261415652771291885473869307392024017469106212002314681580660153159777720333006450763646858723653912336475237231727473532276624359203701196101088477227235068268606147877590409841894453946765815196802112067062788525597489935165492108698054796265203689608112161308697452406601227316990394375523911533976717118155297723169277733577743870926791184;
G[228]<=2560'd288866779301887728839407925443027419602680769892616641828102147264940615674487859030733037116766030422861340679746734664660735246158634162216309172284829376816816711665495520131057736657770522874109240284231168142323981352570123154253953316829862552291142975296716021837478502023001028744129446473426622946071893271594955798033964231784625080524082751667346938841925202572539182841357078692178665119358648319006988386539898167329504988656700387599550626056663611141213508533340971465645478126497785796508128337374252538553741663700518257189042764132763202072596133282015009005195163161256436752442596352169455680670976074628494722932981495146681326795465118527329676726388737459726094909160011958304311154276721934672037448972649433581714641378518507532095132949719294226;
G[229]<=2560'd261785543707769904112868983312277388623199806460468379398195466373791928730507219555183690741861799480237111989897204732361930675297402796136048727046975484478083535069853642170020438798377362695279349352465824374873793691303305736692198473333815374219755391546721593121633104430612027811093845778428064601861159362561512336567933791722057810707400705660437247754877121286860244779424497071373466826722710936831792998320163097568422853330556911215690747633511171926220259455141331681833458955555235304781538166792974398007403345311881474110715584270451296864180121764729558959807550499721294143375777608140927326279604546045490525624939546907518229440989769586097131599474952084433512524354405164307671584129347899809629651586284079465337399519745318607246962020521877778;
G[230]<=2560'd288866806849952828218513490920199325627659169463397388304697593003547991654622017398271568178489230080674809896702041936875788655801176503332919685854289612040004564201204532647457894985939097238696769006242976468575397695540054692935910927830217167648478480412800244334918469043937020004977175817106785335510373064653912570094649598574810038897329547464667705098729068568278620799077708822320827148362347785460275432718762359437740089653111767257537260842189176280198833084598506016643730735270492409268423681386903619473437826077683590753727243333465234954715672536385147343169932671963537885027714111214173766142152015788414960547083881976490137454568095518419627671632022273901553074176502915493005601367919693649016676409750503757221085938208916192762117886094549249;
G[231]<=2560'd290671811064569811978802878580452739573683385617813840918293828149068450377716379058269778311603485653577759387136411074311458800636025620211290958269076359200673873554976518587300901784513022913105016733483239565792419829418697337761713058886193500080637318831752464279926825062681804270823353773967881965575601290597291434562589828287238233142849387386348769304622899358931733406676396498202582002715459632279650835545584183724727425590368946188145571082426071037106723423517365001175792596666244812003558843827689086863785952024299444103334232176082569258811560216827609935479689756380881940804336801979635678837631050686959637858214488111289158639199012553543345994312317262772111371448320729854701944706275070561232886335093154062372179828344640604126427641379238673;
G[232]<=2560'd317753487528640956892551930831839954451587845253445056667297585754098738066703503374875883920130545559481078210584224401090736215989564219510964992073151201782205439089171330265542671686200279581500684783185814037053884484232578840096622186902796321408160624711208359760704651744937294092801459325352192546817444159676156882486357602807147607929163065595786725331329583928363839276574659838644685447299253389027467999933958049087726232038893072781756242283395789982126234659706312961489265536713768073901264816647328017447258342855513427118332100462104997484490017455429932792081763681812681704784539261398331426228645024869424528708362576531672746663443898700909178689698159556308371322387414505319796249378682863855686003737100880665569945753718144611856423952877637888;
G[233]<=2560'd317753487534946304820906196863095721361049656360688043871920598362018641614664162435430931830708568903991399828856693504965212544959383466165884895718453741421385346848173037885631722227599523659654551283810906167362144311508303619376306928948042475204488427239316777775775689843045496394615045795895881578711061400350525640947545302674484824494903291409950875540102316835509947024195755539246535576482675098516069508796038169119767019242440717328063743246318139191101510661876614901740743249320245868951820415520724603923415817212061325618956667696410530667415994850953001290518166060807543351511548426091572333246607163635310654371037108590041650222648832141901768257034933659696122693782035511041816840081431615748348037276869635349793821785413117403006605218923242497;
G[234]<=2560'd317753487534946304820906196863095721361049635716468789376158561418005251405462122663003173329234168634697303392638864890950382230740818640471442232066160458278742919226562859399298578334854099586072417858392104424115943901720240430965803992644703472996350633660937248386680070971644410986843000501442935564996300018319248043650681760421410419478717118433965551488143052474817262472153123881425871371511592416624030338830872422341560160853828155598233093237157815526229563088699940505526578620180320975921089325746682654905149818799857034365052332518219837466833676367603012304589853433019582771589578517912943716508784421894731527331778700406581776860738794881459247415367750368791270347146628488077764014452641173673163170808463287181381992055302421902468760256890550033;
G[235]<=2560'd346633115807664813304606722345925466120590955268164107553135241711410229105460343803143863816138695029930291239723535312302637638495044124732087536449118208536013580401091515188395631836469810850316147553075511721949319069553148550930643220329889967915600569231355664125450328722640315222661840679202924966417446113708606003191529569380907172886678585163212756314613040754864659346367499471473781623487158441167699411603218199376200332153987908614864170589957569611444240833587342549573344201469774545701136323338652570007492007079964881131238295181495944352300053518391526813262381466982932128071434020902977938697782316838151604982382278514466537632486895667201196481714321758120043181921612075545064523786754381365567572390308212203165121902376724600194714790384436304;
G[236]<=2560'd346640140671455967932643336770908411751187455794182028448973678353964023482797298370503485188731832292530465482229455254042050304078386972400869902770679299304822856912225679469522007468432740245698911053047827792055929109042935896014374902501522941471188820091421784304078786110325991206731222806939827524035279413113234632062930178537000800687180173013493993833991600541474094473669868649327846442535330327197126435959490905882159444189258946992308358041782436004994283321926643953323038817571956272184092806582401358485654633411959338726714447911574478389293414254649010451981437918509003840049703488634478698345306008787836598584268297268437438912512796113573605622967854412163673284007095547969272950786742212119059379165224287087202153895426225928443631880814854497;
G[237]<=2560'd319558903362283609294794437299319722185762739584393743815402900440811549555984188195606313626891260603197814920607576003121394303489926926962783142601883099049968794547520523556589463873129352473308065197357183661891312941126061183569771748396866212073929938394845888228381037040799873415290007451441673743220439490939734200913261902450795664551771329182197114989765833765773866155392427527377204593904127926578223090794259755792235158505541679684322663830759015795246513299056878924092980768496219532393913804960821204465577847011700559377721367440163092061523412366807876259234482453695643517886660274164727285562000422856057795822659649293467685165428597921811518129055526503923476355216420226300136264174800701747147429650723353797083882204476386219805577171934781747;
G[238]<=2560'd346640166504466532625293646531712841363468429855998473439919041122008268829779686344654337932926933860967742315936960715237455638003939934529922246944492410806883130005709900079757883578524843668608756517358187192232884265330685006823621520070297236380471601758142433337248160053254856086320680634335139985876311478025031408066592218572982812168465085146864608356385055426811620824642919508471755708588883144512069090454010825852764214234627144742915783705528474575094836439751897622458161123903891661410175657853831582375333952348746504962942179155671428914631210780067538504057209630560124191573661382391225988596659693947511592739096885760250811705310396729305064745074139800326145673627109780677917452549070340025726283455815234707746346686413927571647888032807338770;
G[239]<=2560'd346640168213215815196051365719374220388627347852853552644359060687753556732950158243961029396029608829676582315342786364253307311707995726316143220238164217552882504871426653216210923417635116356216300259341226728323752756515988020089908800583133769882002305705815997246694736807259005644810293993424463453859828896719258813330761138356729876818098255189609228681769148983275076458367926216562045993545284621589448625689425081855703221619913337804236379282069908603432800253190854613661346818945047937842541544458627744053041432573770441499807761924949877342047630626787793567076334380145985654331836233056100879607006855615221718393761621845456628564393499196513478880495009748541504655838946882565489486924149329614945224338474496628306143771502965928328517036149928721;
G[240]<=2560'd317753487635831871674568336370618740935843270893601456383635861227088704390905521266074136399920657789827050027267611980113682219062085884403207437633305100965553486795158684853434026131348595657616714499034679577976465411444027125149006549715592259011800939685759052439683104235929200919697373268882929867739559032382467260336401247544118387475480309035208334159245626582927515076914991292297606031910074626317934512679501990421958683353577979882954088804125217824967394862674942637028472427928509381330807794951043156962858107813777028661905180690624102673977987041176538660614034242406687641303702257310393491746007163905012451919800309284803944197020300786557276218896593175454115824497690487473291623586489389529042371087981901780885628316406642722260224350527509571;
G[241]<=2560'd317753487534946304820808324982329514156719573147504920358151399068033120374315371344616802611882374624057630365710201326569676981855341487030060444446368820952729887121023057154605969925440708487967600213777011719972211779674900974406968458088236443603290395860466677315575003980894797575967120367626874995178456679678582066729142919037304322478962263685159002608596660491313120648424633685077528786002072308887333586007561764314226284503269231458760815522904016547905579754044129311748136322510782965768506460331498522311758402524966210302639771004601137349752734776941326371252117457334057419691324732158522537777106590812122867528578967056912407347805582223372741400785851007975396336618158211327644211894253016781540827960406906645773006907962746808898721823293847330;
G[242]<=2560'd317753487534946304819340246858682500312394912349154612989669455014900130552183720147209677894964172409185024239633126959293371577583395683214086183350512092329604459074647783203211770521242585171574889328885871164292626241925024620533549671996179292665234208426706839133174172998318797910747184693072469850736651869997054445390726508268397316137941623846911495261140094586437988762029128469892875709851984524117477187656262586681848340544379477891131462512017365746844702959026423329827764783689904050434557751054103978105059228956263095114171571322795845814349200824992623802624597572461361474421467547679452189602883858390198737668233317105687185316069831432787729993103655122376390084980610758360663758215835440767199556212152700981328572734424545837325266493014939171;
G[243]<=2560'd317753487534946298406774596573632681860880662713374825203871784740808342479256224383490876789001923965346662407464719498248229013804563883909327895663744073257202605620701626824782375838976887714090437738990040463297860401062140287858180330514917339878719351740893578270489642361690149987658329621651518720270408725944142793491895731738806423796266323596575941846561487522741451999170403814957863916161747592046999180566876414934514415818620314173279381941227213610461660284818447587105481428398949743542031286516793505038738201009897844636228089061712917131839003545317132736583541304168076122494589553670217382858973755309823000948057969820511085062914810482104112060642698665030366955860312121342188395450239794470151583327323010381989147315266794368365131797833581905;
G[244]<=2560'd317753487534946304420022971850474722804381029319755778379669490570899920204618992923194716556560125348442963386345487905419111440006325431566984490355763010355828206362327959850109414899273829977298106591487092451160817622433250656339838101308683190576874259950075995844105683633960763663058256281382573025468675237397429988759605315216308867362649529339566646723874444055012988363183046817326810117471566008255038430437334787244096836214645094845641778920094427274469572287693220829736414222469787905024025674894170464259992830932575228435470799811620966493239133460326513290265114911647551278813457323937485605847573796587975284165357031052007122396806693274698920673498862235505670861500106301807970386792186519831052426552449363148716418007097536901220543001638601267;
G[245]<=2560'd317753487534946304820905814556893761859029617855288594279009145886009901709369308622628529462095656516759098274008764731582372613946352489178844898998773619428015270152144715196667720666256535014413719079539025326207730937683786939847319454547079187607084715250428534565854404511291146873707247942042411650475008548721035830765976685773972114412386612513374727295640300572357446689371975902132517731933426318449656646968425137504644184808968622031419965731894491726124740795375172344433677109435131233504183363752645475637169861777767182747283646549936418238570693907573762437407070721955224774274705412386659578622700917643571198583053485548799656287692538970287894954889837294957684475354606263225829602731872275339409344202535018003744408593008102352424386800378974561;
G[246]<=2560'd317753487534946304820906196863095721359691411162319281936343002134538281017069286086342040967392207211700730031845177039557111461114168356536906915049938231816080135130069086283948192754105438291879143991277899250956528912552926324211430809456420973956867888566584731121004049392995217562298725149446923729841711868498257763605617290080207575916685124727218301456631097865278373387964491271058480159273154941775553785240285333153808535068389146033259631458416781692674883569980638881811122907868913954090800650342120673251790044990011730968404677631146816618757362457649337447345795983223179291498196717796020625773739862873484213920786270523110931303127351069980998168493455851256804520770282666950222772363552742415032693815188888216317983034165528191007038329080533076;
G[247]<=2560'd317753487534946304820906196863095721359691411162319281936343002134538281032333122924762352780547774958672088107546660768234896559746418952852087544378346167516470065611605808685856453589435297294020594679745492849145929085397105062626607936576671475958146060330281563931301352734366453411164959458706219937018553119786433076165469678526112282032115204978782108316890119066578133779039461800887310167527660252551105765215716888166981071965120291626602758516319669537714367142678094004379342477666789700309944572991717133095038019578035001304789599805403827336154542839827580332645252492260864204015747463931770414377410044377558021388400772424071091478366449495472657642097515971501027596469258930766357080708905364985561036198872810527666566119540785050931845798052389668;
G[248]<=2560'd290672196945163595086007583775178341424637251958871203582947346900691342953243384311177692285142473398171733322643100575328497666762766255183903879118342061946299668795787163687125551007788684826563863369366070071324473859490665706484297738655764833093756949352275275726712448624901628979196296744287680295962213197109081716340858398528596187689332504857631913641991633858133551144985034472607992091806248964257010440341555302444171257929477481295093318861142121548583292124690051819819164267600126417771212537545594154930807242507862523878457874005786583216317230650362905764155177399280325065992596229417984613256728800406283809123753750282618620776683035328662971130567362960183620897698137773847726582552576162889344978729510734110280315525568999700564724053157679908;
G[249]<=2560'd288873418594045513645358069830705190882746072404512820394964922756526058960857841996408744325414741996326290199134598982118605957512167641427078468841999628684952506083971873341382095992543175595001539342423603106402141769262175660269942353177575280520062709690290810530931824217454456570778543629861913476682888220206542129956960442068682737189969812661256304895801367697538288330567505627552600781444209352008402455005221469514970718731539764859854115946374958893682688642242964483707932035383832955992138219995612086563510000416595560652844995374382159547876445577406189239800839916525156336861463381393398707168158870610860829120018014063036496425796897962306661355082558465660582726076042679665265371328865564807422323609134193343801851889032115069791287450515419697;
G[250]<=2560'd288866806856650618376266149196992828230901344769810195070124475989712440186637500730734432101534195472004997871028518775251265747544649870451286184992485164031548756069403061657256857496299640980041625143497739594619950255640420570703980138861413258274859280392063837250266605199327664431728121142458520929327180991347831036453464567616353443904419732780585960208790698405181394309554669401493814517817643569138155729757278241806561789925158442646903592749769288453806032871843156016653220492817233137670714543281559820063420688355915254609623114181650272240940872584298250532896624004947980742121114385893588382425008061067839189173753335051882386007296613968225044432022769394462975712482017742420480166353550700218601378922666336249757879453599689110888671493908406865;
G[251]<=2560'd288866806849951186200823815335556125969617539165001141147927011766392144313567624522756775424365606770862116583012218658109586039576554475309237278199426280520312948551758542617425841852576098371371639717010947393981796986962709432648464458750285485572003246874463179163896142377572229455732121918696150572694968446348816028811983574478132962550636771202384336176327129958193920657738177044644395355980534719927466341620650316491833618380566944789403610568657869051166447057200031782846930686262238710413159123155711556989467434347676802402382062822652404843512464914085126276321753666207448093739604772598738459604277194896835661821822877036377965017500910325930511748163834008971185146359624570218123809696433985930070331585686333700509471212581045651595822607927087110;
G[252]<=2560'd288866806849952821804381890624925449758779836803716031103896069753290460417702851177718761572095211962549255074068860133937201460473573320256989675438809688292702885342915954668867281977607883058418040012960079041133293052170482530438462899494756124717939871203481390741657001121140849132867871622374949107250071409493313486510784823596785141884976941862953621535351871185429455347669488367046925854843915803552924772241494692032347894778980454883661405939941733447477883783995918479413246607001792351928681200939283567586659519125068430620332128686904532137188340319712287302327390958505402277522126900937457203434911202866319831993620104420494816639814740592468180094483138325045817485211020435420019490088249368626774081049883400211682698209248081304703811250113503506;
G[253]<=2560'd288866806849951186200823815330450196363768418821084198321681891067064587276912289283259899764264629221684649644156498581266918122102141864141382482941227090930313749583511135612640536330685123973604328988799195212336900714891711925259591690416101148548207032931299026272440678038377953277587297870535432039183763299935062680123965615682938567645723623792161587359006901414654951285298187650529703658232532234989431935786976723043961190352443906126644276737206386116134510245500834816916667413572646429876328625185588705312694440689340494928710796943063364606201433446756870849613749569715907432843655390652847876483968281901340512331561967977786479116901220150482594992951823738975707658421227631903800634850871536158445280195316065202428830333184653913546275002382316544;
G[254]<=2560'd288866806849951186200823815330087019417901282875133422202822514074411421053343516317351130774691181089783900146516070602244424300946432575600732137625821836791731664863897178260620349123734330567590029973489452352272491288814301851113077415822597734217702145266784378168987953467793880761040144759319747870031466024841185001035951667191331749134138413444979116736356645505600517753531012645446029333474891183108083838709254879130743761987120557729807086656579377826159342755069305469901082035384435616035294148824583400392843373480760148462843606794784983627066004917871149246363274224513327645220108275123222281724540005808811645296724462343645112943725356209049647558428533934957557452067192303584777455421964638968017256771912803224170324965256013245337523913887843634;
G[255]<=2560'd288866806749065619347155558829994748867785660032418629910706144487718255251768009000171465173196845750318567723503333292919654841072644995301068276718893067406885654845649878003199110268575507863436117174678153023009414765815635840490322140354538253990323428488285903617767596243051368726311597768793390365922945896944282275862251727997584913477190002505346961584462225289987646667457494613490883819952542033969923250399555890751272300176653360103681546221099252643721974300363631936451004418499847037608580126874133927166599500322915465505560688427460869742379280739176631041368552476265595630861129233885179204090453343332018922204689518468896904774672521687949712839813872669384920551696492560168518723472706566523718910864750895448458956664466314041332529513991832339;
G[256]<=2560'd288866806849951186200823815330087019417901282874835710851290227357013897529629086850209676794964736857525990266216064196636826112978513343536275708516407617657660936699680802974935273879540581048092057187235141931616615117137843287508196531514150333315950483162648904018868449776889828092277057153508940594067486003252567631272596957934245916705697929755248001517419410310979836070602710699189524623860284048390972446625442780858580595146812058310163361517193481411490352770422922190705914915686499971545411583048188484504013404076475301795160158129244902014854771954181712163475970650032339114052664999350696255627012868753475922969824934535743135701667897892052393823233809176031582040282030237779697240296355562733070846656035160082924422940052749121503354171671257137;
G[257]<=2560'd288866806849951186200823815330450196363768087218252565323162462943241697267191316678794105802145149376728691626711116529971847148772814672022203819507979812279555678138754820737372401219529374803832591505864725462202072959845370457628697374952150750026498331747707118772727135613790834417212487435140499848649727295518934856955645007897538201099225485301470186777239756934237363155436448075095359818522992572796607091988975175926768582967226411021040975649390894817484626313553809020147251285566279851232288735333098916401566393676993567558312039010496339500838542127768662201392829839009491893323444203914083226239815063655692592938485251388274507334717947473502045031072038691953855491142172364204782713149344586362310369255356493821863221135177867931577168131515416691;
G[258]<=2560'd288753968354410997286513975322589850922108738490692825520404341418666267093450686822448690502813658763268228520147974815307506058679657786996564457563092310507403865604056895270121124370822756444514703974924053990960680997090943306438943174194018195702529412014504704121608922437253399981436031659688793896641345343895919914999800619165184321320426172154394094478307520903407325060025374749198228025131353672198047223901941852815782533748726945974538298259777699874418435650682031299982534691902027586160256951274858181066692660782432029148901455077913833997285866894537506311478946036425282927213520096422016648227514656316642422658301678200118897561905056726039585869353699458855059530976004672702581260682005475022719544634256511709586237023107243344150966702776131841;
G[259]<=2560'd288859754437674576465325184298362679477532022423175708434219335659064361739247938391509687998740630510655911370768457142252681375941873599687851934475871685870353703480936648600779700003862469179351319960607559512028068820741358480943990702798712629238921324225393462122990947718579246022787890074013317194046560997445357938529515072151951209961066069689193936848372291531815871563382861168544572461665049449732252279462458049804180794763473545986552174815854515423837023586907748169539636576110493961840981161925627331388600768242992815911901905872005553670373614040487150730911176555500511704298409921488016362284981666128539591290082481563996117592418909656206916845288167004601322302655038233506386055285563718474381121224185364824569183341226992872126516133028507665;
G[260]<=2560'd288866366074185540084989624917427652937348192253971142444963996651003723191795467772825051880157570085497946996492612617910712103914352859075289931776090975469258625873647002236173851630573344808598352377360094002072462676490070713686829574755566707413675342381883337800456998634815258233605929464435444990912580375849944482720047455563001001209422001214231217954683315622763910400308306614102695112971057762170517607602842439323256627711807760688009065392235848329492786876857048423077042268528185054258225473855986356304154489757092021670584752301500686759815171058312317444270307700995173925599977809816020085594414466663174243294722743821158898250169502047637883954712963969747520061803127952465890353137809263046045669230406555877871828397588943330114499510460743680;
G[261]<=2560'd288866779301467372710168249295366491349205432114369159506536445585034517644044505990597003182326458313939767222387229808677520419843077369903492395545653035547824780692874747835242837048433751628447454702945494360827998830308449564652236277322395561633723276555898813924050351383773596588235046585780449510605614011418390960770771253762821370629772686953737074772593820683007090070476606432602710561487490349671548074754043622202197116576996738853098891178580346514207259494905481939606887508561915010458508662357840369301111587984979647190504067934702301596783739663781545361641707803778584373780393532396866088576300502934674811694353498004122334508193149894015152068089403502085978179353519120177103869764756134316724697491034083380453874087118458352729928863081328897;
G[262]<=2560'd288866805128197117514587047170309173288089411492498722280452012207287841401659968952497575416770108089621119765774618796224837792023120820273290504443750426080893154094256549263357105037492329908487239769582475169404221254549188878952884448313991837377141947215722314666541589937132659827150521868631066749269107226860411034930585098936472246855475348537265237051321542521851195008239884214093512974260724167154896991174739842682904207755448885106001735630987723285585023173838145611078717632234335410516673032620744058761830112299043558947836354826488687299548757204274708733835191768730933460460449884244235781359834685015840799716343749417792326137484571916888069517542850519942971490642584463769670061897324925509206212155732523981557227402477271447986213861111994131;
G[263]<=2560'd288866806849951186200823815330087108410211570320996007621861642151374733975357001624747737359291639488807931782693343896967867928201506212027261417257009735569120094117393727474010032830033799144843078741403104088867405076962815996351445607197797762034070271580601588566498057301992181646997053680153103818410705551572516546616726820978099742121766519765972090801420748468341975759302383861540393010189570247636250246850145358025858368587461536542788076425206023728843685879842052303360575778752888270238207184698534283473986177916185914373923924622589285090289798531157581166102231772495065888046406700661050965689884547649244912042413545636850301734917186091924239881050003556612808256092177913119866526869659344615593419031615624414408878449460479277871098880355222786;
G[264]<=2560'd288972593034100338246551656083135978626422822274251894609128408069459470186683692279474419481195664822074807256602501602981106734659094959729417682119658610637440683738754564798097428747217992296632163317503805317405646010880587302980726873968512134772973930897304068150478422172583659041109837625498296980689192312435189829569162527619503645163484471112412403909398923628735832340194060027328686272765298823595857820526933850015833131447580853398230456627347456322057358937516685738664356525708916222581590094785423467901370177645156837906312566127853713577160294163359985262218608088931319397424690404876034670228983106738650793202750680463551968944449319547173185180857268151436873169967578570498429611866887194356886900834734683329427987350057042134554157048649823540;
G[265]<=2560'd288979206392363728935646414289956602697065626820539360300630215794367649882158704765439077552394616161984979863403359397419825661077741590252579492986945902360865170995459268876597790498091022080130800477697042143341453843391109848590905268587165358646458907180668407061742920161170260216064825319918225897464353061603182698521966821767102694863695279307793500330115247336214203302981656187266533812128583596588249504153144075796508065175618707534767019293101322960415184463453137414146930237731536892079409566035985797739013994292488351779107879274051958129684589421615337981105358299286351137433635245943513074298921744238856322858352327937571729802626797963665922639428629237583813298544267340668760318619286141618171256065448556913010942374479719031572420592174039607;
G[266]<=2560'd288866808571731527170089275939457119987383974558214811889990736112869658831157526617836584578962982542197840324368761559771738025686959391318667213886656993161035933091974972827903842298193004971862927999962608133391728070058482639388293771067728898391206224799602060667527060766200380769841010611187079770979995821309539775798128045154362257581565701330220567086728552341089926233741539036955410559729814625540435352313605278829623435502551194015846998047385139866344742913572763234580365416051886260591578843154024714249465510368648202461015805276408403932853631579183003190400558329541162725521174368970429697790422581413677528455675843923405449078834088628221405011238823373815430344808528228839856379754338452760219612299606734213181769683060444085480775699979055154;
G[267]<=2560'd288866806850371542729380766398837403878526764636698880405354821774460572051629806908208243964932161628903862107136205383966594466234518991217713763829810039049097782813832926779663454846560872622889655498280808743905164390183472121721809222568792733438012370137776047080319561557515207705847647740220327935731579339487687014813030115009946935348991525041279417524007796579793866130564634208841057488378099777998053780059135173317332357236525139080096423775968696020357330241692480697558558317638131954172660013889114464488397576224913878906142475667116336720019361951303563666021593140115140158474425595237983991668381262225155227674230761461546503942273983579541468926055480174805358988038407628127814036912031758339066718844935857753428974353912954388809442842254917668;
G[268]<=2560'd259980127886738050567702686988765374387463685668492741581269237612928300188544289184385084648506636025451550350289017322002953307527880435977313086888477334301904566662313435133386344850893739429575031195126393280935885252793107524791469693001074910667954726859593859337827640431173805275172856388968468163873997000516384164022348452410826961299324157935298407899820876060578647688201404839739811074916872136715986299843765866665382072809559866946450122194001504739942651115042526950391782127627733776201205449299688729933098037427814204440390501512556393877987248107001685317014031297806161318530204445991211635076598920562063746427166857882476181174970510003304744060698983887496647983036201211342664481043920630484489821728572164479001228095067700692986059954400207109;
G[269]<=2560'd231206284076807068072208925154137932499244762979111942031084592826962664482239202021839689082367403421846017800157422778836767745513475128586423627181519529100407948495094947936399429167723501024157897939754719846169382088915521243969155881126885214566387779670744895074149332318370099855829547497494537702356422968896106596595211605879502454881328711686562411243232974389030727439056990886967885760448443549645436742042755582037687890359611350354400477652440683847418900778243702965204253166863218223498614571488829153570209364388381870463212893737595274602171150241606072587081400303585834532550369858755260044204538083152557376212466653856791970864693418594202670523493451191068372906763228485665152397009456529149076990546131722747561284940659583078366900247890313474;
G[270]<=2560'd231206284076388353160458806969080815173270010969867922426591326308640952126204315566114774180626188682001003269345552202769191233411294597675085320149888359175378115136827975609519612126397528066749981550562019199488313522879065744771609349595020739473572099354691980745074368640336570958254560438580544826624359008894451467627990498333220698169075529616087067680820692456618470032535813361115815276247757411328045290197060101387540762584220658740356729212164680563080840734810974874601506426767866903444414699678214439889651667522772158815487568205660381741767397284113544974692481362880997065421010628365015162414097206795869559462558087648608323083364811682312091368286684564321375610843936956973065417706108877289401289831937419339484171633021250335518073081741743168;
G[271]<=2560'd231206284076386717556900373256709030610308385603339582079664494033135822954795041799202521645853956483294035418899958677300529169315666078520309474361505387453133825796889770515316921102273355268614370136431467070731413640964972657709268900787920458378656626867458919093949422658060739786735338348420880937362633227330405518084629399062766114447973274440390926297578043635288920053593940116625549932043684914930982063644827470818409306044374801582693425637551838044345904364059026429808642112399572703395439811234689259079474818695694078043115273941330278243969726421128337341030925304253930743194328097860184781329081025743971749962495718471346745023699849906678613274806921697263836330935616664118145415981202484817220426406297083852719897737706953518665711571351635216;
G[272]<=2560'd259980126164956170206944910402568357759739897830253428175450975477193537511214202205758539072541944510705842936295851007667956349498338884441766373585211773658374276291961896088670179244196207543280331742764411749213944983505639941838562159550318713209567893316103897570889214801604840679383399364426043055682684102759738582844543572177349048574551992802885261760996890371309338105880240132843955507327373078240168954020568152144459528443774839881613856581715494045710659091779248950790437998583934349458295649539794643485606172400731671393377765082252668401627420085294658472382138279710688357143215476838771712572587001684582403573031681807145999688873281490313825064781274753536117915299900290036356731109052330032787011040081454820081255164868660078505676641227313664;
G[273]<=2560'd259979712937674337581668796455555741546955857889300637953138093237687103141966446179436402153787085687687900759214031696076110782838035426117092126857459535059698871752351293647165499840997315596489933186102051577948155651180955562808071513458125679188909936151846897334798803375168817651365990073671971561177604394501991615783373792713511664197172769297514672278541696344882131997530748153966133720270964841078631506959499469774492895508082819900421574127223481423397205554442353955871233109078200217665086308520376671476481572244677009292611009618311972887637082362410927358915433548643792462754571171377837933669145274275101969235652226088620378995013973068134868703895719750881841279262396763658787669602267576026995896544600585236880107954586328705071952934292854049;
G[274]<=2560'd259980126164956073994873416404387771879767764713084839868115769697150106840967097548740624325058552166103961773884170574196666759042441147929355476836889036914885307465010161558289013008780655111844753552035785853738621853938442540851516865884935594753725048687498767619511090898233527840647089531510188623502524400671990664446147259803056570932913373851312468625094533473348926560275922758108745528109435709429667047534470289669479610093287967286971841244444110661777429790903676842075140551310479556393673002415115328261822164071689981754060754332370049349074751036844544623796514329011916871716601847963906082785218117536502705260948888024398213493285340904726015622097572284269846746741488860637493538949941211904735187033122704822894118521101243452115873519079025296;
G[275]<=2560'd259980126164956073994970905973460214819040537670920596115418876115233572016013264975497022760341401074898160582289269214402742995435381832023836434498918134270752813241479018343110618847102578326032908861798383711226997470467402070189841421695902126119601733553253427467539784650364553378619963200046358355364875833553991477187330633663197941580940246974020682600475245729868755589492200411392413799262023645399450312079331346621994753891190495309177756314301294844968722077346784586122763601032561409730997851367820522186653561049751777644329010960439338464333149758130002755632998914446340847614803496201282764026484350654261918434423867464843242461812404478642757107072218419734386667315146304506980348402389524508473834306966146423312826537282199166769833039757513824;
G[276]<=2560'd260092964660496262934238075663502775748204722563419237099712572647322759733495569420634504956713828313269241200588294461971058037293557877960347321812615908442662872864577076845573936388970808324745513004037872467000682419691993218281891067796749101998703985523906639632996421770375629531771064229539569616846315156104988913536250599360697644407078382454878593209952609356500333731542854933953894722723531379295884347934057925288042393354999776460612463025325802406853819973734435649675132961456141571725513549513963338319343586260679586334752024459435937797673172176934170848442098481667348776585404569324117761840824938503000160569737364584128673329367493890070735672650203912727238201833606486467690115823287762054237823465613133196128257666459911649360638045219463952;
G[277]<=2560'd288866806849977458483858624777375723557523307046579907333923193189318291702694349702418715838387540870116326564592233572951875095367895680569159270676212547522438328233677228936714241600006928960369527023511195327399097328390450314955582545191444686278130716162292880892038038887970019951049201530748756447957443742823233397557311391392338412730620520428074921245221695580678292072519529865150139156214423734906708598944285956002378170050282301444088488103219300650270272776247460470634327930047954360149340743967064497800702283916746999418000342347274250361558757705776818443462852701494062279982720190198610585924867756817068941728804104294677439074183400431185028313282784443833107945738681641476875289694369122417309562276796632136037812456326151775486703731416138576;
G[278]<=2560'd317753487534946304820906220757597944997666702310340914600483378251475314198117132096086744285405134186002470671315687952942109293653375299047967771292747631952511622235956735494338414074057479974124482479421944578103737956870170053665845089798971491212525254959532212499701505860621278977856016621834916902578354973162603568293732661559237865066545558278037241149219402416139049820677912163369051688268885090097064009528260345451479238509113959961625689136013404425416940046882273636659211640381953773487413716720830022636615616997487535212760470550775123154261761624887513545079637764836141726309058007700847133251215244580836182188935902750402764174201878356931787317610031170522585806227280085222136320957517731139542476139142262008240720048985358204430457456691497989;
G[279]<=2560'd317753487534946304820912313855664972681365945055857243956279001569936844099366033337668241316817217175665139972853718176074279014575419431578537422048196320706055417926821023614574034706568674974614136631648404596221608175974820207467028267555528140961658698132427384663405766448321310034753654001299093535861317617134597920700269777586402765804742580374480625698008757031604878045469072656718238256598834666804568019829063199566103401546202714953006330527039606291238932241184905536914134507181264219320426675335728562553113468873188708259631676288272932195269755091136241174043684121525167899700591697436303115530918449321085962392848514237981221317823152159711494164909457159118889760685712013620910724509387692659857120327994901953238397596333795647466134595055085312;
G[280]<=2560'd317760539947222914957288052913274678562313918517858218355133984480458333121390479808294016872729976557907709006443464120715387705431074455934692367292110082219542560035226217331809024015956384077966945217453304500626804187229432273137530723620886309524665908614024640995583707374822529769872825486628675651162789281450665901937847722151386647305100592579633632052938662111480545865300285439156431213946982940105240071339966544199331454353257816570767554742353925268269865411157865026609722798411503806446699703701728069690957341476049973513636153288921870590183392463005416064044780826202857962024219700911216179681651247065294687131931078391051075737374745921831795925062836938915056991209736072814104065826496040408726739045825806873734943845190185919687960867428049011;
G[281]<=2560'd346640168219941423440988578396104423301481539449802853021534121948074949350697667340640358627512172922524706403888604697671410056553996887674398893406435558470759534212475969434800666494988356339875640795165506646675661852933549876043897486022064776921757223760732549642273044228712720332803539585904501758242942227382639206070249380717303530263505842716964842420012081617538984756755181043891394945233883686873286216730350359184036226038064648804285405457713336720612472909227432506660328673921646298071948835036632433794836224833587756170165071126054270526236066095269338256471831463950947716172142017924992900213862853148038629780665776331929401485330129688343156941455923676635446719152277845161014505951728248590963957286883190229424892514648686396088597128139911723;
G[282]<=2560'd346640168219941423440988578396104423301481539449802853021465111213903647704711959299071332830110145284250048598603537797485109289721953132522718287983672211473042671024248976863898350479720367322640242297407109029197988359681530744583600477328386255891991410114549736415609453925336769095809245479171259470162560156618193987380835689880864010880806095006626072514386772650257375035620476340993892425927682048645632602627204344846695989160410369418013444044171908315860278023771140003510715840110797369115120156926567547661710960400918175769715620380559834642144919213624399497743570416378709920093632993844635664188715098968096004237927874844544364546822777390816731290747892815904189772368154952831488325254370450544466803207691421748324666729311428351386061423017100291;
G[283]<=2560'd346640168219941423440988578396104423301481539449802853021465111213903647704711959299071332830110145284250048598603537797485109289721953132522718287983672211473042671024248976863898350479720367322640242320901313943997992422655923442495717101394746904960090762313768277226082751875568884825620916857419778142904351332144255965788973845704792009944449650600585740075454214490789079052852927751649388053851954882129113600537121492449426948123271526107517119031977250112002911040867988387955967284660042771022310264683558193037534237404426185709226116124780655608367726673271417583573887121405627068956550485834352145776917008927007952655436481757053458158182196978490926329984014758780295522293335941389434837397800463249738568758545534885691463169378760767543361707338650976;
G[284]<=2560'd346640168219941423440988578396104423301481539449802857828072237613142319219053929601647797749302551322723410724669605205868826654722004404641882941704886196802133294319660091387576000785252372675769620273959810566613838198345547973166811634210712314730790524621801969710371264119007869411731703426914684768365699478703876970965795874236102534359866645088235844016725795574074411442640960378703326067820707126659776717645001182822625446247803692925801450752642460711377900437404074449107369804056113823786597903153519328263884874518298521278094249492243232035576679983679021611690308978628490053874712688405030396945165036516332731163641649252661516248569509804585764562474528427285539974772027938801934551346736290822384458631307610349157187128871852807642983219686753287;
G[285]<=2560'd373721431362124347147315811083300081371909784719318700913771655560605601436611957779092833304158640157070309326555537447322635609081726979788141628482095565756166985381068023356502526014204050728990460763670842476444244708245024563735308116297472694814990758187941658269015728793364311555505837576614936148720628953016414633904466658782800323609844154999708400226254157174630735365859050714455038235300406222203131958752643349355368737472355717870871871066055875264434821180691243469871169120532575566769055312517309442180468421265067649102681094460294424936177422859312552802169134157706994168119858130440506778592755907747962973104387740012445813082052417973885824700432577991174320021994146391604090939432443188875801191616779885087815089899926701437160024248936389376;
G[286]<=2560'd375519796492659931924689103878934168040649160381747487687938861325036711822610886641135682831421566998159978053986320533553070658359588374738642535909894970017282729321243620385424078034155908460136200883953777664097027243730999661533388438046085173075770957989269014502769471846201737520969337562952115274720104346092211147499718757276765782942107702759481148261191316162059667068695560921864418037892739364528646834578630602521720081624752550728141379959203882712079161276933199971175249857660327923627176140483657985128649760473959113261888932547399212337220407902921550084348991386257208302533625757457463848021455792865405340228011510773538101657182766096789159338178926569426713009799386503507069991070272071540676281316140268353754344850988814693553599765387806548;
G[287]<=2560'd375526408129169253927547093925976940418107761027565240581595152154469300065050805907896611124987064866206272089334022383401282992195518244198611474369284763476946661978244182143014002746638880670967854573410808900732338544526253774296211561890780289605955600115986566551835874849506019340813345168992269510851534242545416969818468898411912994829147532935459167398965413905361840671038850386373076316725310708860341686496094764823389017232380276039130607389608627815212470244256430826470634941368238496964068376733362986010722351160825861205670523467377835946453894587937060491560814926489048485790256874471772574893166168862361754023038045383880981594811767043670727293266822702971859669829885379163175211269913123418991224844523980442641124214546100720164417571813667636;
G[288]<=2560'd346752566141485464343242665695923824268393373271121733154215036415188150942111237476568056988555651502877292516566154085675030597451940531929561151019962591856081400197499188434813090127755752407478985185912082704958526045490450496172615854134765043070040174802726516823701409696622994577140524091967100593695286213935404563909588255378585344955334379961521941291795599318146601097635443666797774380479803082702967271485227572673864863232018062104129841340473692508332073490680335845438834735389686970476617146565063606128344516776451195915115886161177030934888203335921009403560502864511979364826672174303685045255934832397405640887609227234827631422017538399886280818982058410149786524282230174829390387930537479256320361267015838191222832130450155406652940355350652004;
G[289]<=2560'd373721431362124347148875644188459168398915927571499015997451226209997055906817256918814009716627326935660996909025068783668568661264818528109737545023349838709312108497881808517610875315077102866806455656282182622867159621773205120013674159340918952266639154211703449866172367108935249129534701496433695974648463547385070058330865948831677421080417329874530866676392928063595284947805857141795631461542431000010866906869410227833577609732237756191170101452118778470493287576501382431627149370541121698987206082968556190435500160550373580335372449243103484906907493925033038841957875158047034206102096114565088907822010008369583964384955220055093304508193038326147156480505318041463901712559953215342688304171190954457169084196441202122427142802539277079827965770405733203;
G[290]<=2560'd375526408129169253929113042530298889789414982076551930409923439760068482558632605409088302693514892441681899446549774963415278933728174823722718733133277122899925408933200306429203324529774208553795836072766482884935256296646592601451516340407307287510328660532192014204686294693703237492755042186196829262131189339773958437155201666885207322569984255419163719408110157165959662529328158968329878530969674314401961525035110057702215433177642764431926021922562973172388655670355180171115593900576704401518128611247899951110583236493759097901609846858125425702599307922090693384160405274564640469965214352853474146288868734337715495623407051449659263710777081761477175221885568237414413200374534204160464103162698906228401944356186627611169387231773751923585379576584521267;
G[291]<=2560'd375526408135474601880956561520521519737196886325436384754235895324169030419761988665777073679377503397863365000500314179856839278818258852236456209745357574109791347694505947546612741494001113573477244016048691090551571148402015366277436221967841990349451231363594949092508342610167637097913823182453591819743663742123432834145006006849178067448745847287893365070539403770353033615227788248206245752402313832896914583669903408925381475896483315599167589295581679187852508776186095050920406230225082688654425070151407319823516393368413080015441510878151796925939132181684560424542234523237126457301491224043222146040043131664903305496838223187765234208896767804176770262446477998975984108732851532748587819597816292557092793309817685941516003964956321427565808392238967650;
G[292]<=2560'd375526821363150519127485350980216382125986857065812555824160204053813673185976684729430719540720812727115883033741012718423631070949418756474964988463660424895977049371519920357857431938322457214483751608971709800251844880473113018456598191090524687287327051083366419554009147294276221383185891512449670818739002823833796718976821554780375863089413857190730650145249048145067859929811614613724333310628566757950105028440238235586201014430770878956950307724126193185467645603751869651609597261867181980354464632313439806058325102203249987510111589251259764747541967802903133155882431037038854735477715992162923697149266592144561477819593051302154611328876753704941176678242300583980200443222250179696377005058944232976077237706983266668015207679053771634598770250115148624;
G[293]<=2560'd375526847189855633666559015004202244124685344680385286986908383510140360225359778383926600932986682321432518024195657998733254571311601138885626025487105466667033324887713287341064338082346473038203208001683532548277007853417794530552127865957312009935926957029842819875057207958793591223400182410379062630744912375996286346595764920386935924647818052480677703445172306084979079839975779047316927764803536327712249962879786437287870577836751503167937633065039484773980870076408247758254265520475007446235604381450519477738896696205924679890065361908690446806694768636208643154491413576648720265490914546825679952177358048049510425877932366515891837035614163693466313678732028027854173951844096633233819220279493721941519726738860870072719499360753542541716231090047058528;
G[294]<=2560'd375526848904936542061070959929113125243186798137565353548021048829967726407253442370302010655678350364808738927299958539513485699262617651380144820295669769748673247307688971112162148309042557400011196690001809683950963517309353977788955233674633212980233535279697739321895407972240450244800389160939083301065222471205698227064185071808386007682375602480808963127827827319258723570115682130744722535488360548583472724555560929212270949092463344501576238891435410943109365417600326084782615623763794952943378901189864082705977082980265908197387506996028731988384186730335957227184960210196982169409659559792641263085569430221147836016370493133950710215736849604800896202176347209894759097897391214147733628067224751341549972324253546434835495634796314995681457964835025300;
G[295]<=2560'd375526848904936542061070959929113125243186798137565353548021048829967726407253442370302010655678350364808738927299958539513485699262617651380144820295669769748673247307688971112162148309042557400011196690001809683950963517309353977788955233678694581385293626690807966578880572000045423770518189129141529182506889641914886363884940699627779121896113098559384576008483339385082980139506105944585763219514486311406304987705835490695270135178775470887535871887463285494505537758708682353562861653222269689184345862328957696784531518207190004650934816268860071320037860839742985875405788509499391853860731399407327644136907457452417018506246839689364471676828783293391568566536779728445558006788436703616248320736729443063562580835710037118991798002969599137251493959992279347;
G[296]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374651378681544973288907532252361076013666096184460625399781827169719148772977610020867833935195026032158838317745569339018325945531255002668281394175289134992069567765219803847188262940875447481211034710193756054284083414598378595076781963247700374298336694176296505078631449050348818831928461717636340065956134262017483659170151933945715108224488681419244071933931150853042323265650978273513731356627087126287898286059351509987632559140499298677305962929838818147595068890991662436475534209150685066187941648807146812574275743099734355392924225754987579665208658400645453072;
G[297]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657039402917386276938768773586998417597159149295475539205602899633491245905579478605941723007278097492554777844616307919064847940564548905239597325536668520282737166849996844511351964826138914747640122895995307320016870068502197036245286120807295476568815801598894994276041037261027836511059993763468117425239876393218907732926459438863983131164352222629781775799407383010481503767578556193448632884110341213930884539055417183982716567472085382810774105605869408473109007752797907430731421725926151122437824997318661331409208903707680152685148165780140389235223615978646784;
G[298]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657415310196023076925218073824657327233206299304039806276713006698115550748452450408862943291697040146065178922830559647560969230955197467482495859451973224166459711018420976279694516823698429323433530039251591952575900210307235613641752465367851727253191851699472077409305280991582571120795226137069389773322736672190261405666787114976557665197863418949667621337990339366751316000811626871960934573522331479894904366433421361869381485268922025878625569448553630149009730305105886991972523666412207998587243199138503237987206745809923012982271764569890465258721387882486369;
G[299]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657416778583830251925165141403710682348972108483760760444959530553836739439244922954968104308422193732422518963752120017816958167695556549816364270565742410309470784660412881889681199867100629442631847299548386998922026390361655070466133948825978186902654570632102772689301682343569086865765406792236428652306369554265815151318186400990111638917134098570893080747479523738592761982592396804419497563137004095859950674641000457406655072687577916757231629033555527067911899491646265038676265057328732403817690636942162861123360396714729010990816811272903091609242289207268147;
G[300]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832508357113066119326591458638797904556494613371008095871397715574088669727863970555507067396872967028107198711476058364374657416784340807954113454800604208751712865204558928267058124904247147456990264372992380310034971286143486938080533102542529503327138947648814757532578551161019686048354786133786222001384160223697637909504794077060264532835110628172001678766657792595884410835988962785442484033862763246259953755021406557369516173528710655921289938212232047277381545929758557019142581913197999673696274658008760248408734324683115655104846805822209271418042555022580056421488016602067951372133531777161637441893156009484039483856886812587697160892150254082630030760821250750643413001349584434;
G[301]<=2560'd375526848904936439835848580223185723368693707248157100082245105822457809118348087590095698571469869739337393181350835846302500224783686911464102222087831713236718483888648648631327416695137378484303943437167632533436369404056353111333448490539670071129943162283606802345088665745048015127786924780970649583853589505013895673343080842715588017591407115222790310215133293792928570136926696205489051728739569848045865499798068798311719780622578545671205391694619176930945053443916216794194576575640935047724543922026320256350274631671775115470674585182779188461636508280767310479083835752947860029500106679091560263950992563802132672406775920761465473616174596067817435358563544241283821325856111217832102198206781047347664301395876781295355680520868178809398917750913118720;
G[302]<=2560'd348445585661867949275853091035897794748149839136224171230578940215639490914454518039843152578157003246839944395160268608908099119098937901568080856375832185224327245835263105475645818408940631064137985811401507183319003828630070320940670992538815182664927142209200341533879712428861603737489947019917294894079407954102091039928873948157492963581443548492567893982982356051941992225144188123257489009060485290944767822471287531863836413681645623054904008734210991128273930638018544563640090339685999565385101480400222529430565001016634400841513509356451632150296292280938034492404634630877764736980979315890165616368472431826203441893118936315982439421717211475425951619831364761713253575643663325826845652598447060779373524336865438615150143731280742889588358762053643376;
G[303]<=2560'd346647193090432010267956802042950034872640746146855908410108296943834601004200864980790016116858921587975876006529338458176225161212403691009675054665081370652454221438876407352801677217745456613387348009691088950666360349550538333011341841793823262495258206632458665130329923913735046728859917565057734139732884660642238178221274713474142907426250618121605812760024984851743789945026985221518093709696053546609121753118067284308696098338398792181791885601325967876699408151047158636774805062909631684107866471220203442898486100405168062724175444223589038196604749655612514716518143723221536677221165708515203073184998066923632335357761155760454625071730899649540755308674863195176591697600326357032125843163380892911965153724282013672871182996847539952878883302471343205;
G[304]<=2560'd375526848904516185556003642638323394220460995529563298783069367865548540540349160638377207829113661986176614353811621435524714399916059905156634154703299210657778061980939040198585328187201013062808124396403385579164021550406235405817873845010591771897856437457259832298901923178256853356240608899885677067216524323191963235612466331177598795013976185570779912942148109393077897140686259594937430375554704815254823063487428757260446688405317079478717470452528636146863610583009837659453994256362719140015621478590097671317771784533191650175625754629408363481274786482103853738480692456232234736253023019342794975734790470726605526275942391680070703455930780853629796144267402489074736213949005991911391054649860122339760956788252155173927901276154887559840521174484821300;
G[305]<=2560'd346640168219941423440988579889146211111029311278590752312994453994577135627304058425346045531358489929099089460949648771657908088388276447827388096230993387996665576942285140162904845669076679144082551440924803261203120529727031550144180410252400697003679722462655927700229138830688619307145970714505889190260167892611803334569077628999798999118527912559814921104423293503369532790182301809001769278861922074724590017437709155499938523209608720739349071930998661622215119982818015656217160796918451149041125184430656280282622721884277249966595877347590721555959079009776111936730352006166178532393694915652301833499124234522894920215025044807607649801645544756647582956339970950220054684215168839090970174249005627237546778084555195646492754499612590443539124935773798612;
G[306]<=2560'd375526848904516185557569210424016154361537013906935453260438936936445110651989038083759123860745836583806238287687290754724860441261589290052941820937719859614427395109211699569844811125209627892307266329061090947079342164810385520301054401171004877333155035255009624974596020407257677440066085636816585407049769528102693667499570248736894968066906632355349270242131989853521229533754503044952323888505828428890230910040296815443317085738834319074833320262895604571372431012870338959089498350239229101660937079010932181776226036483720065908327487847597036024183673239260232959550667155003741179667665692491338446566745497368985127385125091823620687185653570175214675605957491090420487546726263757228966476187644150886711650583877524631031116201890775994398784957363296147;
G[307]<=2560'd375526848904516185557569210424016154361537013906935453260438936936445110651989038083759123860745836583806238287687290754724860441261589290052941820937719859614427395109211699569844811125209627892307266329061090947079425960239853770036559982984385467456116524404556412408359775083834176693272294669442183632555229719434578127044150689959261320463959677189936808156472337284582669921755904406810156970278640654458130389428211363370876306953149845264023164833557099384472406240629086975014115971819144211885174261202435711982559776852635481429865692633411224340531386240649435166748532315138750767364784608730233118568993117047128546099487489756895001552861479218136295005469065483952796288394776448079727294381945963441917392255229226398973495563490376116708336716125395831;
G[308]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723047641974943817133278623886585272814067639075285614971820383723164074045292231231462044710139670073055070647604676300152927754721684453797438305567538907471867202414181885530215426543722039371047253171835550239111731494467613664552029369450720266184134684662980353364403277553696804778779132330345287988684121520232463922987098291955588043244508765607847995549332978622459149880434332531614132460930553048264279533994686950189444704395265945059760282060303707359988458486018557038977384667825297946669078017425465788623408493459748555301717432;
G[309]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723052107496729862771239177481630005718846648118712958013050939669416911078729221903567595356438561391772021921686877284936732953553713683533859010177111371927686458635486087837259074930031822078156784921774099477765045424112310777406988106209590620258513102241520343523564805679367935701786885123442897082851292310343359021655023975668526290037319771221771776044698344646350459169777207587404316732783000392782990835614720959041136458510834527174229636966160218705708816337736647521009994814436017885909635723445392363238809493953652261277221176;
G[310]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723052107496729862771235061177759838348197284202993201177687066269862770303404057392443898514647609247072966191596754797761860573278479714104322581552656585198353456918961734055669536790294831364476699297219477604839034674406160610354342101736789382235711467157564832497110347588636018353568914030902892610508978303922609837201255740407519890454120617359338299114073807393176900651909508396956952930053240836125578907110692621964716837593867075274367679850155064465214370648859287136372591510594936232757263878883987479464820439160426939238982190;
G[311]<=2560'd375526848904934906457512884634274695250024299911217239717113928047055418501081776084835185353619043949816322333265954340274882158468024849814305507487347853454889731265283872679630686449957595819714142588178606765900382148224723052386591841490623611453870657438563174370053109572667002577531568320968048763020180154273845619082618629380564226211690435244469367351423590419871220667266970834424973878696771591127051561432873154439612586525037517096389998399443211256412901619855546465234714211136371514609737617441472398747874418480378650530842482186453700831188746202791929713950839881885451842957248714493351461205783597237054270720578342738441831138165111979791632901827892493633338643745707861532370754612041306198518742905773792238515446056540038405858310385901900037;
G[312]<=2560'd373721433077178983659774043465613524924801110993599615069992963155275820076615329483546461043819793951744042388502183442891350633694048281361477292991525872657926344144579898310437022143955696896366026922127644232094721293202169792692513985247642791411580721287692795094512308871201313573323488973309438302500259468340161921149830438881342548810943427194346022056203402593617091337026873782899874401535266454498896872089472856253004781580114241165678283343465855848321180349819789605583738165087363964568954099029458726360047846220685466188104585336608086870836608229043001209542299938130751477964980172125800743196191202587941107024679940939944254987438836815260380180782490596554903723616496558229528050557135090554528007992172401917454911788853494198591718952745313809;
G[313]<=2560'd346753005094588486669950423090141556831270931236587125728652429030591608673345959649455955031653811663935251721904750449228090575450056127101675945172960055888461685363580268264044506119840750807281081761388897619368419335049043406834130895894610698270269769161090870688973330402985541855085352475722969025000818535565406556830557157813947815233223762735511540954769754839529322040220319524428675555637680120731468334300409183596759161638829938988547381162408712648125240563404603767590468296055412964293827651868763644635916362592247314272124284623804988464507188000981603189993098272695251365251176740311324143203413323031141594687474479246903753817068954182580993522079537960998438902233041918952060217216840687164484318756869319992242902485944219172964622790030748050;
G[314]<=2560'd346640168219941423441086450276847843280448397878446792590461653617842175617255904587188902547472858215744061801939558330603441485461287807182527293142884159101823060870283554753895673607655605912436020269543783367467791647097133529064074407151573117042646606905085883606823380045187555678723680679579562803448935391735558383591429425455394538786520034605072689644732490411160447499794462515893546241794947868384896336299654565257245550149262099655998730497102169042028996278067220784992976891196907369152346282674243526188841944597236624354454773101839516737818781608821115180028728613429214872851613116755024118242612120136731854521316425134439881502123118136101141965505959363960093866815483037022364575421059606167214102626651403350046428313727525681139908817967999956;
G[315]<=2560'd375414010409396346732629519626342080899058358993871893160616322875534162469465899776576919288616632551578269200109209183135056948141567630058938527281332722272110616959072614031629531376579418439800342801610532554186712003497891829880739530037215812692070587435193310602965401489655207720069408626151812429832963720252982811187524887725951204819700581383676497087019500144762939372633856757179644229107349380387455863669597079327446704620035852971639730696996872383804767960251616674345601117013274532810388601517987104021227455416644442113391441927377043010696711132331306483612485648346697046214095045776441930478060724851917772448464521825957788774391874281697877140970461708234507039035198648164999129368798857732216838330100723128739614158334944280592645054188763250;
G[316]<=2560'd346640168219941423441080691702199335269302910639842536700458005944222164396309756752642879434794206514572032290904665845180323790363793555481396649501267759562705865218498394460832823257968686155584401297841388683003465787073992613012089622363407788145735809484120244301817049590691043170228152020713586020510137609497318889746450021609580376500170437274694148590083415418434832647042954451302782390847035313840995138326527338296101133280059138939314224657543842980133709906860953706035846389888629301867728621189912707555307292591012612543318914871487663181346028017748510713070389310075986373683274168877555357749131345149766306035826806573488913671530078288467162631027582014304413236441582544335214610320005908759414676087857644320322607736437930616089235014966969424;
G[317]<=2560'd377332266441024674534038617167303985585244482812850037864277405454706906936976060827567322522515847482713631764029872220365961238084088224477748256803143548580879818416097378953529607283064010941887788800807396761176730376592468896783202412144193467099377816342359056172163281633880165342604877886285656525015890761329995639098286429011090379494943191261367212608517833808467068225120630835995787715088206658001687663449383568434877421950823754890067076949152201831550740773624532261085565698702696307515517523173673209217699121617813531319638863974336542690962268556735197313854218745381328097710055792149791764519373760634586753657851838388820063686927451090223217865362050788865995003530772930773664610003450671668403031470197093454830276622929149971537197466346590212;
G[318]<=2560'd259980126158256635406865026139233666304076468074305095169198049654743741651397094953947118451600235760294816559249018872235399055713113294672479368369742651644303149117602459630681565040709667717971939391900074360034738822999161431055795162220350713652074458878819684623833748285238489363611154500289767983361768241034472035920487485002951817081881273500699599762242663168971685170457385566076741510989426617725016899368838419737386848694780438810272967072510186519730748321056051679406893906168173172514425350925482073336514346282717304278813564940831046970226549979491771743022925071420018668751731900690972091253436052256487803078521681689591422088605159563550733749468618114292415449857487805653059304908669591610504419790829727543105157635554635299165466843037315175;
G[319]<=2560'd315941019301637840741606719666406898370318314340297958116507573339952775406228458391153395459250582762584154730155643843551876890452632677705620977118662112025236493733768952927130702545747925431295125757531736825927544269569722923832946344126950097332490215582399251696040538520156072621762269372954683408479281866713268152949056611772588120870756657675114494324868484989443638092545212584134592762384191607545833056625965677764043913727659442988916030831092427863868166448530053355539351903380250578657581567654106251023967764798756807623009632303725622229073049735134146559764919349722069251469844105835348409142807007062033081026483547050461020415162235295767316665553949098958968815971386788052285097269474618754722636014034361133543245480516268054674380482746205040;
G[320]<=2560'd375526848904936542061070959929113119679899335218837535980752748966041383386215790409472540008891051625765417479546745746262134113710067793539858982358532168704980829821235471074405012705906548985063812969361550487283981037675630105635799696843133416296996319322761206215587210344018573302701787178724609438997401854599639298057041743497564706473801999298083892330924111559500017281958527232364289045660260654608601705172991965011394673953779642340681262933582337612005157132188598045352152523375309955972977164892251612680441859963566581388043185519495145561341647616756609350235336319945335656034597464813086946654171203608950988315914804170082949224322127765708583237474528729053499981908111331253927734227055769684720504653723099881635396722702515815931061596905623683;
G[321]<=2560'd346640168219941423440988578396104423301481539449802853021465094361192219946495457141142565033507453897452850181595683976286092803514052172074760706681739510818511965200061610304617990129984846043256177511350570258251860640880652062806320583015061806607306720560327927678146059150454415416736147314622973561432764072563359422434596608665527785035804915366289212138832653620871501753822318006497490525815686902382491329036509812759014086562595115424139709060711614487732371136761543375240319835370715958140482142817962602704550055219524932831715459181515087731047335403964264810513916701825419226348017738901395820901281440184819306088236508616823137698774709479043196801944794124573324736612683534838654435454115462362681973731199915966058616792880897460701747695179306266;
G[322]<=2560'd346640168219941423440988578396104423301481539449802853021465111213903647704711709828827940022100936906611478783216268957939562764555288225274973611746392107185252721190639162962180130164964029177284216985784244453299952104949753710335492118381791155131842906935767485498729277712287017043249684757671387459276787418233663991592353172852986355538450570825600053759930291585796790995671951207760298035061458210539146948426540072875072240666284227243023702372066282974865932387859311390683192190995295682746561970317698185509103136405238054149203395383794356159946455506593779298837038536864235005996237489822844698148403525154519962307860908577801323565385210282856571033500841691256443744426974331689234215901573845314542391869954925090227334047745962270121620355321807402;
G[323]<=2560'd346640168219941423440988578396104423301481539449802853021465094361191148479959009337098245242486631442874245980576612397687610053193040420820426021028752497047976680783540743429987919403100002450269510362213986522570622108902775284739914934905919306001776762900270396754856194035154215714681515312643378537579207795652746400795811399851342512817109215014537269089309763844835099222047246867890362472484554955183396156267984388925848147149892052950654319418597765604801263742690053140946263709130023340782575987191881207227708671193751401131362201353931822561450797784321050984334944254352718186260151830655212088882281641886466619045571081215145932957328400865815176393177890736305714660492463608645598860148010755101835071559679226997905060604997190238873542298473603841;
G[324]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500282773366044883679600277988783080328995310218200089877372429646475606802734884255207548651553430591519233595158598425864076146643599585119309746315205823590098202634844335782132701435117645960070280869337191146978736679013038041664194722638845128531933714093155286445130949464312190849549750370006781649315134518380793965947533579202329638863454760271761991347379013596704377721705739169415432429181549480307470269024551257567795895257127176809791664667105680773746252001678868849689136261350204269744661048518238451588732412715234575187525484489075654345075088641109380825634974002069363988789370869215449753253962345886625085726859536091978316005378868928749445514547;
G[325]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979699112508105382867755088050408990184665037417058460440429474492645488999355748919373060381364373316207943159628206614875076560219440309328276727581979869315180385012819741960925185380895340998914104908715704066102999420046604102879142903973591471352937643612950837751330118585455803687330260388047502089502333821476021364995091780388390353205108444819474592136580346234316958360226332279537218233389572212849977683880431582668036393847077671527441663071028162850164524743034383787426415422533576529409945787139819878214874927741002318767662539548429936768742511936881189660909367968127042367948732845290833427699208751572;
G[326]<=2560'd346640168219941423464477829862029498531691690635577009575698627722631792078647363085263079588409114283765262656054865106275795697842053424395408592189042852404481499917277659289075291717724433915799482678770567422184585568855856127823342343638569452218319752471314986026872751617862088843989562149607280589473722184439295330673221902545745124288394044657617511390346868302409914202413576426586838521510737033794353587470586750853072309984164636651029780956423522043063441765605738771074190646412091908546914536079492059956911902863128050285549465669791208761106846875308403704081093745889880616758716404124086604056411172557302419612230713837096345701461943183340478997726570489337289654095030992426572284870869923008089185175908786875225097037763551422769848701459437750;
G[327]<=2560'd375527287958923489225323248330674559346377387611524711638634604634970123077971587919760833476594695461281705758322779919142833332497402043435836023313169488676931035304276958499035353136160949225262753783569358694867345594133357169585681147863189005366124658613748796736257334697624939339596796649348938341023444674343861611212738746939938521524281693838987960777965479358136732021709250893317888276891150828999133989812944621455910053175507442808374763945233285864286781541769572062290049813973322048383737088556945086693053414396550589844032774025018940179950313956040778532601560017290843277244567726323892030301161205440208570064766907258361091524555390409480736955459067620957278982098700374786965757084666300050083213769343149201406035544775802957907459189518675302;
G[328]<=2560'd259980127994347679860592485004220513219339050643260884804360016519412004006960913784636810804791333507154208628635783266028628230259512502548326673147421380346776586409466930890958266309055334770110689138141094551116272496008570328131224747198448100145273616212045843588824344111250022290669430793377486856382256077828058980814187376303906820812508929410868783068750313204141300628675900014067973590604335650104205944852447403275059449687049271533580576308902639136609313503016296206977045044377208168602945391892247727041543536006343464687564481371576464296663203331754841609028535947021772865322338501495269859062737198975743404004975069961362994070416931450407046849650149910794442488483980900135756421899848170481779541525606293929581439329064194327532021724875896691;
G[329]<=2560'd317746435129395399141435557912922915528349966869745531896178056794216570062245169126153431282803090798434426217887605962511144850857554686827662706009533631911208691926827595304492300910046310621501763052736004665215142337868771377624286612753621676901750661214658646746348787633501367745053540288240285474834442447244215202891349938541259508420806375538855910476970051852703559444908954335596460874223204840103450077239624768693707703279766491187991001794740515411593395042468017446407427594961356688171139363430336202476313489791148366924625336391017611217089251856034387546278705264224233110016029687781792841108327076396239232007202271307071319166538794928538364779084087819789011835476037302033296320809187152291003986808305386162929496211804808485326719305517504370;
G[330]<=2560'd319565957490035109871043584065289681934422485167754676826192542481141305833073855039119864435517249614909361964957356725230637500220812425243906643748540363248596504549960062295154822148483878375515465197934897164523129299435085806695285824135897744869823614970527102557583381715977474112309982627812871863902671434822140780666881572988361676477604660099866912088149750953260486228403953113472636263104319770344395240118525199447374295416434649970553400602873166156972034892273898455002956337732608121199602242429411192313774929809305041882702707014700975340884369490720620420811820626699246897694871907768577198259692984960681568193678179293363637852770364915126287239578552204181811689055074568575486229754126097125859199648683434543495531928491545054205979102411457644;
G[331]<=2560'd231213364138034241015058140100484796374131443742472390217035448534456112496072872961159101447784732140566130633039000340623129719026467055094909058685300602162580624333429619348088780409114397522121000354162311441543048340410660709353776568341463975184591528256201143628690909740014700215389292906028908381586428988753962142259298575654802147287825902078797325541455018305971637941268796321896883631502902332321099229777748606965616960690107610916752723230309229655365202539957053062562144755282860104858285033150853909753312977112444912824622768554708899815906229838832918693201300622951775096312280389037862964190304828712673578469007868709246648042232997980183832071217928629470577350464011996602124940243639537434205679700022606600704690999654489302287007365738575000;
G[332]<=2560'd231093473142809652519523677038597848083139368407209418500205612149754757593385154884838765098567465601367013585000046926510336050548163009564920088799203859748031568393108301337531858587748579102693570737369118835432776166505922427928305051347262924033457960198119599039518308609990930412394612691091576231986260927679999855846865383453187396553880193995450892432294219832448305393237558783263671327427086377645366377043617945443613054767241130569603458701598129417223773753704867671036878165324638910136549230712668261863550364536477569531371620412183365081675871777889484211956816010164681873300630640832138709036218642257068236813553448360136253577671019240342725545158786001626328187925609875371780660085572374100823202433298799665044453215967328997557736583626582905;
G[333]<=2560'd202206764902605022391067431222359007799262993461919324246545821611059319041744603128948280439808329973809388558080870997266049294346752451668654419565604041973836748139969024045288101576186658685711930412627214143013602014883711051258196630987556747887041772363014320602269990752844265711942885097616989459559037907216752911218529127769768030762764973470811481417557002933306134943535577300215441487167107163375951461564429106117986126982827900669129128738474908651166346858160589748121681885528295329666589650836837959839079841688652123091766647579108608939408818970409683038218867100721355927561076168176395755954856741609727424984269247810964453829154269231699357460284420769909132702075946685603426628212894998844262990535486647478359866939861876665349350082537105340;
G[334]<=2560'd202213817106356880064049139230372479690335771558318542245979225956319614209301758826160575330499100989788001235206929953773713185979867328160907803062047096912555999828486132878241292260985017789540409063100926103036660140401929245755641400370242440156125091551092802482519812065794806622881987385726258769526767018004320428917197279353854546287156599475063367880889231595918700997352512958287019139814420858686155498856152081383174147070766788115435372317309141903173546121567334626142957994969532487551884659067482816924930654004745263859782243555190332796561929349080778783238893397146143314116920703311053636612218354230889153529613976715696284005308125815301328216916124976192484539388891409682900885773291587514537345382233429252782786896508350603510545315804239271;
G[335]<=2560'd229288029658953732121682396643270210793679112876287959704719155356122284956587881513729214842816093146060917911438725994345069828034162031524460514438613762093228769251188881007610297185265257026896510996058254430297747611862890818494921260346239901106517374359741597707580276940232581409497188374812564053979104936738307736478233730970897493002322161549597770602096764598844740598625169086293686868232437090739647076900315416592421550399588267513878105497514951115515643216205099396223574154246994860798002262083824437407881455439055700149413245778574405226799440899456448989445048999485773242607955597837203044090222902113197872457644521436584340057185107379282292052373502523249860967423218123654846296622914977522456592416072596594318858743698162966153778706137303144;
G[336]<=2560'd203899369568477836766056595285055287061327936298050469777005617163204429617265137685121957730154756481668046413655476154227019157956216510248901014202679442121094540461818008755469158372462371094647283228048329083850024088880832238517561473316735167430411415727063286314128875737258383907551739696970301292879479324146904560595117745576474463908532994172526150437337251949866497972035906395605524898297812633730740453029526071019667662972978742793962025494066532782640187258299866833652885659308927076377945145480086841204990552454186260537028579376925642756581613062112965934542410670585875781150217353899711626913573717640963317877331203208877125700649318839828226557496137779156504247172174141759891444585719261922918600461309615052982494283103178983105965029086231201;
G[337]<=2560'd203899369568057377612861736895361760200859565282768434459588093221777683577267322315156621727125531170812870950486435560203050371179492722570982094832734265230081786938662713465652299557145522651898841177148077920696824713021489813912917425931082723285192833869280756578218704131868702755522857523142473294832868550546609572016395388354486051730494008750943930411950109959841573747886553609017318439774010906545937247293468072096539391611037107748013891857205839174558770539019612426228644062088427900191140131803013438970268525196059383947144158095268961260413353084274914322412254922885605143194749489978894743910853124712149882411112057044843877859905015821406339590494221164409449117040268065651729783511014866140305870615464949472367983187418510731026189425587180723;
G[338]<=2560'd175125501659508611091062783262764904567696519346202955976703954639031329085300366075741684755028344324125037084524439586776232704703765563793292582900517949139998618455789554993667354767436315485701378219896216230217526702842088462493805512682141646962436606619661190350046719622612598862943390910583860466985736717409047146281431233132844954978107097806695217957070198210087871057877377339284162854756000449107672893588686333725480911881927918744075394426313590315549977825794625488839900842250096049245189330113229763776881821822281182101575798716068155717652170341101887371928987027418358999886298642843789964955975562146524614365262326380578305104358893422912181607594418526357499187021836527279051709903080668699143576681263844838302926845510544057666374793623946331;
G[339]<=2560'd203899782795365482519411348736625561287471747760822015351949233954961550190387666658020230881197431834214667160287708251087276913909470734582862567757097604784719543222349049627346167112966524711378405315092616226042851684229190888818322531072280441926811881185853561400595592162855024136922278015646856165868074603087228527152938915247660410170112077434288841454093930923132579037332989317458425282698267119550933018732063224740366038932361771771361968432578836257523839830832128733853138767959936296589930552722552972291772591727728028612237504290134855351187270833623082612086341638144956569910350148883189391068982386263652624292195646816988748809272316637491130542047396803428677590281684453658948922854638921585644540217740292912715417139994886984226146349171033738;
G[340]<=2560'd175125062699681526300176513193175894891206165179899961613962716975545489034451908493261700491911628073648422748552856978655300583055143460590561633470758090458660263230849982534328759731442706885747021266315313311058862109341055430542593198679403116740151059520580630265948656736744968803231598565496574947447562669887884585280786894911623205497951507598621758249801484070485100457876508104363290869884216541797734088810922015720382058129322267463624371607130782553573604373725902688919647187721228847932648274981204418734509288567289926468978234817707863260748761476875847948132017618757752927166878677919506869574900558758822803190907650773224220112040471449427116501956434478701714633148487111941195127818865094332549785421061668717187410377960553615236212326975196439;
G[341]<=2560'd258062309079705057649129236559732929448858679835146770035648688992295325477182511194167091373109335367841203169153887884814740480771036109857506036165267378572634910339449846160554183414870101210686517197184239566157106901876084758014144859286205069037808504029675161960175975751512619869087658555052853481449886490933777550530202705311964238901317886939371800564314678406829611409488492697787924095655845328139475129957880297079970392651069758054962498820937479007648174776453122727750368734827519178908029955805306174504944062827669752213758127887363397481084757615506471946076546714427570891052746996251629829705958822821582190217360877679681453910544670816775076886065876762684259734111865720774352489777683301663703320189551404710869967230824658368870453298584197973;
G[342]<=2560'd177149074138633769353906881315947183979968395198623594946467349968799734255548500348790490968646930242862562811738295079761892641107257541767918544808954686351654154825194381375097541703955024697281519714091398650343551576210096634256780359215271243638544957257694487454956545109407072922795844466166781802073561908572952654578917871121375532900856402445098693616999251242434865950730890589578108568232428494093550384536019430771665222619166394374144790282657210528796672175274854368597724581648343673467709435192763021101015419607574492190764033034298234912336929670593815336706325899426463467519663526306659785377957687562325503891848571552275978274296366648668057335709841838529069075545666960354865770132624894232118614374957207054516087073703576400268283687054138979;
G[343]<=2560'd143274299016237833007690268197125428216797836150202233068653579675122025926587856618466493173159944219948666549879275945824836397778556224792857195600963423208684606341540350403281135100811945852765427374944440053632168955128370836609715702941158087155700676469731785188797950648638846046203662951370708752419496023667614578953341698768340345352062098471234766592933110990797401674671617774317423703364810800314375588129162958418073054937321771198795522769925049507555261959807760357622589451327766571198497109324372779069808075523966126216507344955840558983281005614013388467384427661703635612943247172742820653404513420135285302860447411713430712116780396598821674356507078974985212432260653704920654845485446951062085410735959100933898422144670865041840447336524438;
G[344]<=2560'd120201790053917272393622337381051760023410450845603600730654865553527868615055119926463724584758926560842775541495884199624683322889726253740389581569158835912961651449538450834428413262766944568670934987164711833745391815234276218528163205326849351348504820660059599436896496677007545677999018122660029559528561171115816791909644170420727052525577112404594939841140326918798099045108315942862559448080773755211092644160829695886629653093544214663676456686333146258540506041222924947429181212892621946609413358414236746521254266892696742986312232851649765325945433206115014058704422226648162369513442928502617211873266133570539744328912093734558940047138086909728556910941924324155391550264482201621538280242361051881023793540993756516150293297318699104065812001653;
G[345]<=2560'd7613497445223497781101466999057813747485980472406612769620292038473717438857983851964823216654939849034781152639057338441474446696420814417884977344693411405337799640288820660018951849486613474584561079206897797589700573349167294967223233732251184462196649943630427411953941268109214444514364332369719321683432636900582391245905793175708035048834850462940487468867184534007041553277755499693779889221113770698295367024348532364592800798041995460341355812742155116749213137441839772668747911836461109702839181286037178863147912664791668099403152270308862265603865520196697179843787575216647375251109921743378795810526715909893377905654054289697377798802892920384467401535174800160340147915050991040072316922649097893045957672178385847458660471003347858543728623897;
G[346]<=2560'd27081269040625732417464653287115421125953690598544427549292347881595370241624010954936334198933735583434565431742723273016187364091205029932879456818244044057068327877029397113527886685753853923398174873253328414750521917045592896310354932899830624278916874450616248198211112669718903952390670303407874076176353138200395727592392615879735722520424369069000977754096996472741616403615259298848904196124107782778789332273382688723490223673804333708081301675682221833346626751439826000759090660141512916616066326170143461687222227481119852853317918261366185216075484988260041860259468959478537795190400004398001115373299279836084683536513870384836964812330381468739915955843104365757568248761425916603233737798198128106584529913866380594108865489795037518543984493515311012;
G[347]<=2560'd112405434157560890358499200341965259584002578630221989362209600832654810079998887274370094391143277033420270463083097943596250754370119088699975183667417934280098664639086962350506633127422903861513531301419591085212698060581961201547278189605107794887339406970056654882713071899112427238201591719183115718905710264590431254528880318688470586668296183073605268047646820895609921282090550188666916266319130708410650502844697981446523911454444044175861954651309589356115892230753477405381776012568826570218509206522924658099801070432480047600003484376135277455356923383071636780506590374196910372164551747523426761876394704015122037892763446670743309846984129174031775959128023041153321813823892827539734675157741830300343289911552231723062086499038606017186957906545780;
G[348]<=2560'd1692584945741080180168639769507371137931388075081459600562560036027464137542465951709212441783832476976452891024543055661413835933783783520463065306862150747185748140199007552492613965440394164749546128799331221188278566034403950045414144680033652854553882558651633061245924852675154344096132661539665919076139441102480202832458516969235939283036497559300397325516470657223013017014798581676744675706180269720860930631773726859372507798941943594089371877539394026171782253312885876297823208381437555581666094716259621231527880095893690106297441952863114583962394476210499818373652503520732267807294166831872843999529729142312214839826405553647953641005614695730039608527824482525979054792282093348618306124306013640671082864294178193287527273506838625832435598544143226;
G[349]<=2560'd1692589788222017297576501823972598245871106886254788143216516394323782424094606953498749069192448427543505223121410157754810543037530461598141885770874968303657695295881081277349962684836879462662009347873950465589675647837912331472395730196558317154460852193154102104104705493770843532323665913086329441318744463016110015341011951673431897801546027970251518957452075938744455742416319954619399034231254999463935748656911299580421803207736572905050705221486384352315608830502791341276706036785666791995794246859329740606687225228313506712293574731353782984952475230677615562395659049658122883899080521401632998489386796763508371869563681954029811296234739606762361498558474650620814700189097135664467050434124913824070193963360732604902242901124501937928658067709395019;
G[350]<=2560'd2701258132438165946309670587038957502927495619238018910458773837813198137029635075074521890120764520891980739699612466378086581767556224116323269489490485874847910992605688940676767514727803946701742632568324932340261423809962499620051569180010550545138894801707399655602754238097078339960043321882283786584051075275435239551990369726687205275350371714601511424006387656896768855307734255700454040145592668147656694261376584992924544412286404827233336933419878024568253782783239910456193093177462752584902887163727918189377529656583661802145695460749105294070459439874815366182060547781708860029122926636650147058570911048654602388552314951652526765605884491486600637530406591960930913519653571607582672699318042337358864584435733580206143106599181558389758987776792;
G[351]<=2560'd12305564096907383965118454744745174241888746486041722538907866859772013926850738682398951830824294517329787788621264525507362418291483017471118379052291371009177380959824187825489366226326320796019203589230800926371681666800204962015793358513487814681253109336421843384134275440079506963730342598417586798390009030759639916119522867586975901460254017039876482220392793420760953921774508306204673811753075558722974700535562824751894285192315251625420372111851746007679123380672090248466422370221784098848981008679444776542323701059083043960282312550686785461539826381120748934765165721470546295139267718808515690116202268845105842601481473139901083312414378393064946347912600009724137736213718567006708225613017517556438602785109921428017359686577773019039567825969547;
G[352]<=2560'd3137184666812866482646569288086007109229579844593183884807664840349731007910793662576251725821761916990163466239305788150407564691365809219975892797043087405118356353718410857335600548286808838955686482778588246225835990622444497676163427953656089959559440724366959563390566241536384848493233304500703557166713426375583539470524998265560073510606419969279316824025602089547421120438832993031079001995891764488953366821292995068406228897764269895590411965722626127697269200729546787023497541995177775992003008942663087260014488839886005287413268713185072422240446893673070641353501063298077634010002660161905738337764260007897734017594604577587483539206164885942036428826275801698303915573031530295651371887655324460060967762438697583150264392781780143594822009308517;
G[353]<=2560'd3550311063078637993014447135988708937736428788978431972435408056776556281780562112183194344223706610489558629884629433507165033298303721955531596908043080383444879721292908878985503227961104353533320550312760803449991714041732177611084251507253388716081516294291549411510276700561902193741142898032145416962885768826076969233059215122439316943046726706661242302375625418968453070926760610674514233845591724360398064749671294887679712059596771117927663427251087292198336494596505907851344699907337114538586931516236633030391534867951016659181393180488061798433661893608350408782519790960348786082776952368083776647153641899915610910024631329811064076498651311305738290687366161847220883526022590317271830558573719279229990094596072939075232513621247886043249190974241;
G[354]<=2560'd3550311063078637993014447136072159522392602710432389950934599981186744173099271598362305211224496777713328191523732246509896775714719536969459759160306927677032986222123380129993012003130831161457203330312127740118501175133554992772007084866389991700231372243472776883500168001368838377291105890630406608033380658896997324222911796454142815115783821962522721882484606122098416193226053909976662454951128279427809712867188211357278189983114912115062159737941007424939723871970744878557405832080260412472365051430932292159419225701517618786712245004368492447093937651878956721789146357071224019500614896080126479019521152299230382181123618203960883559435485997771356755434289103254716873143427055307629929232712748788546361032222350445788259951053670141312945291030582;
G[355]<=2560'd3550311063078637993014447135988708937404825957345433452989312123858201021739227759742648469604645754147182459071368197275614832284563857763029099390395387018749419982418934320441202880814060550782080480533115876496845155411111383827295429415537275005271354011097421106307297675037651714593437422949252515465063766303258201740353384162009224402123692698357351873398265361809979364909473933103926205485909755509695387987718328088019704029579022769633949074485353409027999708231160152841682178970216217625198305587532911756359262760728397457543762586359973935670104743057946250428748952885078529958905452312128919753520301309794698514945693266135973558056181417440920272947375992085372756971139283596653792930428772592719498749742509962371154780998352030042267440928070;
G[356]<=2560'd3522870188894440227246422038399077487991688511324486384609522584568205025544895202205796609207873468725147419923017261708828699326661912471573649605096160597008166563460602052010205453719981096283456631879193509896212287336060052734009944774782499482433090609053158176449716280915070627621079482644645283537105324175973589073464090333780182144197410923377621388665333855939015877230785250113006278918700250824595651579533964045225222283078496829158189775666847648235471494120371381750618526402511723988379365262860087902485632721280447852646481758599842936436459787790633033133751661266445225629221483528563025668874070040855457275172939561924347038296322545767362973749332926199604802717509934651843587628207517041402146956246872347274863767226907683009912052389920;
G[357]<=2560'd3548696894008979300910445659659907087439347284050083621140114254381180679557545443296293226957260287489502840055844856415794935349408624214725856591213527066560112241826081028663065228752617347994779355386557503460726597010443954065101028830312997798151757188856218721503127251280291051798983245568783292602378626959404746486530432835085992412234742894258332363654237366290575919139607100266916379334041063542471533129780301756829123768954211409722137451508737034454009526819835408626983051980131503500086867809124433371120173419722043848462349281128611089526574433546457614040792225951083906789991335300021772411393931983331140365673154802843745177260327277283864093964213064216665719717320220960492277906667727189031555238998584400424494511966508007336537371984912;
G[358]<=2560'd10573560685163607337524870642605558137202533465412531957461118371702609577667444234275259288954141196803580509521417584578863637617557989557243157182562308611225705478326942943194848099314922826459307534059264484104959815336108400852699461539814732165932599077414089859626843526321126567180247484126788550904822924133721987613776011961672948334653963256156094394231227946858335165783149413304257354116235643020508268571919644030497472605574702293953841450362275470339498814846936562045020038232432550735427606966497705737855191543002967094422278289297423864310791113589685271384650435189622851540749018934589107250866649479439565396951437030841097964667222727441979255130520481110030053292855047898483416003021531329564360570841935419840314418493444106035518178983939;
G[359]<=2560'd3548696894002588756433497418880088038182367602582547460146395524231554770187800651632611413670330814170079905587996436024052677029998169995346728936573613656058267117786719679767236619354255698955474554756145729858085179547871122260605945516341082283960282759597932799747128435235071258027789034853359351043619875949293421549546313018948110625338876881956882395938014298105718673167893975224869385314146112522378179095763831789789715989077402605203893261545761367970900603017627593496485926275232421386312425918097361362817272713665860929829100437631697479123676114679945721137299220247531689784664401570893961978072991478058970012084603625586577969771852615173588883738176998971583250957725897268717408728237341688658028630117789706284622691541145348331268804247825;
G[360]<=2560'd3524484357977680397644003635615023943254120525215776711246447596300232328984564660091373151175933622165939569685771267841123534466550308144051771369911864601441674273130822666380833139170268628583142876623256703123303602094795703442450357166000344844227942037318474769233632329497557190341447969900886857633612026631717215026046423606921692297988251133937922054075930255529477698260516652105821035092363720871174881011049518940747598330127818461546070008707087335265234271832197771167655618918175190027067328492382992736970820339097205462766290653318570110910128751077312833505029031509396814460970692148188730371022571703576672880367642535585508729742418380280618749441356256428640409729825025509384575890411113640099320045794622173685943647863592891939400305348880;
G[361]<=2560'd4376859868590985324370685126902846184393011801907854622851068234864274879369362524481722797099566176540787253315426473000774618212299299952580281920747444662866161398605750620060866508016605704165647709202290712939766647018376706140353579478645702998164096369772992410035401904301961015838651617401380108438855215797951901605069342207370009995097217219836506283803279400806235392955569491403451530786826242528762187223044179245215709543936640795571250539318124451497593515474195766640490261916130516048767891029171602211435994244469398907135636361641795538832536933501217957141070057207039398988840058806676791839078822219492522789415399134525556630378338553695721491134011036099726123392646700355907401324000124435296153591053428104872930398347680130887695948849410;
G[362]<=2560'd27098809920412622913081527958890090270555593111636312499943103938055012136140259060448948384484900222148308879169244290092453286096193162113754022573233976040476130907337770356012398952243521160984312598178736392269348262734417794044288130205655063015808174790814538072742248724852498359840056806599966035481665838117912646067178650730063709920772406393648331329494667312192550187884492443858755736236952414555321086300399111689680688961122599483290901856327906610012824312077803457122853977461069114122273465368074207044579315738440901350321836416316071055979182080810905902963916926833287611559817006922033640116430619846311085449697676747208294157763900465028206024430804151281829617829242487974111686135245220683789922036912190142045474380373088394325565038182535169;
G[363]<=2560'd10576714357474915621324981377013977593336247741313076091434256614000551182353773535984846664931985636513986251677962104004875621548143434962562512807447099941237167671161660660188324210105096062495159763677944166319122232394258504692089556421582639182829753395783048385017478850953127261554153979582928176210109318355370472055201619578335030111984407593240021155667506965284846016899493371581677060805533565997961360610445010865612728008400111539605698118406878044829690594434851320171205627393965647491876085647880532644970233497277122519536680888658941775377301890447169548770105208431399177112311449730496402868900983990409437439374960532975193695690069941342839414886332074040837279419923343912486380618978524612504189773996106478144568532652960710190666331726080;
G[364]<=2560'd27092200411310148886147691466406486094798151457873300244785359417196373449680162702791701962835432321825688238902761297356736237540715895370502880446112789231690085879699945692540629523356485412261287728868468542478323432831642064088983787657498866867647033813520848851197102047961519415086635296186608753241612085830578931320224419614710287161892260822935391127206151745925996505649074163514478842105887054307053587033992491924724124413818847180454864249159357702898956668282322860775008481494365554309777331809767810275705732455318379185986852920974432054906252015743874192142465829783018501578026356651337045654571391220924764938900140037730332602816515761717578998615353569956894498309389257640687963455535967772927562030596052829684063563636760661275095923439972864;
G[365]<=2560'd16779892794043018800058536356847281845635341092123483811357697625583236672588164988191702785858521593240950989620340530087401582779048464397597063941165922330702537479712557871475953626950496216088468698772395550311623382764603947464416697111529718140712482342704821369724959270108171352077903065345846665867955334816266549163209984072547323521951217563698183358774423672472515107983833247126254279609049437433805819029731945132925695923860646552482352058287673773732068587305844890441193185907469360457527425215732405824872785105270411475834235564209340103039655734644507197942315627482438615737659518526611418404906159088766065281117101953842407559116685350808139349389690657642848484060823618775053898011682593287537638537164932104533029440297618664210049639916049;
G[366]<=2560'd1711852125079697282962856169020494542296527249420747694139009962828797297051382313486418101207001788196081425421589986094090261898597598298590352818155031244124813377836212182414857846276267671392576782871888213304977070184873190293046280664236218294752766989114681959418295158759007827977175576935030287270897308645487847230601710474187355485648881209820904533399971809475604394364554802358561053168675452044547607096257753611155007834299748699007652119289034216734283051553179591026878525036877980056290689138916340266430037701249858908669130256897338341862613064227716827102628855265736499872111653272575153174061054716983578994290262001777451277144648277564029320376124082940716399293662427787626604080109682648960357084223763454906423410647524368153701393934385441;
G[367]<=2560'd27110602279193046132221003166316809846262049193035654484283437390771407327040492952428298289840846404031684971656287893222966546366782906652716452058675608604616365884830494836378482529284858973159503827199361679427520269693867955027705287286015904979379880439471640235951745342978410348068110094588517294979858777525520824882903502562416151641145718550084247704289257838305705514553047819812006229178349312730174153200234667193461457597297990900430424643711105870421575787898555077129892910639888937036450427272205809980355676180037834084094680200827616289001675560949621972999015043602807159917472081843303974482358353162207591117475403955609059524423481667565596796133034480859748453484069575632402127524039966483648231360054710672879899657567172783914040499010273281;
G[368]<=2560'd94207886959121087535283553749586685319992172369941124020543116429115270087301361538459151191350620341596683314066329195680081074996787816816010562539196764494074026824389877695815908738722955718603228533886114211152854004439475242823397884604942769326043014986863122080110915653142657188904719863861611797898015426244210709516698727739806060168160594896413094473781793050105669163012921740262232924194156265652000457084878126445932843820134214408307513969669462320315100216519348814517031820020691290655731171366728034999347312400662900904986995957057980859991221543736471524167777691094504141531948724647577584644922710413951300001216587697136336209444912306170845521757988138968064185679604481892403286789583947204399049678403821121793;
G[369]<=2560'd5563451585595209175416538786692741015271238086729517588251877848071005255856161728748250345327796585628852389833662419682196769920416057867950624600803806184124481572319898520017260410073324961332437833144624621519081653793046553245631111811965019068609262133188440363948555808437457254971008607247624609212763456976230826641348067364798656001180115574629431403547708544658413750841052265634879237396970313047782845398201229590390515402662836321648401168444431576135760127261128509267375608250413083800195468495647036278015287413197617717836514179322643633568721065110958424754066815603675334841188337343188087175474088812626341614349725610985772655494689606070488934000884830341064919025937925387457649883728104952814434479493328417280;
G[370]<=2560'd1363549467393606278976008390815821103062068714058435599896488595889099501929753530770173431829562062706088175333682611897974244517513745338691196088264229149630987751957195085415665628832146467942700244644309988442750121121727727606553585463057024931961400749043110158212240610851094686455448343901851349091623361304045726555221936735636488986881044717512735388047391366483613781389322557929178801287297518948244875463493442203002624838023986332881543213841412300563103026311453438148492470588205223455862779553177670122405229445743128442565190391152266085084964384403177767000414575330856496167173162797781450457449852959933437209095024269218791075790522600219495486276955054119474633422526956979291351854017835295916494501894422784;
G[371]<=2560'd354903159918391446548098474093260125879838002824918672182813326543381924411288554847244226331211156275022321376137195624801437177392399008634648996899359966851329533429307105270284305916876873461113808654637253438933836765091684830408029862085958887809653124066466888540327120713798616575427554345775004075732044215196500342464912148174213945564865274466057715447646619259820124325849683067707589830816042421301942212784432227141416709549150464614438017751159812137011260561346220194047570877942670358239323504345202448541749797905772871598434655152948108834167560119466401392705886670907694274580838972779250493667512003855405024885018762649638219097278684664207225458763696783021794678538676529405271401653371913048438861734400;
G[372]<=2560'd2671564079244667609839417593197605206056135824187364182171406412902281836209443902496280711049957116598049022436932769006278204526236450097461426406178043411541084988581199708546454282297003685103268613357200669861128708124283608735776590569136179552904310701247921259321711241003094959725828291284100533823841702844368930682434827712455058946684978674745725499987877241605788435318339542575125573852270045603772100903263580969470593377504914495458497692072537056011459490740646818530293947933431108370073828090645521003549350116490091550208176365126445565979069755477180763774686718106454527759879171189163362095922652397531030175664553676538633799616882334485095989303038712621643506550417004319964872151627319118281962430737;
G[373]<=2560'd15811968010149373620696857058364560157395978975143193923379071207405439786211493537620895136724089603888334335972571369856062770780123405296581693326015012909969056777373971108676456188435345659721872592128122283953444388416365047349738532603214107532907249823857903184812714926382382816505564641232252532309324161530832303575989262011685085203314959415810682116841938876170532487358236853380772471441843308129841633205079126658043242523300454524575140776280035027847282926866753135379998995551441644276508067620432844101604642059903167350618977440906249562370078191404898604717285155986469981243288338616151906263136930483378163312301845787953658421809727223782587817807874847506981336193198317437753154053959980284937044001;
G[374]<=2560'd40842962419026583398267838919353303601451783888452366785209754860268773926641134330802021273555987269511660904093199555301352784077107657886671062296994262406056540947923359090974155609806388296902005643770944556245761223659808829133256044915606718049952438733533382146047604544415283650112386114431853234478778709458869093056605532798675213912953386962250840789667722889683493178548482474988463861670939819741900956054137109758774415371659781697787729692645255129333699538676060415496308045652887151957351883030547097283136374320006269023441797180782189709973277896558525610498292957452159641408958804254842429469901699961042251330473166867879635055675608254925454675552535689176657146828036647573934250796236615358362112;
G[375]<=2560'd82353202080926885845223337108165536555809296830591425626229192259091583325297743564420679470064883821240187598063106207441214316582271454872924369390769593810591020509355680085098843741966203332929498795068276874029309240669404631014072204682458135481538246574334677814261490172853427570261503113808940237395262759834123668948101652750510337972706826590501512681653556132496696844672072331981331908618073315149197780672114176052661371508277758017934891329652121668245213802055657176622975695985426784487546214348686524979681019954654757666238634009068133468339850405762800211430185934420469832039146958894781476265337691161335877405168203455612272347580377179552594952221539822992828995560096221303436172334014119564548;
G[376]<=2560'd4826781358949936194836026256926746496512253851588476544305925792164486316928721729005994448691950478722191114030035682369702576438773121323206389537163573893395015201642128053741957307091443137985463201650364503218282274030063127664305439837420368240068346985867789009626842859905915168660620652187564294688064973698685414092014276019172288094939062862256521428407034073231784142912034444697528726997198372972954726391258167363786788901906981185909954570433047057345516468440205998489835063746308689712070890567023830537520574597375354659395734882518872660950448013812119667577682579173799529753147525426210953834248381334315868798487661898893252195078710727504601981455238468452618013483854240103767355221576737899027;
G[377]<=2560'd87148741318084025124055811997096458145160558997076420112497220783855209730030143015244131987176440242786232940037080621032926921358047821726582214153591752748568200540307976019625341009074546911905089046957771266895631115442600863725426841910862069608262918873581028392221743505031956218533255304758802446281733994742422072048685367061586631060822378535669552596881305370080625697761017076007997127827342249983889066097378324159344540387757665323768970338174238224809500527636028862379605765510527971100432706340311888766250532160967053898861434650464017050503161689273990516346151833987286280275316859413997189801922581174567872891419222071681471119809987821921426549883719762666289087644571183635660840937533697;
G[378]<=2560'd18118912087321698212399061878847457579665563100085248362949864473457717304716929089247228164545746223665140136209880050906215991351561505525898948189465859460274126483485924118270924785686208126899157877983839420685414668115597800381114615765381926869088988924959267219759554809794512064442567292247172875563088390403240605801396696912405316124638081769598675038328459068772858208315472177039928990044890431585141424495877063378083364627291915983016897781643443977208463668087990779081401367915309582782497627797726132016922619204764252132133067240581964155748892791351766694410096694994151057874007912453993870311015930050966711979066052280268968473364427014108489762751382706439836792245939030141421466065833984;
G[379]<=2560'd18776132729502845738900953295118508527321617869445447832685640369894452072264650389360019236661667124568518698628886498511430505279394553645416782912704654223933633933528488718361210088644740752282610530395057328118452602242332084326692320096750881885780679935478768550661490824694675157256264038526184090439629342743322933007160654872453504645632678378920048433643530300330480194513953602493336335460459852899231727836413637281807888645671655316083174109125627867760636070921835502931756198261565850037902028648226219420864575449698772780484173829970872421931255245843829099900448389388471712332721316918450436040903407827956610385535639633756843368111632619788997703756913014909562761034561569484686225663092326416;
G[380]<=2560'd19170232477226286970019011297562083084679009847007189129621457815850685097218619922960723222902942963283897963069250433231430100189796467271778930293767049125312173747561259722059792265674871159864029039048540738011356171594293507294465633638024024618009131252248553119174351788449526192767523779300524973112563816689436177134692959825905502815122805081793295589431329772536032966033538676006355375021017736811759399745925912295306141237500868463300712925559089461360162093883676382134882362957891728347823685459437442023839895012654948707328927644020050823337399776510433037051057790247160840503177442405358569497091703551191946261258149936182400253361911162706472834308648663582773360403592795282296632508432;
G[381]<=2560'd4314294691240418387816531526335713783616456948575505491860244906147635242884235747671870111960302767666933568401845239970966371898260638334310012871953637808313820487400088377205017788145800442189562188475895338666092619843532862013699752367362049861267087542039314118118272832601451902266677613787159015889714839395355089167378971264935317763728115191493742249609925793355180281497020254865172965233529740612175703205048327035639283853646500550810549639880729602308670723987672552569589848212847045944895006382407572869831024195938445120525907070129953954868975205794254799160457869104256303084542802703883389101903455547181673847927182971955272651554153259331252519952335301527092375430471380420423377803542544;
G[382]<=2560'd3214660180265199669999223687560067855603769167660064781131483644717957419763782827263551814254821731197135807725540399068195382383235653391166771609396822856093602345340817810212246296991923113715864363243846633833274566601574219835653711331422368062862513222726252407066072509231118002222919570933860272013554151262511434757249061996313495134210203268079775692976180762157419796454252139955693677859190545764499010793499203270322902477052105313109228011436220423055202884722389739190916475374129161480462925525186553013259810597068242366403505295548164677906784315693055013496806465315757349029352916328947080204655013278437716428761030807463142414109851106191307075927285704838571967053363151351320576;
G[383]<=2560'd4724878830212479338176406827669293450660401657838242488917722710388292020502288625385418137778623826528780637279263124575461386409337301873586176739636873426986653017247055896226576509594343576793177271118457212209978092115729009341085479490644226234657915175257783641309214447386976518615623852545145329700774049154392696121869499345490622531939279129511160381140022893650798354679278180885867857073316570684580391301138892920833332614485629571869016795839754586158390306588513231850482963960785990023567433721703469594853017926801663696102715014329724478672641230707560750568171558809641087722117793032359621802877699376601826643945849903625493292877551920468657721607670128000689925648719017934848;
G[384]<=2560'd67244596584852928864970805954253963277735896813354258169653861598808835605608722804558397020020597024322678630195093516171675580767150088853580992794213405156111218708831810873518411429510154441370643509461588253558920738319510191868626129332416161574319127264405628263355461347257305217188669431221117547056385183006152194346122935635015380386486637182855657644020560564995201864972381850718596184788820378530277527037841891806717616604612404738043193735274637073371400841335171600140529709218236003445231131425650886505216608688227358624241629532271204492371173969837859339549480715301374809593865845546763823398239044208568428631877893057756945799599573322528199394718587285204258949374673030217728;
G[385]<=2560'd279023236836088257776789828493352527866902977639050336686766049498481626183876556489392998284608830524409589784893769205386973676968020401760233989727361742580886776727372078693860214068569071519418200038519542171498220816093421164300830328048660988283425851472862165520616129158257527538911885310514900562682458232956275186752814520305581135419272546596366314091941851782239735887658631751686575860813522594340148773318719035763192029514595594500876818415719444248681030811564285740040289953530137267490089452796595492874302606257220456180643617205632608164188866431493804553428059114627097811316966598823071236001936100926755907137231219934641762080429824672264620488566799246455844441393287135232;
G[386]<=2560'd1089935489575696979225819286325103146118529314825793551003120808861031248781224032683469569913387206222553737481258158397547602000078241511599330852817476012151620280409192027178172612959472145652193241626274434786432073314361281378314464583810377815113966482529985051039687033174732359837840749419439946115933799654479595182036998604993912746826161261662172199594673706439591798250464469426145723836967138549009542441975316989731327944441003256423655781710119098604130498218950956654609150661277642198935796144160579714941511796220685475450487044777367728865708134603557357768802146085078177547454948702421856933396338860010269112249715273157314501582264927459379576484224686994905730485810364416;
G[387]<=2560'd96211974004429108142940779256930945246140557250370221326470107241811593578039555559184917287011937276993403556768837374743637664711225207464981371260317807550165796266567678196554301818020814866190657786627264953896383738388255020070064084664860151998700379602540555373223269604777416606794672657411695910106024818824649717936193715842724205515777677515228505482199470281384821151871681119325608185975858102603356352851578610744008360836139614382255146047972738005364223064196032852807944294990147467812467302056101757199065107353871921224350095720641707059708954914518212869636748166757344874251423051544674689929555871280065560629596499813532986475578906771102266339374140581294116343351910795598848999122750385655522769502878353582235498921178081263616;
G[388]<=2560'd16631095785038944292541898347672254812496280370455955245201706520103338407192103421865674209592451071127605507359053233092082852154635204165849878981380962559594732812643360782989895268702282954796275008535437556174029586046717159685795931205461587323244120757350392830753704914356377498401448502063868662616736675820835526814330981972432903528624792386599094464399899926758824540365085829949551222145880279655193605964722733840068556469305649771075032504330132229122844428426801135556349116339832476516629975905826934362951636375702405758173999323345930904944094092885347005988827470576648631032414871602784397702188614626075079976722161215260784248482750940361657068107326221419833563545600;
G[389]<=2560'd400785353137346596115460704607271546206609682149521948579808627057213119412188085727958431154388211259822261408786770645745726083133916144104295437061404390348168006316328731761546822202778088146008197833362894141141784363899562638439293508081225614323668614463832965046819778262455556293535185823039098975714160642334983405125044471188781605460675859541457051720459034856226661417940901726169854045480748390135347593331544336672303492064318033990701231579784826001555660633555494216194266268874232859654644749735092567566318540991499844493877072758738873993478450497179855831584937286150863654336170361901448542773829895945780561408841213817156678330581816225776995511102819696283864711310495331989602201355200264696645782189776205112349666046541561856;
G[390]<=2560'd6814910836440051220989838121175796600596044167191264580326951941449685698583935097348428491791338055468593440185173067299972164458451551391865153115833797569934111138255577523565785830846080066824830096018271492260201511223237845633115519025473564878889066129922843456174039417601902853721944918667444000689391353387669454784906836317868336758531002504627968860482541297275747554941045442607487238261953097045116393843783147319230716454202921810154387854665182220798620595104863267693941635798791194651993764993947243155821884773161330290104881904111295476071479777067955523358708158327326689354253362571745295948571314528265990751184676202278890311342058013544958939980506484988719213487026929161711658885362162319311868019370562164898588754523661008896;
G[391]<=2560'd12804767449820017847632614557476467791618325434020036711819688469167638325123599566963347271174185297355873968127254398172218615867118710791307371511744660441974318768831627692975146544901295738944411315205926547962429608480506932994783628188603622563763397054500094932881496725443491641465338276351649700623148103852684074627456394606475010820352637068508299873410409650036755934253409606312670882281607182648791832821337552684360996897046518303341635350834554042945408324579329882691628749997748395681218060748902691735052079690598178828700471071205369170041922432135094544307461405409913772835395158145001796252409570504109173760838879486405049971903184358217702943902754528945550731953381528802806557919672596744791246891246594723609281939571027738624;
G[392]<=2560'd109016649699360587220748275806004343607459842709646176188026838200528108551258290603349913465301215685443334753417691083138980797350642024284081232100223858111329124426260085796009637493434956809916478724377389055290096660069014867006814716025307405458441733696938257990945249257318153913093669115616226997464330614295094654728336765438091094276047952985611582096748424040540851142468405363980001739134123477671759832550894209703936136511459154896834578319497699427711964188871344695912008152335559032320999120002765610784544471933967602222830588345284127612282486286924590172963688756617287913367501549309581336489604996503499148666130714716393149488214308487970697550480834982855332067475448919240921949824446450626906367869851184707787149951234260074496;
G[393]<=2560'd6815008326009123663929026005104057870288774140356851546231339772638052323473700564093741694483064345570081619497127089564232539616992787799453659673971018211697959514940243625284190032114510904985443270559061299493046905808594763289590000211432703045550604658049374427622781224584066353874486085672565064622437117527045056454236552364044721742586055344974122508251809146765631204467711064112154143298830726717747425616679949478818853833453621554827670421412156581188734785808783052560356558930025200660126873421363327013942106494159585029976458483277037444381245488874078579883909626616123569647834133482405803314161769973039704296525615189170275561380315417253882123229322501727387275135397301608791722444702226564304245778279629404912595871540952694784;
G[394]<=2560'd400877108025885365940578713010340976505649656893603798842761878908342338019575149885012886291445349865050995366855335628581295944219534200990504067696650973987363725621564837948302857402506152904432162759772358530524469458203534511931919725777223177397333545278819900209940665353679471747872146779288323323683074523445447687900029694783438919550520777099126665943181430931755803850494391928470231794595621769947668899900468052378165514874522542377197635551996668104389874093066769038677353820647645706483807144463210763478178981749616621108356253625002062910523990106994283044185052221368868738393096312483543761766533234970036520870666824460174614124481129628652321477849174828256239683257763178233428957866345552724957341204926044266780170103317069824;
G[395]<=2560'd58856462181295883324680253694024899352254989735633295466412893232666729575246432109908426866953915920006242715329874419159619316501882758222238966112789344691612649366724289343290628790475895636744992642242701850323700801548124726968725288713392535543378423498590724205833865094280262526410513637910273973215418716279572765493206685811504732375759112454835633528574520214686661293799633298186263515146326692899419027647964828246570178878778024274628712833575187006738701476986781812537881185863354994210893744190074649778680931204396556763453757164350927962581260420562083419359353701345691889123517180153027175683625697740676685457679099115028373804616157595333846833538531328;
G[396]<=2560'd3691999855047665944681715133632937924044506934294680815005636931981691470830799321858431751119487450525758397123407679253587090572888832626994011655019311029170691296201900986664314912049440192123151032718294501551039070020946098271723838599283909252340795679836384029272916648843502144512354383441393683105591504579597921968366237739537679874986201798109096626421859551311240680634669679339093757289248053609790663960924050372231619330640369532306563311807094664308633130157572444409471551548860681556723566006713073067474837583063056301195945678795083875405795440831934127774037382958585234012882733688722263722708490298590314475597446266960028174854742612458747195461468160;
G[397]<=2560'd1493041787808189526630419137355951764459199019333429443015935368902126370371429788383988891427451548324366382609437907753494348981960929530884290821062713729951648007588764577745777642453336035304868597309243034515779773580781037568904313532153816616868253314399116628674584251535223969897505558311056474776620954413639749303175458656997975893806453781042843561294427646296584337384264914498698880782464541447176651521326205036151561144211362293502062755355255740017094585431055946479500133049622114663338174287501079153685427639985307221518125203999306368109118319670973906554296496843139547729537208472057063402015036398306294685100852847429825992750989417351399625359232811253574608940020459958855511545839410828845230470099402976629876588544;
G[398]<=2560'd1493041787808189526630419137355951764459199019333429443015935368902126342531814733941902575051930703646383066300677952518675081117793504780131392184545663830876813420128951727318137704324816840792592301199136641088995574495877269034716991629847722746904478434400765344597978110390315371595188529200975601064636072304680733160466512449062311405592395463902280376107766080034526629301246617283280668531211879081814740565517357215372565854320413335957061095623575794724360464243691348578124944289104154589587378426728125998633421902439144837364280869909553594001605476408749392777519234059519282010161107817695381295299186855116594704542912596951284454852067035320097296489890029984834693234808846446907781425770010309781226230676507239317608857600;
G[399]<=2560'd54454047507783025985249257063142195026691018582892565365786824158889650302959761759180363897621591251521948313274797990982449833407559604944349502940533962502369381299584724940286923419699354573883902990082949092930373116668398679784286224603364494572808273102925559774446201664460932798471053177296722959937326546835006846142180113078723117580550484776456772984374565852226534275969927481597958507261035366400867483221513716300738071682019437557000852965392601759132564400032056601877665150605198023891388146313493871049601755693239494292032265553492358919227968916707778411979902724969874877439872794146036234366515687784151811999045463530238407890855010649642891380547718020595712;
G[400]<=2560'd862759462764354276519207056356300960877884527116956796681339931056244773812638906081158618238895711728754083025286869784223435238051872433757054367596226583910150172085478720961770777476546273004505274965110792530709132559177565798084652881885408727913952033726062130865007654523909190221862688163458165641653436175460413905884290996583855711484660942173246588170448639010104180380327473852227021022371360199982029955222482213284335725933315261720374695790537414486304554455181683321022240992780602861268465419576655232688360711332939646276208178139051039679091422478449240058712760342083005167974523575465042020534370465181069656249995538013338768968148611659464704;
G[401]<=2560'd3554603770600170577398359313318491409345385255235375741860417243772272293790017744001645857931504379755006249473795577932539824954125306864330577890584368758013338038103101307081301716644586797485538766697546972443503536536137442561165855962935021005825369586167900610089013654343449143578997308316193786291331520752214936145767257143914879492738237767147654725580662801459241004136967250142564283481954904199385253621941068873955167965846032095639596646604299903238602838230579435554750558952442598537993623555121373961368424157027098152222868771504350440084005714647430168032939239148434149968588935997903345156447902008861953902054899200050933047814854967033856;
G[402]<=2560'd418146076142072806661647774440807452123948664284203288376519325514438189521582194352561449872868147790510761850621086506514110953763144797909904410645465302637412253107126641004103563274583878757802906650286099634225199672177919735025738165016054704430320896976079302505577157913026787186447163376211696355710903684997410817051110715308774091792722237752038368168336385506908947492695925276008464668328347564586184391925591471218445367297540584168425782296596016235510123578500991687048806855465198068833010460803823120160912525497228753316709328923556215289308324847794652060033684992981342732087460220741464254883594111350926207417992436079324007970699059658752;
G[403]<=2560'd13167479080817040158317739695105513500491895454542910997115979167292820195696920533616404251527491186426867177057225608403896608408248335354189062585813760941864709954626455990421363898301080045936019279706926196438282720170442923430142066628426366117391058293643525272745907854552798688703559870996250962326282863367467349547019141435933923810466928847030635403477983800514532592126032773014143377446660938007701305957908067344789094647492596470531022819466292975252994266221191694917670713116701840927325428329188921832988139788585887919787327559887151837252732079061254242576924783545849552357118314266722738814521829216638251950139142628505327216154625703936;
G[404]<=2560'd54251363602570181252200402101072270441645334662295711558434758147152296310700554327701543364834569766098235576887765112169166040621638264975974061154755187852906479232691329069871259118329358968588012093477697607352580753687482965276787784609067773615828259155567849206328362240231894051474670416773187840127052588991850975537476790699876625135278241200058622220597154919984777668143596954653712817856030630412862663280675642358101247497615164003951595970614249860271029973054643758196022300814254294649955695821501923274052003173483719967864746525346632723313039739211068688363711080647401716396689578219212743721400504600968414935174040097922110823329693696;
G[405]<=2560'd189882796098496690197432474845988369511029879101457572603431027004697948127467961557584046909360805703173437855544355826340532356797590507037232018858089539284745944792754241009232201923771014060530542223297418704772419623788887836408891002658558443507939492804153390874411832542176092414541432788798916070257166706398876065050075288541756928526075484790737872986221161995336548765344731461844559487657345652075581910203262672938715641001682246404219195692160199889298266115712397784815571618415877579655267679454352382155204635513879458827250566235503350433231408173864520639313404368842643930713475734156574902521912486776468869593530462909366495808061440;
G[406]<=2560'd781990368303030078359196724291483127667839304523906606318060677197288051842131535858223309185891565727243167235301103585242432915470394644862287069768393393754050428841534322238709688627611574996004619901301424771970092809178034732651013120562666787837981830455805048923731314762511584336029503409648873695810950445741019810722259275458675472954591511817336384017776939941472295682373320793478566849075722067721347834564846175947240416979298658382096520531076192693280573289552646063322103863193605597519619572254355128591350970489370227587104596845271761004112849762525837451930429835203834816258600977425930138832616937270622897536998763392645449383936;
G[407]<=2560'd48695455434986421465480414896175926863966434814920069790906724106928764660453846758748047903419062512135842423890629862722953816598388441996964272841832181624027960525907523456732487124402244843662386951715642673602166087426309100793895899555301531191279476625746212598052620685588571755395315278063990627051923579093045254147935218868477805306295802705190052630269375857315280550138378296850387721940646653657329796615603564621544206500802876089207513742320494498435738351901734321478984785181980121111971057252686250314762608290851945380342821995266465558312797841309071406472382783435258521212958350367311906272627316774382383030278985393919701811200;
G[408]<=2560'd190216292072548167607381701222653857877838928407102084057400236602703050388264941318822268263946740728901040722991104747049284811289893915447741657911912008086623208344470697903757101960561604210081877074834478740048191368341736356459665209752166197425784936806567620291282949772199094594630865540197405570235464249364803686001173607994797500567228726588154909404357200860054197519109674090197004210286864417906231594691430872478844328934140422158781547375937788315612212622116046236995703996286724641891926355125371085838718392478599563602831243032822672849955733331170436674489525979730378063961719122712876206206743612326930400508385446560014532608;
G[409]<=2560'd11230671110092207112322984547890939793483457866417335729882341523960568370673023966672873401997583746144008755164710562176236691139031401217916345998066361985050273038758411432005134175803783219653104449129375635893636981383007882969823911616836858429596598133265508112683078490569929939395436413793687974569253173003544919253353204206831757835167597267509267879565251332862125347948162722000508221423877634746311509171755932178267589341181847887960892297185827363604475616487012344207716075234104317613668493681193784358357875368903963650525904459434942616093867550820344432265514910465385356033198638971613709827226755696171135023447022204142747648;
G[410]<=2560'd353388121884157953162486170473692293843033106755676087273748106100233176799896360171866443962667266649679229861116259373601823547751684027736982723402304124324463863361671570226908713187134891644810607105990961294095218004832258797896030277578022766244141141685474971777941317326689544093424256758239223702970758890695795463110715546109224744993439659338233886456932841831833947590863304608903664035507498009443064962643878294902320518075867887969790005263177146959025950057168079088373000975069584286990868449028923274966111899194279928871799238025105364677463671931798508877035303384730962799179687079971267923061467671772170270192870820413440;
G[411]<=2560'd12085291463313101001923473518510508160510972280974237465931984750726764640495820801284879731979505373106210966209950008546549388061482761699909171283672152325614946937928951453307492573075289882467878103586186197382086946656183351648086785728419204462667798192712174746231126216073728477396308873709988215769653376332383777899271268250628039171022558894023655996249296141776896310621564442559746961192877545135360295359292809820868952656840674279630347926724736001710896045408190778359866726286969516131036226219415995542447102876460560352492519743527064381022344442783422346549929752441743529590584363042520215412138120158350234422631645315072;
G[412]<=2560'd47208169778604693865393437337901749143273079816927695950337891238931559863250938195181259520033206864714389471265285147242173263354709938910992276741853661147855324523948741114372819376372615876333304947125181563220151496855116573475046526268372687891745512710046026527847014299448747998598980917746634162378794762676636951900553810831603973890689117073947694861316484714413893885617621058257717931618976470226251229940604731105991877826391935898824271117964516286724222741115546524086971352809455356101104851359824997962339144314801207963760224373563824007846329080463362242364771171450072239746600721806188296094167973724704268431600386048;
G[413]<=2560'd183771172335377129023147843921592167878081122243790383649157178779758889576525030163045210922833035117036545910704782586375500740748153426846314657728032983590027498156398500995553018189025833812918389334086229955804617671713580447461107232352159204069729046159436277889237833755713137507432582276284028315175737425927781574397791603279187046398264065409609046083565613760781100579052842988901216897391691310413992982695692571287698271953232968925395593081517426444066843220040703108810514365065334748681006881825336261008760093341186029848052371947739775169219664693826935945948437908547964926540735293440320573401449995642922194924732416;
G[414]<=2560'd1311661331353718854917495765775617134761517580504000237568875479528161307181331061450898385029366481654917465199763421378467039217025845351698951592677747494038609576224764487869636664738053762323358587545728568196800942939945741357456377270048532963172400053917309953352123835568396556416500946388703403053158877778295441658265225050757742588707603068867848602825282519774463461354922055006917176020113559478500457281753135271403055221971828704026423743495599935211263805821146487249084178270959264540297678030135182316354427994764685826791562494575212054123547022609896600639513071872240928059036697154433021323469176007035090481709056;
G[415]<=2560'd44866008861688316278356006068964728526741371832743000349787040378394248413834583187340626873136985032338087073322660614162118095190565000515771061614600607616321129769784285921326420438255548465837401734250701135840311271226586223015864143481801959281683945359794265584261220780881002365791727634060224624047985868291256705646837672948350827888091138528823802147617226143387625980052405061446460506100072299846378643137502101797451314184008228472774286240093956148764741179316273150562650616003959354519691529993950856722732288914217053619081726368111728800567043450967359701500412632153087662146006997171995540404382885503667292602368;
G[416]<=2560'd175864136882119903527224338504328807497403652721420205343223799490133997304233735919937300633600833428450955353744314569238319116277561670618268334410407015833083941438580630603295365328137207150476726551764483421095101364930967437945297732446531697029381589984910527966753537652146128460354521189071554493384282344381615183873611722550090664059239150563484330184241310734765908066733073920906600632932012176790541750003444668721011933240594536272855885412294473954365124395260740612835552555598908171691070572259210219524970775129511503222032107807962282355045806739440626102438121115859013585325465820375276145314060011182151958528;
G[417]<=2560'd649207456311934671352940814733672112750689567363545427473052128078848310326531611439229755716718070969601770261567649164372808129866326744684818560374514336635060378283783216639930738791994757776352547416055095177632690187532515156509592828612206923391341454387369540309248217582218149434033538571105112231272007193235902768778186347745635043028411983678496469406945613538902169476052897674967606351786028708441638658211145258864353209377090830111363863572486678579510847471637792343171658766287166049053401335463870707181473229363323050639233065009901808263607854542898179794061966201431597080384154360893259947266715412600979456;
G[418]<=2560'd2665581518493582600192521270334081101956713046680200175430111130889646243387518478478246034714540987527472272924042021416848175724195531196038795053395469885241797271509301566295030820224070756221328215937900525240994170653471551244069288720996151004766783098371532577722260462878360038742403456871550955564435288417934449186531065171261004783051917347886871930115368256638997141674308769357807895302620342746609470243880686074374137765714450855650660287182268616045160897484899014527865654010062716134340385057005640371513656699157328376683883652901261581523810586246529042702940693645861941789935511041230101142506625394802688;
G[419]<=2560'd9867838649083348961383117947360202536396008939205073965512728078310014870626085008376041989371641204876961233619957611347703981695399055791974777979382030470954822040974702296514374605789757326223717667637663449800688740919930345726594974795556558094366923045837557848940501070310892767900789840137685410160156631878229284748968434773367657670104493024526172123652579168094815531027933872719908578544621827036576398362503207623551122586254076690791998775555062029399354816692299324018369660841638553221265771459859030077633227863369086944119742110681444756206893873719442172183133846885492408634622395648626722818804739473408;
G[420]<=2560'd614621988257817817252073664607650570613140151124293041016620088143030603238392144095700279357285809717791890027775161125653816895791098494220034456077935061116181084330367066340934392087843257999570059396866554916227568671755835573183713964621768002199281068882057705408792230349463664375440469383040541386898650777206516977096670993833752927490137273026186355028869841005132956393485393173299982775514073590820654563766208381116399549245655446059162954976452019357402075829575658544561454535790073770944335004232012114259083657353810030906189099940089792768604647694082171598613700113769008329924171476296811982604078153728;
G[421]<=2560'd2417999329097099916215676087533862648944462021751167645542637104046497836941438133340362126406733728339249133691338694733596367999266259274741288846763407062258435697598738440603767340581688687271498862974690878032767535932725257636021892161030538093939384004169464620957105193311895440532742772722208826852458989475618587303477115647210651108350232799334596954201902683272622118822342195514431527398615759034440761304419137546445379973664580914251313866701076613922592584560837862625376437039869767674242416677764351615172135844235400490082731256295860781604173986057243434159268335671269798398428815615968391953159028736;
G[422]<=2560'd18235417675525524868871209281670982779006540399354570754025529795868144852742933602160642756631306787029371175704850299852179067074623843443353606822927029039164764131457576991336930867184636567017876748676173329121352757341629629934568923965448059989496293245006699027986500949605335212953260589801775454256283447254640172027437690063017541458095822780852758151073096918403866664517179410429693689123870443251504056936719552399604698170452828491037437082437235265215575185823326838704087222103940067271849223280235443036995650775279407822983365507612514853305084136546393258018679612617881128510275380847411110896205824;
G[423]<=2560'd38923444618390563941556505296694389560578653808393771560941068577334132681075200208915958090407251226775013832213138599031286959407265190077714142760843682863622244215497469491914972094139573731607050396133733741563294588495465211729424245641532628639571863455121117045091959947135404290025395604813230579020803139795631902069910361966250000858615530781872895832774185852599265282478080073471338958642490597667890037958682452680867223013751049072216531105573777822627724928677135045164560659548246522645135930753035170102605263715361638494861604766954630765398608865513147818065523542828866023877034597466796653019136;
G[424]<=2560'd144122057343212079671132011789414135931280991204454263090950091070164564657255483536170107808426531268903469411165860395565681072621808298413301611466047698927223267350492790692421706942764594034849273683906725717869183897938773685836521640861627511203205192410989499359428559786344372057409920293592718680938653350638789875675494665908132518125661471277725011864698162006529182662246037167371705058974689269415222812784200041320252205710586436227671255632422764974334829927919195098404561606392146402223922113612593547820241041825882096090939213896954647585646935627156909811137303774999376313655315087683724771328;
G[425]<=2560'd8450823270356355490187389786611762758450588210052241976825111696492936573245091711890433497840335510560843939682415120607245132038268750384218851663976491491924138607028759401176135239482660065257885658868360242526045147657782990270396370273850112934841483869930152565507272987511399111482020911183450486738407547103472385544362266825617082343952303321492774305959028442787370638893516230660740018549766884099406683330995968448905637553816010011322403131310986666324240327031715832654822196524193920483291385958572071949458808568442498692134094979258930920863337803590297889360129142902395304612316845514625646592;
G[426]<=2560'd2191100219964868343251200982822876921781413438177563934861127948492337007413222619309883803106172037745626381798764340440249651599885233260889092911340793342237652056894497621236095827740042403390128307183398678156723379034155054191505406613694711739257547639712070058926684114029254654385704369412834662343522109788614992816744301394178616164640458641258312932160372411843987147995705380737414079502805493255251954291598154862859113256510583240906471088126228291983573985081682841726325280790936563681379098616281778153543494873226680854545994538785035002274386332849095011025569731836500480726871678864326656;
G[427]<=2560'd136975237328983873300432165710633630479984703493298739902506942820231052713503490548364135586207913138359005798652344248314307643931749912000002178478296954895781898183432667612235486515067118942277646223213258662605111082258110741041916488481761326700495739058363109826448939679830316378195450612959474610453631816079852722631299811915899510839855401088692683200988867635003237792185611519804374604369116114680228916097409952748275656857424618434929589150111896197521994779766060728765942983304863801592795429302996128834507464857216870720770185028378842339469930401690786578807605047619470338688084839759872;
G[428]<=2560'd566411114964159908047287359688443423391573498858615818056383364505829263757837967020307449623213418203262481513430531647780764250369687203663271195455594628978621616085587381477388458467450607020828859546339109503666956431796573964893651483782520130218515272497266204389537773023521637791279066495949429330219806664433968279060581713214107898874434909234155398451371396751301549606867514934957195083652307479100037227397392443540404787034058772033749737080552465888995144048507475980409448175136262924100343380046469879100200510784675977354524693444913966032590991674458842238938711795743384149206914564096;
G[429]<=2560'd2097253821942714468063510913820096631963095166941195717018050536356780203664817510245363507143976140654040353499192640887328079816875354406330418753363298376920539825242623014667538658933024083280403649918650597566809866274684143948499866950775597384029462407389340929865875539437500713144941452173866663253931670699720403857715077757097524789774225530404189305893794940811427796776354537025298899713961765724076677540575187510541862737458805721641608972963173696428292687283585973181656106273425505686927108449262273025311582219768557862085469805953877323221822745610188899013041528761219505517498466304;
G[430]<=2560'd7687724482730840618268383820127267030730070676450039415483200355659700170200549796341013970552618344549864215537379960261350760421840978023404216512062325789976672079802829121464851241684266300417633880926809433201750266176610370928792521750021667817475932561202390123194454365540710304910453948777943312576187654778203924472932153877354937792232408307629314952586061713353311875516936398906207171960103546016411214668421348164975268347151472117777455054721711256189783807954322735441644266343328216811984531356596831116948378574724429300572656762089610196606640441872833965446993306707743875612540928;
G[431]<=2560'd31884733053575794003346729589434869157750505597436664408364970179656241472878201303875259579970962397245180824548260505993285962657067273346464002261751096995626308156241718086019311569555928426921649168156274054537882232211323778370698956561648028648976766466219302015686981752264254384096780647754625585228765459969801369389052626201638737401399818926383362129163871891207825957337686907763784986151700685333296241038721235192664843997540106682916024800875373296235393067765006597086113997168357799579158180469807771352277201520909353927374322700410706260676176638202250099080328935620458791829504;
G[432]<=2560'd131877759614534645267330563836845296388429128579824446920848084090195112161362379010441205437109621906573958512030439860143039708037802408692360803534070185383486440970057646046656608643135867034047085245996525648402304532936316353096396280166812548028797853192307236928461783330233620262788743924775923676220736133281863631489428184837576793176521352118664863915243714875684068405300471750931161544309169325180953705194177197321385844205986461804659005536819070308923777232228883006655450452857183260991787603082045761995140305689247807385025021487141819483052062564099334924215563548191287672832;
G[433]<=2560'd7786147748809003077865386273987468093383596827728083700393910443325307034952244738668825234942860792801484186206154572175083519848122068072796837602444291474667965113428266101789678790476922132619923401027073335640137358346069912724420633462352078215022614221944580486567222758325522964108430077117326039365765652174531209281940380448398498818885311042701762787032612067015811407685101850725298318525941650902080548629707173764918436412670955528260017821010630978973860521119728416009112897055413226131611401903823759604166502826454716473565228634331140419050687447627766971773835137718071328768;
G[434]<=2560'd30414639544226536895309685029687086649362395516116202492744441808548221364087790451212783193374492241457135205176743358780434757224913606965069503945896283878619106932566888263162350632351302713331304163403122883631924516438050528129281911174997946297946282774742923941529399096076554306780714971010173468469806599546328897687815438314599278351351689440943938785009518753646254416508043554861252209555000282631883912248874083638180694906114006680537268812121905933415845777979749736109542328389455105939271035711661662362812579139857105869954840785202447476279582038157594146706066726096732160;
G[435]<=2560'd6990457168743211582723418222802367476729289544626533691963745739293933809366777811000862428187889141585579068582525624263913883411090436937357725963446149688554104890035764801219359771251935478881853017435189419968868153827366682523613712384847502615656903913314499978456863194490315896664122329143944598153226775754754117822476412219817531581963609028009723942315901305706330547429407514143618096843390559138939504432497518320650063876379046261832273253883610292082750263323667025283519260592572539930769089131116030740892707428252663571315830018184526141164590009432546950823300084793344;
G[436]<=2560'd28998995779671344259817188915661462555296675395702768223921343744674997946318425798789088452145050893849797612965432584695557673507444627203556173679621248989237652480720907714424751530311499456214880982776939460429529136664137590515322892256972874701877951502993328040631281211245379192955978526529498664287676178928159675051973264957631204952022680187419879134190944026698832525941469050774030682635689972190371062635634065298818203464210839456948652304449896346860375724780391557415155330651433093126301244031408205772044091937881463021276917127442583575255772857289003050566665895936;
G[437]<=2560'd107053298293772992817906806111933465632776443445406876148284359593019665757219865135353440137897821024905970720670873665986056686039305324692686538617563329428302521918565318604587999491034083920414689888884106800948729422980985241864957862950473332495578249989047612390432814590522053724913229864928881481453055265163165586851415312815782089219777919840124385596301878025755674858590400839644313716523379093336802988253913436418035856347763464508028500644535431373925287046617657475601557957426940456008536993440046790585932642158207329774100500150311071000246704682145503224359026688;
G[438]<=2560'd442590837449500599981519648314114960093641655172812231205515249378587410071819495021649560172961773669383124277168487870973619621108437753158165560601778665873638052087551115812889825330306338494267331309469866346216495490921579382482391120546010424497635130073228457893540655284468019290664830166198775091750275839184607047034702270940193111652594167009582276967365041159765683925748097904594114536495411385565064470586849584792706513724061490390555105485921813187137044944453031958451238239531438245606450699070233505692854657749446756798766023051268257793584640543739922050187264;
G[439]<=2560'd1836084074759532569995027877138551484048119585985326447504654387268221438123886574512173297056122404125318094939812144622209495883810442427168664038679916931805049959924655700821838609628816993218713451346688342305042997150621059694749573782924999690704317794823099474381561060770727664477945101904027270860972731151805067591763812854992811765037938987842574768232630171276220528274170885949271154430777108563405169724628635070335374890255137581680229139506755479148182945454109705622121622851875318133295927925644584379106939026320830438248450893464291373537225503703854215069696;
G[440]<=2560'd7172203393448820939714182774628451379751224834360858683373250956031558924054958818272259236568806488263302590605085281825522145015913216418399755097815138150142589086005505407414382582472009339184154197277452973894425157494388798774208484502057360359724446838138548033026191095906795503059560510707575754873337166153925889684798095042877475943627793736976068439276366019562255256792018504716825565214621666588817927643422277807522305966911063021537454280231213442554164360251864334137657122507612734570179388574520503482977307241639640578032946741658729458330913045652246102016;
G[441]<=2560'd51112161323069988331627226215827222810092816928409239874812411820556793134322393338217069962708418068657126014948622209920291392850366686974182010772284083326429067165277774785246345211735949470694488659743275161792119008741628719344904446973369798882619079809478050189881988373809286836202171472887518966079830718065197878244957992205926754554045229963155072755242164666539938934259894730628535421139887480026272546023914655791437124339336305451694527289413181989727887507159184559112033946521268625581521018456962314377397122657042421521451303424802110104195268574797889536;
G[442]<=2560'd199633299587486091274277558195628147385305259888871243916227504553796778955266918398844160221078340375231776234956421507132802424964600864660159912504969312107286085051618968420687910863735015452642798986872884446822380282160066933100700878308086864392159845065230765925083289740913649309374780144357627866023971570388018052346072741615107574723463931156893761739500533868703738759793468404305305414078951972598720113410428188182576094314795078805195094645953670283756623740343738269935183724149455077801024222498050107043194023630946165815493720092239660676042575518367744;
G[443]<=2560'd6415478822172442691385804424849829335275437240168293701322752372327057503900417050541343527396990503974898670459630212729872494857954362082170004982706656956925551863303332218140471525641811572039046133428461077716281897052893588788910488599100686326334033089646441060576004990791483220376234374952984583936456020945299910036920197815516684587181656437746787386748154614657246160569700781094623916946066197409184175421777597671565318194670604008893000879547727061061018767085370404826212436957275054165162414118517315735899995903152310092126615478089476431857256081915904;
G[444]<=2560'd2570999922049101427810624589757922076799569653180204733358992781382799042034878782027424319379434527126711106117171551149820849231125946237017585233768738121193778266252791000378300860257087733325107410648821340658465957308440578972576395571558985679268447875274704790428178310495268345107590139168180888173049096317510385420846296267438099001960767371512879860882064859191481110556132511437870695747251107643372459792575875225539347946592620706415395067012317184;
G[445]<=2560'd2527395763998834195447003244848063853665333801896035250464504235008559628584988606457057043391706961051340913841968946793436386768992044479871328251927540430740023020954896510537439070230054936694674253566460684334529257272752629298340383757652410215916376914369291364528372575686706853451733273427170629313580664947569149949057500735577193153869988367960643908268970077847978355625059246754232781167879206258337534506890650408101732429948292547848462450458540097142784;
G[446]<=2560'd5935696575181333391653631137056414439340741311899988945558394590919319454037270122115077384345331547087937985971750382275458050433999320639461061995483760085053624170250762512835773288766513860058263689479693350236960683056570341106030359493653640516922874551547384147996969433004038158275433630198222485042248453056150621693368885138432122296719127741495475828027115937389169777630326600152391562438904949042308021339316657660068371138285340444453768298345004159439708249590090494462880662379424904804118743910236800168956110624698868447268260081285967184146634570366344757248;
G[447]<=2560'd200240922278232540849726515757695833016074064105555419586077630674078073359514318033384219625193150122168030950282630606867592104255085393491958604773718474647094352648363794903855664756699434714116340871226436957160526197013399364211831905507210508045409892893312341364304533647716195218987750301165238567759659285078087764542160703426747556715326353842951206742901561002656841753161672699767536430899852188456551060356317269313846188062966881735718128607110160587767231994332562427104851927236608;
G[448]<=2560'd57869626538409204305571641484234199088989820139015679862063956769528497758669359196777502821589668255915338558485664205284960825507918104779834777395979336882189483220789055366193760084537380160827283436113619141580434508905523918099390610989767888997726736869313699447215558021063504025006291708015275842406498319699183010893433815568650257945683315860947993284073273729181650485169854497506233756559308889899891682511465448535207213464531667866873490879423646759183196690874184808946024613549178880;
G[449]<=2560'd223914405314576582991685433713546748905705260902739850180423393596558108399678035280180151434251953352637256804907088753327965315701802562957564530937863613210785647445426615686825083683696089505693545348768098112684166478810457971752033251679791570724168813627946858772294075761779951183656524424816787600519774971155957426090222917539845107470944389707144340089491738199125403852274498777952192244344631076395361307091049422656443739754085934657071182213725428355146331617016768522127235067426707079168;
G[450]<=2560'd237091872442920152429458039367608939986687657315386814375555048119499810060053352816308669224658846729804611918523629128171985401248856992335427189479149862153785207013764160488007349662411632428862366921316759666813598808021257355094193753263419490456857542851165644895394878959699292309174130902434752159011097160599792861370321499026572315743822508282463255341714283397009530922355067588215665133886324359594554947456650506667705969021228502002203847444631195571579513040549243807053870744542115790848;
G[451]<=2560'd4061368405060091411110227704044861789545090709218669599457586256254496920543129079902935394722253174313662485817655351574376771494226819161780984003331040582606465770872482159202435105657528364394183256761475144899660695053983219273489416327456784412833395038033819403372676704943418162402731166079824586680801709760109775061090898437123544459177644442376735766817438084880986221902989525428921662530986994536930294787193979550284711062865650648379864727176270146942242454703368331634959967105830679852292272204773127161145982976;
G[452]<=2560'd259156520131924496662368514636484344437290429814358704783398243833470161404677611549870512400749935984893921870008731899233925107730229626619864164916558618240972555685894416191854863021240697142237734243612834100452977030662461561160365460934370587370356304889602995806363924253383408227217278086387469422872614931262942040095770856357080739739822755978587261666018170079733931707699720227649913660438614262257692560446445491239210658059281312737582945311255789712301657946798159612682841442833810141314259171032214536192;
G[453]<=2560'd16926499725022794571975914886494747371974439387784807282019307431864964265911406749959556206799291061544230678625365062275571946026228528077091783261259112728384329990120349447526568103320181103556427601764802547082188117005492716176536678741618413383994214305115317610161338308140666537967583163299692468339032057094173314934075270379801913669294789360184303112223178585359050403033298565286165638276395224353939115878696832777301431690617494148786588580196301593645181759300667686730419259288842327582632898273895915724996608;
G[454]<=2560'd541515772144588423057452285801975925394797829064712875734575371062907906953358582554950369547356621068875153666306127853440855746986163865803281295829285347244030475702826137995850150326848233779112182992229647865043260417259239433585243588158167772302086877932494040437064270363320796579997138102633256692453788297917605428525126072174390292369955951125134810807734305401662221563039980945570482655633571932241499172140654308630043134364436206382570035368206557380056516478054961172138212637506546614935380919414034502319603712;
G[455]<=2560'd540458140260865429959244538885814854235108406854623886198861409190371681419884888546841942724325271033769763807297470112266964463367966280433310021803130388472860584415983305952439892110044788453940946906620985779191448836095172447328841900139599851030898357926408808999548188922796351290978112355019360798677579149329902902092821617895755315230124356047771913203080084360373777181176112441917882031537708788344314192837488697177614290615770192077985858443284813521473718556765881654774585923686240871229499064154188994544926720;
G[456]<=2560'd5148396096422391593693210985223229948801183492992608227369323946046571732449655968919144750263120290927731619490550057069169514345803180878355113508912121465536504128346048803546586007534195996790240386907138137368026304828291887990441335709457591138003493714347746164547597820851404101231841895168911536784805676027879155219118696168869726296715744483106540587250810835727427548367510321337165796419762013236770748476360308301649175923332805375842025558938124132006931860904076809850148118702653006059094398521235458194321649061180156519882184062741023555584;
G[457]<=2560'd540457881104345298034751683004320939014265623911169199561708504745570910673736170903213925449792339825345750192013605983694165758530947280051327086405010051492853838417370444458607632787479473060218366957146366110660774592202057061763041465001401252364915258442078583278461471470494134514084600505158316962565080295730328706587946630768500645882606181468046687315183785766074886203139043314224987808084068969458297234494087729837585691627385264981240582397539881024729763879412402177771913174171108858789282464123835819663294464;
G[458]<=2560'd2250297766757528060363378293585466094909643757097628584125300212809396786629648978675107528687434264065805909716933873409112118247433758775930778076439384675731689337155471411861268032995121690307207800787092740597213301550786429856410416017749721412417848999335223950243971096448926576861247855530555578028716380307447389791331162274252808261912941749327504601494086120642560843053794888031697834777840660844978720039517007171928392204101521100026042446374465452998548131278070570996302668278579761812953604852192976971862815836650860506189662786861020749100394644879867266621229343257607630926246192445393300775292108800;
G[459]<=2560'd38255062034877977026177430990952923613463943870659685930130103617759745372704032637476827987681779675160737753933531249188867250244690365388104509712140232899480083835658999352571950696720260952409822501085365349827937117804683546192254384938800250771891269892497179022220514668245613993539373870265921013852573923170907750019121586404323920591055504721712651864328251702819993793149885566851796554588648918015643367246477721539934481530975179833165695953219959152462084162995328177145745075330507698483385044226024248983221274726457028958479685408077236747864240638236189182396483506750354101208191308116604791535542730752;
G[460]<=2560'd578194155599816621627484493316547994268548466529555391497606548797487059581520526075940878236620957890209353950297575690556175103117663551561542462052201473254458502115128946391261744042331387817731135145890941409345007598547426028425781867928544415091719386100021629981932435004259071435931439494790781193305616426386684126472251490062128554383486111425018437859611377744598792386415548124326044221717593243747513750025064469894055034739725294218157593084968185397291502318249261883934395706874407678524046988114311979098929017852420577077718466482090584482629755137352603189377113791443629043662904000508604536526664105984;
G[461]<=2560'd17892249913945973697835124540432957712749807491727780027002857620436413905766558647575242727400475129058422710362796159695297865768634597641993173189005032022900344170620083372229932931555900900233805991461453681046629609408665910581346646227001245778169129650961853874742667970141775720422309770669189073661110631662033577056060011900630219334749983728273865692961263206599990422799831371834841450793640376514150784295731819907930256460373216385771822210950292743875662492176289181869548816135839621224294683813744831331352454831735625921276864671776085794556530825349708312683769634499174257890949975652434684912110386806784;
G[462]<=2560'd156692734094860193899222757338943175120748314094222073569812904440837945955972595370509221404245306525125748473206089943471967458935088533955787882061084148611031427744110168865128689161021328336649808362295261341481725767962178651629486466824739306633219152542046466207329410193653492170953509097402419084584210525608428976247926379427615214535186680970620426607785328433281200597400076808352703200735908561407380080130278771413845946567565301317081733474864794164371359952173548939444108917494159155918612016938820113051228941719765085071377178731999907040607467775870958846684455204464841587129296566820763831045568179732480;
G[463]<=2560'd9096567331764575249338341290715964118267998127207668515915142038468677705151668321797258846832086143402953483332016347708320295818309582269502170152122135215730839937575887007167754573580630387418156459133592515261019079499891659115918560837064983413153343548161955237997413851141898324311108587744271240287263109761824146892724952305591134553648408178621174706014987682113866069432547209848300997373442168830231134757952619282305731709241808433702302441005320463342821568831843217460932913872605013663433926023167613815694263600809543229800137869492395570829921238272843666995596398650945328534252860937430188303834905246222516224;
G[464]<=2560'd26169656929204717414879891957885217106950231572101753495264102900232206525635509345928124578774994910368010802724137634578476214282485102568948680360294486441102000474363655577959478890710134971395886786586525915476696523018611854066384990726898682894982011350490140953015173564970752801234095414972916446094718266466234087062132240349471780180642896179669271078426413734504248898450995291224479643576963079822567015236304476860478919588896914823346991060471579309742240161411359100982557654503039978701150557468459158364362405522770909527545844991985620072140319633216091542420813835983855331969024473535922498222559449501878089216469838201551521313449716768348322362480080281849676422040138703872775489880679263936434961376802404556064227852669513372794880;
G[465]<=2560'd1715054636911677635422294878265538158479251037731161574604105718356279101409783205953049692816438299118657994374097321898870286526331013614230960603335725656586616254418120654962298556859794952511078649399636590747283974665215613257068199226126740574921838220290266990167442461057299777591807046188289133133211290556218280942878895589031718050923296314624554398254486439055641937607543557296087406713838944170721268238585767193131173545456784895374440365902236068622358258367343874512162649756470436427878385218819397817602603560152802100305338291256356546476287304171264853495818787168097062778826709549727304950432532771167175317503718562274992634450949341197121260064011034734677468704687164124612581740832367441401765947970012519977497988489419359130780434432;
G[466]<=2560'd6414033728414507668645369341665142075358108520508558082234834044867338155889710105995792856128985261600988745265221856275393748517214419189588307890752554074947187066546883380326881423311668835448145264103047266748949461103272549698630168677559981574403578143000974764554918602723865687680340648467313015841782783612473444945167943677027981711854909069622788569746056708161765984251266938162027920354743680129509268877792849737399280771872056357521492634561001284470606313346236524202203231516574652477184166760873890030918554661468381717008222290060127293292186034814326999124281549636911676365465641302946372395526721687216330900239041770001010629658495661854938130475696917686602689008820980489015641901726211289677216402883498284241714065648402825216;
G[467]<=2560'd6389076400131688952283448737246274975290435855004668385233278674386290748764204230094497276889901313533946703813967616512256509906141360196470898191656577380832601357339312133202601711473785109964054389581026088328713863340002936265435676944495976982271777489413445998019768626966316651603491862154849395272150546522331912853391063666658350323832001889167793429705882870329774606940912017263640027597996584628948686643433761660068834592831429934753875971714149113199151936262500844389968878238166429751829603503176420839539266974076770285930504219411128090813460205980522965913560232224247819628386479829829793087875370586529369191183673431108047555451646469069972444080199137047940758506212253031761486392001344724974849854320286547531830937743867772928;
G[468]<=2560'd23801164324326889450166993203196462049195877899178066839328406206275736716792504664642063710205066084643322872620848213614561601660001783772477809422605512390736123165302634589293089195442460444308410851421125945951614862158762300053357048604453253880916180955048568963820053477240580850934817888146521886579905366237100389259701569389902820802133133427279047268203272587974854588844295034553673506497922399532725525333834216782648932166207752239193302564944008473612930443121924826329565003949005700743238481004270316635006550033208792426611688737909460733116486523906276041058317098804328733833351519965802486548788175237588323104999781756964340554307177585472071312976426155670174131959592611707445871312406490429381380640736521506545565958144;
G[469]<=2560'd27081263148906986145549132614622857820845587151436015033669738248329783679323429629872510413382199494492709186654536608767532210106738659793195730012112395735875064192337375474826263468810581690072685153017114718227072447076279337753460979798624130612745892234837033321824899755954883426479591069775961465157473175112809341949148262702901814114130602573293509282855130693657938369835981434617094344719329969453385033992537978259657599621605978723002198148078542842974230807193307797440240968857561044227388569244428964116502940960923455811308274048173173570694058871031736512792215256899230153606581613961237473629820060525195591507219258635848871405145016572505709220268130159801775096176868125568143990558979713102273766163306916850878664297910152278879836963747135488;
G[470]<=2560'd6725704456905100107436900048412759051446299402703714083074994243017234843211107378434145240430525672609937421601789231315900479047501268911321559462641114195026617233795307896913564805300462710388341959363099802227515220758684483681310646768843661400853022354993244658153261904180523366887949995853073212291435016647439759200387183738751981927622746791856499742595267172667444824245488643228432681043450662292387821621260833006625257618524211554687692483898785293199283031438948853715817889874169750395269592259370764662079808616643322588441263111486645820663872892665550719515230323653885174085306026358436798135165450985959914121447509581243964168147584666914205071264400049879816013129857323534572467380493525338767337911394834063854750815642495974100697088;
G[471]<=2560'd440775767288133517749010930110449356177159600153185550032804136582307805670599195049081805596033928074933671021719689768955141780051054137084572029904856521059186542815108973894817421991055897505631055680565700999994633116682851293618142065572897356338973862059602226159204836977437376683380894172724569948986324863977870090875979399922672476029345816640235462461081256477041409118414018083525460365110255250530420301761340596320729697006630785658312821731955024445406998197917856370167015754964133506517734395657592395104564815111739166081503358362543111203460626020623946469423799277496124070214536286660603188220171599657082598483565120385783711173526425027228133893427828268134739808433877543517901324853048080865902894665317565714731471079651193816895409094656;
G[472]<=2560'd3611274132885632135436222191347075631203118698096356600648985584328936621180693956754555293180823117171200928931701583157963201801731682546419537612132404030768448834542013502006923758251949339597895433493491895572169507480979610486985863655617834465050224266790704744049937662730905926714669294747418932929313686987688225859757041087127400701404117380522359737207119131232584467932551479850642956050114134392360148804254513796552079760718214645274404159039969671959506689988104377757742933399398305785377907523582528078851733420831435337189527324851923499543710989415288240646048866491272997447334534402835443449000581200240141953695612846550736255799237619302191000677862988998946188262230191157112225784309845513641195804404500113857345825931690912823450681577832448;
G[473]<=2560'd86660014506053368153161254918276319667183510037263371593354515210027611401429623672625597215675157899760712413517760997958564418619600281571547909728778637084935034672857251246792839693749112915548145542685818444857227088007325627714861116120458713585499209342042936794773344711861045748706322617558313667420892598163050002472872269106278851215981414249468888004607957032695424991168796820876406026156325229276845529372747709540454003415212121226887004200574823528865633380773427304154210251210589343527590591761256034761211453735900983389447241636888557273854170796060545411090024735814376945619075864618963883369611255492026438758432358144423691383019478638445085191155196951802192480187198032396200776404514624159056813851423807681314771815577878047372027531318263808;
G[474]<=2560'd86547203451807617339068553175111847483203248429525817925444716230171122584077505336460183835223075195579935896647589667133775787201358275844452731613147779140537129034247911693420752550806061261973057725215330401409033465691871697803938914915113655263068197542397853451087989555341815403220522928653818157559322257963330167563703711463263885229989392884626068605532949259865373988334412826892472021864256403583468650143782602648661390489452248002291690504996016593855628566407889617696074888433589499446425289001575419692008989639887918721426629920868010780816114891291026836999302419840598272887033660707446724120907226112954666857493306230856824389071180727798032686032180872448723532096375730563949159544707934969684197316312878433630220650703518345256768219543240704;
G[475]<=2560'd86547203458561133094776720231015508752527147505387292460086214498375829629551932836911835896275577965464817477833785305598060528996253468261713745997404624106324712400663521481105869744200456599545208802379383745249173190579021683556204429920843148106805635587726913121622068283165672293431221898745970736783967907619829920329414359650313262736283960845644333173988129907441357031578420729082477973058688921896173598136859333728585020920953187522436364897995680844932021656549708048061875559008927817491694370254625643475023601763131742959041611675894143951646797194990810082448650167324845751021659095157708558113519576871361157719376055521086115566083615468799861375315452082371507203293680567223302095129145936686004225646219965136980709808996436443775759674295451648;
G[476]<=2560'd86660040339956985216789991750574140328768130912269355472458207818984045659242915299202783393444888886316129209690444801534067555373274285471098050284345768275708984379388765837105087551760272404179220484070260130423848984123420891784999930833374510064246408335304760194229149234370843041347818532553145446760503689076816956538474931730074912955624086515352456264005203796736461987329127371138970312808073275586643080160221521900215874088308087151430391115296474578781618123520388513670775318258078420175776515599932057241243859950600833313192587521907036116654584548033271934316221360383456159751925767842149674219732180632699417586668306525048550749366162544818630319514623358779834914055883641368035282951172861022683715669023793912938725123934282708194077433273516032;
G[477]<=2560'd1805858318579483045713064751585408066448987035408982917159919296859136304684080491199319840028884211477879684904936965410629053824698457672046460002455490771828150619974613129930207826667483937841491443815951129866127363063663545412608666566569821928635736537937780622311883129271692196759134108362436883463159456512173844725107659450858608079005740265757836914332449670325469891436971517070905648850610917734224650851319192168665248898630412698243516839105536130787388163133433573476694244574042723196576410667036292715412942124393647446949737017208463247622953976289183220383874029773177014767316834831289053281762083789570306801714864489694622840786445210029846334231132873311309543160930524801951663805065014852470136048015129823198847267693330523168705110639387152;
G[478]<=2560'd112866144911121476921100899625632082105588157381888021623574623197200442956829560524984210130458348608351248712090132552712238043179535558533917875399335871662421718065507316209705643625770185742532915013819940976433564500234704765882291728500020550758347958623217325741616103375150028570841505310007477673497964698261959530414947711685285596189574114939471200916108559784974455578569820721371883303329896325457033586972913269076510382460973800773498364929066777325073082646511761435584929387753210943856199219958447228804208457138161337743385079455450588125736176358226757901739853186090513075773173209048583176523712061455822838726734883102780071544996594068497660603192058808262103769048285575963471392551347918787674089642989113900106226041334102416047266078995507;
G[479]<=2560'd115539642779218408837167996247844404590773723290894636235768497392070131583542202839647541006867163721552951857953958893643008095599012651641011047574416935525645942940295295744116384358134284863418075126994816858464399063340182012047213379958540768928600247887661459645745791833523268686004309794539286451946497927392028946903612126949942034099983131999773666921537807691959767855179479041048218034668377844571240230257521067916534576385927718641842697195122054586044890930611030860817781199509136680249627942525625295591137684281082009408154434385329447583426483470264273005397812444036162345925851753017128247558075107790400808707708747607676396549657825012208205636679800160006009986624926029824784248751525041306101469124752377495244697508595496469801708650741370880;
B[0]<=2560'd173320084109970711720494289198052211650740438203027516077689659649862143493725683782486328302616943953466672165309524793619658785190347252447722591712549664159625675664650224604670752595972979134294131742828139792591649887812380222886897358289271213583401051430472000582462636123383600877940612198146546979821905779710513285561350675180051651882002889447609141013041912101708871061651780089771477575643289430630959965066442758212233198347520473616549188506370950799970806489509943039138652694681329579332798938950494503403453276383207339292204766616315269101009651104608690998598991291761310838010038342516524812817511154628610154992468807905459589352649764334914435793507328479851263766351633550541905524756866694157583001944015264900332254359673123139716386759774655573;
B[1]<=2560'd173320084109970711720494289198052211650740438203007828217177875666530843338786299118461633778026724839448259586163977539656354413907908213964490148101181445934151862392354204253629554080553630890129571280110120751109176624498780428731894153609352810938994883454262292413716286976227422579580223267292983168531976982262009542056952689291446846524601802087596315512668487646449718980882774078040283055851565184778880974058429175830081161258965791768064122521095177023208580855637293098233583236563675682095881999746880973331205250941743199289043565234841660968457654171980855351311515762492738399006709550869252110324185462090094765311427709923507836386986373625484119968675000180611314502743993937524583724482881573659973269545366706702497678056132091484619034724968781141;
B[2]<=2560'd173320084109970711720494289198052211650735795682407171289411421624922929077728256950965120755952274031775601325178452213485954039079880168231486770553465955453278718862492008995589414630454360645774817356161131583449474932157741287996027390474386105784278333121316187891408794705903950732980314517118121036057291448874232541403781139388079835184605789087491619504080161733859863532357154524871971910117849930088777697202017530638983907804121834482584329134662526543099210364997618357118855582254736038495194188933042289643589121927591183795542083562638676464093514437885312430341970199844406038112952840460704159887886649544704081989663656881525449554250888067250614732856801622284760058120225434035241400728495756031079825331007319967999795357905798206063195050273494357;
B[3]<=2560'd173320084109970711720494289198052211650656211002835011869433538234118271593113107203110399624717875276984167660117641981658420861943254809063404979882881242693314283248292132429047712111767050893106652674634980650474117971848043216521094905168188180986133147595269923345254520624375508412103470553586815142130958496040808489254870241819882632507776312309444070891030039269527238486301692773546468677102791248827615519713574356422605802866557634366316444247561671834854844890296827272799466283411776477581851734190946756324096269658424558715207691313622334440246628206856589988376742645525155792089973721877495182721364186911971271784386756103510241641031230858796735698778418217731635356110335296122644750827457913147003065721874409187974406066280219394099972230838834517;
B[4]<=2560'd173320084109970711720494289198052211650656211002835011869429223939992765489752419159223103002252843797652126980400914265990883224682294223179967314719456578196961536109441097761953329378960113936256086193727845082326131786225646044397342485572347097685261275307454163737304473711751891980430650747994681170034954417847249008275933726992489272405385393142227390853208460940386850133827199181951510316977884984601626006458513595637208028015573849342434615979866432820259245506730890772312872394732729117484136302715786981642202891521116921240321390101825901992325492692673821141374664240869798532536090861951577160167496322716539362061959337064076467535178518333086135893168599965311410348042184499095680169116387694867825414451068907694208265423747180637853237141730317381;
B[5]<=2560'd173320084109970711720494289198052211650740769724881738649047274633370102096933092344972614463431600781221786003800645802921504545159422768568658485746528330112212104840729118515608006659841608743032416260986514956518068030590018862647223707791966316094548498410768842675775119994034266537517599926764508266619312928627962384235186995929135615905803225444980895727814870670871964128251421568453632258509893393701286156577704030973396331625777782815842965930450755066620901783383476631227714187158642999226250972406609199340011374400334907226807448616558892554578132852063441376280846214977769698598889307954143151064443510130571841227007834220856427011207561279346698127615934242432294383087219680914113790084618931841710261583903512187969039016553031856488372616434111557;
B[6]<=2560'd173320084109970711720494289198052211650740769724901426510732546618839062381307311549436799747381490226331993948465845761319110480813439421894096896605589110748448856432001377352793002142209792041236928805570809311535958656398515000995343715810008576502257137890186512469790614845864897665141857229784330822344387321588813332643537535097542742235948686158125111669330044865983280650746124284191076491452311331083289897619896966700832443382714368896898364174133862735246990975705488500555983151501958246980296081795943929277975369382162635834547167854602139311585554579313197874656529716112098833405335907816070799598030439617905892525580589735383991658298412384496936849848859452346983495921844983167237157071773391785523996208078032841659479293388859974023196822683866453;
B[7]<=2560'd200401347252153635426821521885247869721168684686909202470915545420030226179911476063947707838601313171577192558036855014346861151705121824362324650299578309066475891496557140242854383205042922495500079908101005000229137475111622946096447128475205288646500323532461757842619763751295952853708316044682922920928578971607385535087434087391152370857723337680033841590464642214619933896652058646609428832201184886696116692034158221496681774354924911934694325479423584797603556665847627862606446373583148010277047248256514966229045279613073967703537985522208811329240538901555994107333470484515846792873546839985522376500318293824956429438725318876292665888986199298552505988028001528806509092085781252704353192760778512177900104894917030201800980763140312312817644337687254357;
B[8]<=2560'd173320523163957658884746577599613645753931379924037761644977758647394904611435758102979031047081113643955744970526108230722874397877171552395173175469590598179066490577743646517741445188837686920658097068018434467403745747426178892336773137925072715595714171724168554228829506716311758171314527635874337350260435484498514465978279559075426233528373074956611799594732535844501781504720875090614979419826618903074310216395468845237588463071468560998144272747349986269992328821555304130032444700837984300031680752069535950655067517887277110599031748292008695899986916839533465989180033792174200908564019896941325178941328662780789903192060113707329890573334783408419601982206749574491946948858938781889244349731682838390268069616336433510998228819107543858631419126305019221;
B[9]<=2560'd173320084109970711720494289198052211650740769724901426510732546618839062381307311549436799747381287369197856921960190968869342589853960468996549745257647175182812605221847920225120086933282129971310881270040290862643220720731232045558231021267842012749931876105117626966188938099456607146953504480516630532801697068692121286452835586527257368851217656097421761135853140502591054365709484603358108176978264287909661067843557948479185669453215881801198956977853021773563115248649440902682238765939674084465164389395132162708848565214101049643337864764995823434016041933102467353940372296990598213797876069688304822144932799382012192269585192701653401239752596166838710453527945662914086124605203597456821631768931878468899548513111176913082797912919750461042960710866654549;
B[10]<=2560'd200401347252153635426821521885247869721169014994417274403034507028032665878386578979036299707909850187292325576579854144088095148383967359378295581048705845345020116396494520092311992684952128268779878697509572184128714380834333098873617616820789485581787406969975574094829380780850163731481632821426221550781540234728866176364885117774020693518157155250627799935863444680889722529316302252011040369345106831943559928317468771741221897736148162085805726503691686407476202725598958298212163109158488243967775710811935184690120474701793256484874935746398112285828731052845016104821247477646799918944323542828139766561809651798047173646848922910923445935859988035807433090262174233827060262281078967440503965401488499700207491575036426067945156659432444767970969109761709397;
B[11]<=2560'd200401347252153635426821521885247869721168704116762618466922543161692555101516325990059681612906655388039179250673262689354350391700186230617424902563442013915189664886328208727662100819424090694873573566948189451941303108491035728651935490557701746080962366028684961361231017024306382145665947320297731495035625210506830878010687135294246527369427453814629473511886230471316678092424421235620052025129566710308516866054826350190020636806011704493174327419315393198538797433301204105997967741069896411356220885170917441371551852210927882162288480360859155144570348361610689384647271459347149881386518771804887855085066970364956823153510684290301844039060965905995906544861056318284607826571108071313341224580525069810375376716206976106380567470036769732680881065052951893;
B[12]<=2560'd200401373085164097894249451940124897460150689080841067542559951706738176126645573368964979591303422164224614814878818623624131201402926422899814125867230128279605714292471595236597868153782055486898765624547300972611825249927490994020014772343182299470570303397204055665180171799685388300303296509941765841867075022944509537605897220829853188992873727935520040869516640546485585121326153200561229423339757705188234384476124059038579316489566555701399011888652437726590208217613777283893516889909160942604417825332305441336793727814247142241413471164802365732755834625154478490254952683415684269657634627833617829870629907267268444825546435663845700508875931234713870616659888032580854697190953585138260278735246955350419305949919497211959459033202541560378851772333380949;
B[13]<=2560'd202094365258832363251073528361014799363143616950530887857110288807834663966091138083193597066946990191871578463267022968701832068015807109584884280919909739317578598090798183344688820761532645117981504946118831304575535865765233976099462256766640087730500785862484372482381606198218629498730480819586469417992399634158113796384370088049735889404553585954725441980409548607234524515605669842498505872079197717592827615456370554513439244794165134815328969083169202305034494514275910532259257488804659124671956930612520653832901373006188431788533006333095738248298312045499898731536465704984700666702551050595464870887807329356494027898675241202229631827224046445298535942486921714078144467745907948096002678197675596354504510213157621744343169298057797645827818805584549205;
B[14]<=2560'd202206763073185489371305093129486162870557601501800149222705535682517108448561107281864280745756175391680055396128989493757594580900534050338315346559970848544348667748023639540799726465670045502851751184267890664957525892199515257516551196527524899643056374357330464072109358746362111612116079281568014287298970225226495910831112803538401510240796379905528284836214272756241785561950754318754301115628830688535656941702780118507644969951352821072585269300747905058307050200430416981087466763599360700306012654244025436695546726799652338968806209974422161016611520818507566567590683054483459967131413526901759955292818654297882723488971613554108676575268607598513890057267651957856558482615455919054659263068564389337474576637727596306669980580677242540589239192255812949;
B[15]<=2560'd202206764687354559029997197130962491672407566980473444572532818844512543757589941212313017270308280688903010896167961861455860066168196782386318519844159453468990928372821614842128235820202063424453332628564988242106833280353273575125955231951034957041091047423064649636037489819407864984288700665761011030241178655906522399880758896445113519283485912337356680142647021200959432361478234279176217197911652821479967828530579189101715582891234618343706783669906296629692526049263884411045390412684446458937390019457212138601302172663487219647942811555030115324540461768602866420492476942125204539106445328101596324141736962351746238955673486633992727167869832901456245975778796434998900687795762319488312864730884235464262036682171329586686509173173992945168765130336720213;
B[16]<=2560'd202206737347365941685899685605957172591073776685444504584833210288214858210914066515337542372412565502417851350958559882283507699191588139828183333643568712490533874942258653860139393897698628630701863617765036357778007505205712561349224253019686227270713170333263154764354692534122155497107915922153194927075589296329947938063897534414962612527759516985239531099740793274062589290158540277996437897307332900539781529133963096408373374315964172837105364718230091690635386487893593162337836689837656876811104271575888619336454546060393740424837858163081121314801275025895667964519349456220239073751254520016963306873624449186740573647459512712735619987816720904065777229479042966275933579810097780032921236735007260332520191665879902731229744490149402395420941548571153749;
B[17]<=2560'd202206324120084109060721061228016999317482614145080895029048720817383419099532580320460992100368257515426994771787732191163848546878269069067793939406647649912808583472230369950638807110736820223783885035258614210731574134397846643013524491823641745824444964019898550020586401867898657289852834028882876176651059911305392514268775602752310347677272750727951413109185771561628975058205686896011844729681908953200559720923525228897217468680072575347946794771590436476601921887815756808243744268482383368638371215839922454017771394757267705305423255447276509009955532828056531932770761522517955862976943372123188452944568065662762067883798935914999194827388742563258352982724722291309495777831575032403106623284133352117950433154864380249576961012289071741894847335916459349;
B[18]<=2560'd202206351560958293258486829253114588948932027282526915976112534571305819353022757138089513017754034093741259564706164884778867412575659955293866130895869457351930922656246318575721110895216713829077962143564624404635498852409837494098054978440190736244286042557996443369338924625398384984569869729330489674239173271176522646432866741892358088985202647757932559934202085578838754395451275041778213624459564497273561746363141413671098419350851606650353048708027381340957057759640130847916057294620059215699304593902319918021900731090296526066067036559906073602319307829993319763627810157248838193244718200566278376384604870941332758534442272165186126955934511966195006730139200857082555259288020798676368239021752894463366630436765006350024286643359996807042552678455792981;
B[19]<=2560'd175118476681380480695633350018783887950929558524776234231894537431184475367025408469812162459021116732112717143580285115201097254154848005280688238998408248568423468841338721919793969202370220774733761781794183382357003400368443615747345358218398541415002977642448147077732231713832540602676411810443149010067134536949470612430438066018421386515043266520442073764958201940866943727558161088570910737346880461952890440172135653560172563418394921972207376528270247058555125971726133459232373049095511527692009481752472396303097634409812499401259470557914518048104058512393722064865843901428793838377174694046191855776601470545267135212469055366654915482407861601612175177247890701693148897339815065731130264824658820623814201281290944507971528269658646724500390381272520021;
B[20]<=2560'd202206764694053991205341683005793479875459109213430060727411215688381484612609884477987386441629398044502355649380423635405478018602645723838911606854817536817329337720388405143486161979589542139904129652882540907520770572637658056528524314642042892891435524465793640685370907487424294218667439723534803943268947631329664347493410101994414941626008864884574299818506554944998757993747670464676526470674161380259422748542126063957337412118369106094211525816821038706566314138864469801971237294042151526000276970526397135236039400994350840431269910851869011263352905363054412063272284714088710293490814023622819219093177618246858020805923398232478744037206505032737992562325449327666449942547360492531787923646444870511415478074741448799766363770693485727181275154091431253;
B[21]<=2560'd202206764694053991203873604789173079222985986987585854055255089095592199791430278830818902151814537576878727521313985029475803010124289924853140585069521477706288710074053131494632428631665105079220670715839372924464720931389669166952089435577870249618830015167341466263656367559991908467413600550835202379388925741608553279222086267917995224565795708690032966632344435296777811478555010461982353127372284575461676076385751144909496715695198209515606172352914423227734242663258934779392837351336377744442985256590022264139356160113228077715234549007822842547060712557925925477212434114282091678926063371122536541941105193425843957854089156766850959767397497154706288464289186133830817929213386251054309430639086785965217204489750712846956248562338787830556024092486882645;
B[22]<=2560'd202206764794965728113788340927746986965382194277223847735606686154726963563255220994637680592777097684954723693382267542578554674840752744378565152296970299621213076697571808874515081038200299721388278563663137476146874947485663393385114219548720171247574482142569800588378933873500812740211976226985512617187903710375853244335017827776961126508720211990463897735632064993783188647781265172240412747813132158850730427654488433852176465804226992112594936285154241850730623649240432388810211419579477238225779938276315040888029441610404090970245083238822309590635654704350162971763593888950654696306075679081211599926320235918414065265943940748175030656295548194024966569710666216905819798992186936125830428696820616239046504844924781348009259917091051955607843548014400853;
B[23]<=2560'd202206764794965734127042450885099919034897806209601908361349453718964527138527363265189991015946043781111017212354796297537408602033559673564186141583754985253857896408074285929575477353009722076008238936701384860367253412781098669415457664699690478265904892605798215559855025211420753152755611755628082349472137811925362943202852346180256662406524262717458043773939506482581346934047468536047903344918378679771571789138995596070934624406640735750757768988530810790233666094930716894138192658868384524814830822870103456850532737093536859659168927090711733833398542927331332716321739737361880205073231105952745620602865607005344533886878776446440130749050324879329112641417106140466549904084416160730281289247994535301181180683518392850707807324178164674988815093549323605;
B[24]<=2560'd202206764794965830340570577627524862807700386753436559830869444351888922235728940854246943591064520341447639407484166105069219431530596737258412150665335256816557608880501721021828903202387510441557485899136405817262231570953321771895396441720414081917989661528706580537535656163681205155116752504050138833743682147015053961855077979923660597533547544181638884091998165869819108385769310406394684260334803115093977926627886539109217493606946686852757798455024279994650879596241943477767998902669254053867672475793670607298689713119459177745169207425461480662379367042629441290941137361996982688743183589473246123318401541688344963275248531647822267966647235040492227713120546332116961558487916964539054526607400262859806800077443944528801702331321555504773540849112143189;
B[25]<=2560'd202206764794965830340570935957553853322601790277296203371776383871900720459248542889614029063245474688875311723092753928932254175627724874092570825664657921074681759501732290115082860000243993441314899111402999150496556188635124026097305460020028803532727478693206965746321796346844925332987136869101002265586296130548585475817388437254897696916794353549029135714401804179261043389002552546069574638987198511199598921257176545515434262717188868714260105344919822839657070608945028974326551732390730314830884211630905859682056255887339743098552116950054220018891911476380546698041359633642632381868468936806026801790459476912576652940948432033087352922194132975483131839226758415199107992724552270557490861174935824116083463743601360707331154236173683949920796649935164757;
B[26]<=2560'd202206764794965734128602666296483752766366803903774546222643735983062346572858974301194829319971448700548002944202058768914177453150338067526843225742171867010760695139250985796606159536333124743625967887506081590291271935802424719878624629321553472685386126957589277424149966746432682914826379078891143934143439778031849931356727965261192341556723641922084361525496492125164067753240125285073127034084115579500696540761645100115898184053640165585328784464815051609751244108515907473351336186574387875141115690563520253825054563716691427445518434562208130556235162728648198877875361861649334503627788448173918299239648563382259346077991975820128398327655253884374972611176627506818134981335603257297916130770428114335539203580184694523270810904994328964617988365379523925;
B[27]<=2560'd202206764794965830340576670731060913570883865082425131680936667570128431678221175530117082635184321444780559148209091299416894870318126751443907622535346349964817798734555331478869865150276534151446570702692783486264305194151045933944099535702226510203383096796437737327804431472149728330472144097131353790859964460315548570611650782519219413007089245395744156433699349077555362081459978430349115773779527857492892782307206290949670138646331355281108117219912587955770384592638408496799553671064692727958010609436615500598751889366416468500196983956401558096516500101125188143473007404457973989104062070782812452367217137384591555664417254131963385356885616686276129843240083483056741094870207726725196971270209981276738586552686648779818022213005794160374977727084975445;
B[28]<=2560'd202206764794965830340576670731060913592530898012365232526868639179977409166464439254870778110385053655797597082796584845005721252703445465551153204053571054089714574508283436158879835631019559602425181104980860615405224781934325348713103867546291861009811291322806813114855110943273492806527181764764905434357920709418518517769558304326401953102116859643409362578452588026595706710942032734249723449001175896057252967822103421969666749045574487650026941014798927657020532599165085098748110987687867481494969022877689796183309514247941313560394538030041156742851246474179770973639329785808174482890467058475752895118185395573392808231972880972120342541495303342000159059480876993391254933349839636810786122285437943644144434577009684200582372923805503081230418330535679317;
B[29]<=2560'd202206764794965830340576670731060913592530898012365232526873223117485759416612622059346957163770798462417627511728926167378575235605039908410909435594837030679680986503069922038905299165546631543222101430470105585024950752339979648966796385251896490791037316745935241842490651940632084298690969182316416078264323164128548019720021715262012125931187434062114871188753234892551914103078541358103546074968225734236864893725398763788765315613439081033969371865917055886317976096728497421095516406277859829814961429258650433347458759985973617785837061480923673498490389396799569230088741626687341659444501643934643458636416918759444514994834027042873021619311522247676210550226909769310470175123349851565439961475116151363684044197666582997357209151332647594557944750551684437;
B[30]<=2560'd202206764794965830340576670731060913592530898007325139935443594837432993897933044017075550681153738200387221787310719327124664086131399251798035867033545295956260494446326997196117426185885165705508143178075239182915128762006991837379391038493029871809979577489362686211634537428642843000349930161369367177879480807798087603210784546718074296865267501992341836029346632952365900241824905118126348511171821763304799846863398027741420544974128410004060098165479100269918056024530108742621364446193330022942513456422985273224008790725666692880762712706251524814083057952415116830229772829791947419692477775454901458593935128456877189484404712797446220118323095897850467188381902405401703784264351199286480321734134813965198742092174661365016470492814146265905209088803165525;
B[31]<=2560'd202206764794965830340576670725591896054771962012341924175949154301503570762962878126581705134155171928672319628189072367984495784412902991321456192369254596988583303997151455282670754393415962740980741037093507627515194375265405715629119149619081126933992012454429566675914136784868623683933898878564751620546530199142432362173094383893560279321979098737451197976410850770553472775251910618231413291801315393978908397388633883256414265374682598855871562385904556441652726399479385908630208439989405720441913928630974519077991888697202802762228340581734348657870651058656452717536910705317476914416353845892746584151485677628348141032842758520247594028341001189776050297759876293938563009737646402560951945718599410091148084601906348502872726078786843762935389831260624213;
B[32]<=2560'd202213789659151069214043671894458574850299041947223890957517075325885562316819695036295687403170701507946964831661644084765093600632223112209280227071536599368361606593020745126396409256131875673116298634078449586968116131091854380126297541181744894425584005961812060909182442945051012356216173133745064654503290772782761131551111630007125715798879559217626349418720312975978694303552364830223540226375051660545646430762588009038301138116014239842354612581144271439274220886179249564387558826081831805300574573828097467740571700953521940627962754089094834528454696441610047269878608928985971761931539671115560358045147851073939454698939413018137894930655570304365546149288705804023426174116947507037947635395526980159855296356602101728665142828668168073249983076133852501;
B[33]<=2560'd202206764794965830340576670731060913592530898012384997294337231972585323167483170307173062653365130216640577863230090429368438819591775249374909354139588700211729936549757900244436497870145546489416791395229750207099093101607983013756853022684515691154923069711448390126393938191839079101974517431611164904761606226660249537051436741065746603185263455081545838839180461095947106680490904381235921169231038267479522230580720507292987147771273382453206752173875501131326987928067372043611795385183705076781400697555543292861697869560650026492294325626321032391845269803662903391956950458900243424239623594534727015273205949978019735514774608120018018459647275290520215774056869082672609390767261323664247481656738713992716314396612377916400341039312378422184937554577806677;
B[34]<=2560'd230980606883535186778549355461206300292360907320963352522779985782207697803711283945714893626865679090884241643704347673776871908449511536959378316409430675073204144070526218839236068166454630892323787798856508054924246209913373666664508248070627767323666257530698571102257008282442187299625587086000147548714774040348043654152591978924069620623464772442745826323482850423462687549629219351507105217588569223289079479164259260357734838791930474032603988849279996390424478781149642166701438133873160990203820573824573409984687262481572543466301426045860839338029623067988978065616934535306088834234155097795905826704519525599002763896581219127013066918419361988410989756936029662133393706471540871869098075197709162859141976806307455926982653601392339528675591251134076245;
B[35]<=2560'd202206764801271178268930936762316680501913123149753827190975487463661199777358925810981294323799646496647821245805502336102308197098403639573037052433858174412324867419580473989761035607089508834678848799142084440366795484425247254948827342769353384276185530873746801658068980247358919524210748045343758908533140365148495496781036966449969948682953213311007586069015325565796775282659732185660677278706080827908704461756475339391176021313086760228806741587417008084638916283016188075463495042335019682157423707604090422032158811604674481441818377803280662080156916505608134055253266636923806462669988664126248211993916841268074257229460668187113722401259357288382057907262895418997781618551746211898712117243729262951286793220142526499899246564529312396745872021118080341;
B[36]<=2560'd202206764801271178268930936762316680501913124440036060349139015084950453745997695516994920340135407991105864857619787931895133404820962655617909399275944743160680922711826708740477261371339877461570474185886358370851010826408937795610794607904852132139239203087262847538553786868334227603944547585616971647952986107148239270808518428800636215221264455637775159704106527158459570205662549371784565474165512427778339073049455312968097079711450936914370204996981357390469665250345335503905345841466939390146343014626380696976332863074786593525553852529775006503473214588459132960444999183640317612705053755290879495441234917666080351850697480410392377392018697227101672907122626545364416306726692067097928069497723791856096873858947001493012707714931907480223917370068260181;
B[37]<=2560'd202213789658756984968613285156043859243580661198566360044121930020105273351239453361281613503872080762900394166572975866505964548482994795307459892105285897403083648388856164074261385752847214328718383534943309802127548153957709790755618343411103936613437511085524607493711202915571749267030161493495485747661818255283211955740794981478503597159908027846298782984025777353096923582212786859424668568333626706147032013930420727033378827701895238485416859337754686093826020198055328497491711486573695301462739442985238411219942746475508334506421128850078033152533258691371602090376375661631215725424820291819527572812130848981865034147882361868745772003457379375096549308594292888399398950391101934025570724823345662918211928203736409084186730615823970381730078981734356309;
B[38]<=2560'd231093443758180607991387474662494864812347729789283720307827626785656952178778992540103747384500298034675207520620816370866966858999890350640112811467236123516148452444022396529162378014451296422495308177140400693430007099062276702956735145515524177210851922739187141128428738002206390329125989313577833723460812864528269487012111160929920466227685506179728841102132281619404420106611342189476832716936683914662261136013996087633744737866010210386574151254313356318983795201497818962731922767176749275182849138740030742823516865435658504951399615892564393754344961989485418892373567456907864458645098971789329667222419604447934912279533512117232612767076321934265703365976252611311379753527145964038203909698679586148087195372319371181228736026333150833352944706666190165;
B[39]<=2560'd231086420609444089875711220739080518513263554924192661786838362990022805210938542442883197913807466674669632995953742548453919897834784732358561777578725155105267020345760119178318534472653622079522565098902111343619379540862944517161547056878624938733232330682589276390869127292863228153753553442364961974554647811975303619424732832155405655520610031648207321802112549235388675463052008983403949036751443058025307693060812957456678600393902773519766517432057715427538695761694794067099819797664480771595173423030990477410602403066234032415431520524705519013522479434266152548266888435457432765541365287298656382578546109834584079020632457070972799410049733963710784097236382323928263370557239694232462930802950514166497105806834415582887070876889268832268332650988918101;
B[40]<=2560'd230980632710240301317623020884896050788247970985722704117576476345944950044006658452649678557118560925530074299881074770088224814408817728593142648615593306364671731292765319779960336735003549097743862334973791878877948147300147231962332087808699099079922151871899606887198971237597241766381473562937172019726091161336332043772026790214325077382662751667608457016639285689497350086495637152505100349263924966207066179277861515420892382009250448056775697601503553684278090500262019160760587842937107604521581722863416469821055166964105823549997350229652997475278187776483116575653333588601006740227009043524256343504742951545457159856124876155318428501119749786167707308693565705902260588780532608505093013990530266459659637868202842913848355373898758821045194294975354197;
B[41]<=2560'd230980632710240301317623019484827561121960356270018311578662001248674074771633495217158703861449486411051716828058005454651590415676803020329043411778230256026068265646507529730496748562278470326092286013867114174379936069722939642430754501807280803335562555366453765312663308672763136632703238049617450685343334734089351234651716435292801584907022144251524680328723225547325170777627695064435851392292240077877511243273957793508396383418120173616470254918079630814309690179341147172122209228335386172453396963778756397315479674206941732991864170614273571638759088264264384599608931811933657856485159804129596059900970625083362193911975153262059963391419535592711013960125967902913815143824213484312528422232336406624951309024758903806647700118321023588865092669414921557;
B[42]<=2560'd230980632710240301317623019484827561121960356270018311578662001248690213474753987975259448740392708518328148513088837213823943627622563242392116261644552789163810261487488399961961023629096190375498949001620633265131129996540372657649903920789560426818129757043996466597533096515216931769532946169620575392726961671227914318807427582981704914807803606791241767852633910425123912004083571060279449481313494260243094160539104483774929076915417290214438869782291161699920479971712632912160641953186242298587316859246173435423224555463257868075101117198653446272802338565607541220791426890841855702876759522643748462558597805950669962638226727382401709956262843175133819348856033191731506849251416718618614742312083936495328274618395721828657245554670758375077364349430748501;
B[43]<=2560'd230980632710240301317623019484827561121960356270018311578662001248690146769683720453359121623535762570994545777749603774745696489670451793714542233074466321864946067722059195346867119807886347995008639007124777726346459113578995306720582582115158593309870308374307006506949116181517266615481418322403722724249745969183712000563364965996902692255808772122941606041395884672540070335658322667579383855163258224579554683556005543438797729538801847470369273956009950364717525989435600141153318775725433112624890342516081704579824011615859500479518872252318864798367390336429516793418685646742621458672538583163998848635857365783821035060740896640598623527728776819519511042044622194448773431508618081110179687228451164694048548081292522083113176975993261808482116289223284053;
B[44]<=2560'd230980632710240301317623019484827561121960356270037999440347273234143035056007480543284574342029287443019963185656516617056429547182668116251109140540236566212629350042480703419611187790602650981444967870301378774377207752845990956028513650860992018988266716279780253780830475805824333249913478216518217823280258420787835889306088911403710960148891947901624716630727218995522604672980881192624464283454414131219141326380358253020795737347060975301263418128075498091728625384224734518082124860708286938287135488219114325864928763607124751434361184744033228568458240648112268109845110681468197424188348481876780860409707513951075139784741207083071518315739599442749742845744474285995979711795275386468897429520311233679407442273906461639972390464731850360279050003923948885;
B[45]<=2560'd230980632710240301317623019484827561121965330312492806556453423110115847462127980444132733763696222179599501004596644278598577028957482352110931636662271349589227513989410027895197517933609779605855678601099885232242353372253364289570531350375154051323408647353195843573588892011589698395056905990419364140532869061652728674129421484774748901868656325401622191296296765934421877802273420780113309147324957872225556060712607900057827809511956597927005161158665666693205145285011169722598719963628622598465679271862868227508940635864242777815737655094648476924426511265417274596858741686218755069953119739697911929252896933060651471367056391724285309725159911999871415926021725353732732234202744980873929468969972427539788805025597208223587889512425359280864975577773593941;
B[46]<=2560'd230980632710240301317623019484827561121965660700938835986305444039093455807109537437885590747866579962162314825146821041641674505677533985680697217271022959768652509860879536415161015532482302750315562330487548065557828443363543324846092413848003406914705825907711566482091675490910804232076195023598757137261234857991267307215422600797731177226789551140029880191588511045810798646583713217883850457446887953966224549649420439107868549445413373474661385999657222268057076400996077034166229018022522345851609777725599310800701280040321789602336945353214678377732068368577771770444510533554066651537916047419077215487575926974023281994782874470863022585005072024450514749811323484688914622561576681478389725226000648475004023599918560269217480368029558864239760306129425749;
B[47]<=2560'd202206764794965830340576670731060913592530898017444778048969537987518775954198568010997369232298517219129125398362372040699510355613824157315323684431830756980173069550102410701758112125518452707074888861589083841454384496379692798126584658267710178255934486994261553582137075283732759088694268521159480133645728574117466279527669143093731681854619862241472110640869980080815547627551025687672730570796558651974695413432585215913781087848957429450802956254472211023799962844887274872182401761057986875284894342821708492379002884956240866123357756095204702571287153553405511927669739591049845499812711416152270734907626887616124234894202979859555631810871344606934341698231870515756323207490528041751611315230833784325845125113578357874229339861191224463619830845191574869;
B[48]<=2560'd202206764794965830340576670731060913592530898012385074785479413626993933146218396321194082688850437600159446028679498895092464519855123157665711361162644968895105445251082620276088619585228094307185425194836824922966512466252160153216188918966386296654840379422636668713890354214967188512825363196894544096548915105099455897490781808721958369883962842386188108965089803171645015133494468806291513113561391204460890729449936907577730025338922383983209062073117158699893512110248335752183044048786815023316681391378454242359677815384104758447955781616618131810987291511861688609214512217465870746890208027131165394850635969739932057159641607314299577423680272322555729993028704921773163122812439375631510322866249457327938450800617094820076529757337639202572805405865760085;
B[49]<=2560'd202206764801271178268930936762316680501913124440036142363115609127410755432806889857121526695194547413906578374319053867981428627721656597191257775938024876113785604589550235934005740269950326636327314670623364822917491556992716089047571980248684903817494900789977207132821474356278465096413115667744287253610766683817828996404147919284040483711481526916355412525342573626879967154656140822034710545079891761011609181204330524044316675684887065220371966973206162078050597367995118230933084172973692718725445201488866245882635873157549753972196668473462120073959375930951024619074898693220411097598976683054588190780723024487638834454733378316222376957956155740866954953858166377325738855623212890844128696765679908243315541913117954048042121075924133659729616311575467349;
B[50]<=2560'd229288027943454101998747420915437413802551520895326069903936811990357442384865484037152244408839607673113144789934235207007144393645427337639002946648870077974099110006020047318177330981258249790651309000920836558330084584380546307970500945797686901646094806059863782516055469868486117829841571202518779462662109491113194285352646588351057988702303774222377749512776327184201129234286914906740559998307227660611505983979670900480851775213516951581796893338932008905202875226035757601703244666905912811771481796916630693398546972045898374450772817596011378221415318101947841539868729567904683886787400649029320038878602853300129447286552286831495776137510369104825307112309444810992782551535750510391697329698022640392593963979762541840835657279053832898117577036990338389;
B[51]<=2560'd230980606990727737164129953287392767745106125707382919191740582820729121618546105376986743069132494567031022494040271328051426868643440665413682785767594642028286979060289820475927926609151319568806564074670805416347648395654785027719189655560240088649122411341944172081364967152423849030692340671426105004079520416642522587671402925682320577682791435371138035481832020690240695163022980285497964255572911316504242833454190973344630190971585327475347740477125614125565845705895939041623069831504262671716323456075709446425573687138536339747649681104306713116245718679254253521212852297823648681441784750016499081095553988425907551883291247157284422701779767692215517694925425353177520667179313477852337987659190980764914394905587656276441621565505854602049877022111782229;
B[52]<=2560'd230980606984422389235775687256137000835723899279751539493465591981346537249068140399313399381580108569425400925073263112000330453995111805915179495076087088856269624787971414221836502329228877153346054272695624083436098237569305586385910496473501135802503112147005526969601598939085710536659573795437487835832629956626727472224327728586365109396423043757442642108031959174051914568214208290681468255590221778715019273559329257087066094060933592662246142599537019577909192500849789341470005522524881929245530661896586007522725448519434464568656391707817821519614285815804036579591626012978468304842851170484014072070191586256977045622200989597401953172902246368587601465635729777233445413068332603169343701282680387019475229661686739638575442342967927869844151956548179285;
B[53]<=2560'd230980606883536822382107430756044730285608276437334530914845942572104947793965555610226676041627655062009812826874019089776404817108810093283421527553156630463492160591405456178143686066747700312124510584964101614082191253497677076411625453396904388377204674715594786287726219795607507102439706146097591198228262945902747582427228061225393339171862063103047959460478605111157563427685006649006116885776558365399739051894928374336664218065669167935420109128653329514022700346423603621567629942823746611159673407828639179793211159994631326825697085636472771373949945788881087180581782737354918085050766181989739500926804082712365995943574548276566322970662639180983452735911030596441488519558963985383804074674471166032894693421321545199585361688338825494635347784278299989;
B[54]<=2560'd202206764801271178268930936762316680501913124440036142061524895140989611232867655298730268878461102922901801102325947517107756277168514450111170827601597863755433876773673563346799430448234039377166300988894633329498904782732620811765099220952143312264896645207508129481721297482830160081064188700325344500146935530448100279020107757157443421640191213654899850410233183720269370271140749671829842967914405703844911698375694380524034678268417760772442819739736232013889157772255054436752868422555627658168538799949568453758449359159981264111149628959793400976851807620938947608192318656828898876524019318673762300181620292199572868252490524975109001149679091479447832869131037153021382190525849711541620067463777388853579707358834303919157088917696335837913540454258136405;
B[55]<=2560'd202213376437780500295278178275284528109581876271628051508310261159263380567411882798633883634330854010958532646856250895254075285986904922440539630553314258195116651566365310300407500279195864767771949733965019921459950482687030373295862292084019017086862764536429122901483966736348157771955918210308420871015641964114698061784970747544162252813305969409959938157399827956249625253882687357494088592225505378331752660411076643004780042525667553887472754064812857772716236175229541230001423100944119491264455899150551021219003482919664541533925877237538542383422564907210164626477515796533866906624660026534752067526916192243448968986955091146323152806380809062900263893621833851380776108241251507749472665088800443391394152998815423015553246487877607448778966279069717845;
B[56]<=2560'd202319601675916605894340440841684455983341094859630466043351556822502660137891323271203431391660550918490901504971255263809120320389377304575640501143006740314362209937992572785449357437256268099496464309137222316035416244929452282277449485917868749046613997580887508311100291333932280128355543825544643854550159614324454283876331259988928849641945766401472536126279496353212503908414659084576074658938301919562360173081909369830792865695495546059030793983262889791558216840170918772522722512573613163294543382854441694864359098361313050784754935568383511436914682158309363431959569833705080159573521032971094827879647718731964117432480542613332209624861043323112482127331731514884579153693199458797271720517459192998180707415152453796937785717948317480513518936738059605;
B[57]<=2560'd230980608598591464907716166534432588571372568316589224563879358805705756541983582606164723057758177837458478456764092297487094574500051614640926987511686537004044512989973759103444137839167146439138454419476105596589200456023699641851767175788910084086057955772472534487338548046905876163721882353199572253067878455972815390186586308075703466129037823282900873231784392315245881267283950061031457173787061911801578802095817445921140105808109195445425474106612264509516690205785143726371594757561297739985099356866815911723160085273398519659820599060205021420280334853718958436036642449274330359741740195026607601456164839796840910022568517753298743467456180921892131128746340690863054572671972477106532427538765025382399942186429775076639456901539288613749878357103039829;
B[58]<=2560'd230980608598591458894467791257613329637573864758405146680090501810612808658750375894476632701453344129012727127574455216952898108306121757566607261681325372929265171712312067310352764578748399346222088057839052100487415785001381005381072916230023580905598120231264770762734598173727835411881492228867589669498346142183135346256075760644598696362785567183085029018343634561576793816069259515855597241024226468217470026755904647254870431050768697739466641518461112453604825477799114667848786540996882030182178730062532695131632187702908479393817371560785427056596299295860733589770327579283367573239346076461457331723493300408109418262548740077245469434095785099030135027017296472815768830644060448721573153329477295344097567642072939128642339654517410319128450770696229973;
B[59]<=2560'd230980608598615992949306998896810096738172516598553797306828942122360662742263172349441006147291038512609108879952437725225553654060177019037811341771548266207249367615189612786410701795448121080464254096625020955783441251022747261782061618968041778872697293466464501989287474948228441983844644008227048856708373734187731207784735787873766350232194676168384738152415871890209986639183115611159026655664559242736280371254399445690828784161071215529187041177580273269840220720429496716864369602788851673534200093712535388837265680115044335910419286191873295903498155575217705294638089957803234272316500830397483905952734852062895394306999905933805822380723724701071926687702760252676483522794220896217302419345871595097865450257837461599814587936043493470027846211060716885;
B[60]<=2560'd231093445479959306944437454890577626546909842460847252666772871579134047783225627660134201728198309388593888739323707678532131948851220249503961741020036471198354127141592256919453495707627869552096088678368541453349613294546872686050646349823008846421523158881523319897491106015467194279998769668150386756356454054213303272406635839586842242742222881575757622257678158593789154659440678925785059501408837493572396844448099719152934567996252980967573809687304052185869443839535321488005657717853160182693033806969755907844829366289134717441819283213202538654737030402366400709967218827953634189236283361384649561104527434737753912379623539364789612383241648944023671633785738905682237504714582414086930633637210294150460529210989317126990965575677856401698269068300473685;
B[61]<=2560'd204012182236866186518414106772331384000448770185091973254420410939643722216880615351593929768923123632673950781154866876698012645637243405531424017814605470569879817117507928966565010121666996387261355905440656624401988027058958463967356679505639532558054139212143112508916433180380186844930086966643836222856030361562614172621301587163987916842898044624665022461962125144534811841139298512378397026244831831671134276903638260328858524821697422462876711848017278231427712218457374071660244034307237624236076999997599842155232024133851123850228439759047946649827286437939417935133561992308832274036408358415958470230247552442969272713781546270525774241090321557352552782814816476065315677954421426407114523124325684832071052589856109503397961440545605003010606148974105940;
B[62]<=2560'd231093445479934677076941517742998995419104503847914017321446981694205820477650025680859945715074566725052583833341905823496657995274662374502075169198101967055786404443137015169203096377248720563503843655491664574784751706499802274760608973023436184716959438822507306986054060622532506193391189673642489142820460021350663893412463525729557905077694038777752281406533350878347211222358771272023781452575185101430749076318275817240251631207838408166050699296554710923858488205896732216738202014365639733290420717330368259368586763157410240566329534540282202624051516374014440083447808833945375638709931095072169102389036577843106701866049352071199991372298309793859975204216934423045559636887453201127543548817264019027467583404194473217974930751332181403187542240338990421;
B[63]<=2560'd231086394782738975336637556715459257683664107265420008571446264668341044791656985341242791861694071283765550980591474089182737416324035678242718398831105017845825659662326318637629873413218346406582462915703363112918236593694625571497941223235518502469555773165685869166869206619951520573359603415953158808530857724396262418056813440393329349940743919186237451472140702350151067180101650603570315153423327619338663638995010591757819806498007667438665122247233302690358308331015159477730075872245446733085262158719758849748924590011540004185494498906090640157019338077008969281547683085746598477326690104214080358464834027097904367786646876514247094861297585370946457660957394601144865674592677778154093000709923537802102405835374449023918369038850437140728726428975453525;
B[64]<=2560'd202312550979114982409793762949670346862078659531243200430921791033906496229995249703646306373799402472056572873820239422886419341773191574560447245661040154152568805839708130314232835962448878506965880733900069299259403913087631297329224514593736792964385024903803085136968182644899128093530119159141281339531746491851511199716100732820037282076065574030598096191572169461253687809877344215643777775979088212099903931366103365814168104517241554900772391387862742637924698939572768494635509663030497076962216556885572202978205974782945508524836395939638581500983352162688640009853301776630629920578712798055356454470099986160213027938742801022966259774802274183602886435843355014022198800367740431144125817901248966838357335116224549121307346229459575362063081902219547989;
B[65]<=2560'd202206764794965830340576670731060913592530898012384997595854637721978910296941106314967173762525340324870452338729731005851848696378710119314738700498663353194420763755957829354920473500845357271366154682848518692273244535802196999585553984543803702689044481288420423668962980405286542599862742370402059525254979351202934188869796435053257293442151122831462123712977375429159092276509685997472687449915095849869803913347713017206827275984061819819422688790816791222886127849494938357616492025010311816444311183107886012597023690407944484818143768914138668349655708274136632272139822098257574017248699484868195482963575306638382109748629689166445861891961634253960214333221720176514154647483055410017403226730659962274880519489738145494045281675839165924219030103802598741;
B[66]<=2560'd202206764794965830340576670731060913592530898012384997595854637721978906372155741008905860611891326562185876198699608708893977439210593341345117282028249267554743787855396228451864840130608996421622380648411853673506974561355258387314437386796042842784646910007145879514333480831891088593447677591476827562773786298821183714662891788503947480800499719863354982905790351143572752288230907561961468034155994710153872022485910901519943928120792197753114171035384132527418474661296414131202382469058572679203834952894975000242403093792075411235454725853822607717366889941599497002694274518684448964298399505223893161353863197890821180577404280575734462758741461544379182629484204048884282936058814882682712231455030641042551216038944386057884392714193178287294282674145154133;
B[67]<=2560'd202206764794965830340576670731060913592530898012384997595854637721994978370146327264807275263785789640441805224141483895259364224667125479240919553429889596500854043831630903898058014500483087465359994464079494799123449145754203587058856778721717528106490591896969257097751597986351792216023905669235869634909191014536355128191034422706999549381085235777639063579396600435793526750460935793008934041034163463173727802532746101457428076471497764874080064372413802136431124659725209229656518921844793226189709037447123640689930103794894193383470396976252255250225994027039901911008720432963701590587492960290369894060192363917999789837187130390437449614612911701662666139095107901086818393072843891533771154934143261418081039639305500718781153495523934780546351083017295189;
B[68]<=2560'd202206764794965830340576670731060913592530898012384997595854637721979910626734559901916279644091768637006198086995792373741421417444834333590283242240725929010682485707843218093741606074095455134455834250108112431571276795433196389451551542865660011810048577006888513478972618460192087410254651286866499520415345747683070436986325815631224115299327633773222715677252048549151480270681934627124026147684010295447767378364623413688853520327323954264330487904453822478071501088726142347759281712088924835997087022669742330559512689011218864776631288688052169388783977415492522060558094638696551581177665432432990065098805279417580655208115042292073287839765138601942382285696096566210705648501972447646136306739118081448280548960975363373656627476205102250570652415110174037;
B[69]<=2560'd202206764895851397194244927231153184142646520854802078555218860891441421341334396618649488370822874438669164793392295005024788699370720554325683942788056978349820898136096055716029589901109407724792682618737973007778258695475638297631781236902360225673631772890986781566749070310913774367951500227892492026418447712714863415587953842367487951713883002941209674326162426012112336770794160600681505817381145028733017622124517719463325107104900218448353787998814067730812180959792665001536290543111719315520639718526225255638059048865106802744409288084237116512908064287137068958746193843317991726576404290815791047676923477444735512904311977295459694074749877058302223690979827277953906159562699873030030318402652062998738152657852079306164077413970190119836239975405671764;
B[70]<=2560'd202206764794965830340576670731060913592530898012384997595854655627985802619839562260935171341937229663991544496816260050654688739696126329011252236061622842553891107807120563987035457370746537322086197541545674998088329315751658519690720169920461139072660513618847236033674611231983213799198559915990582278633219682450794053877317242910263147657258320881032670298445864693372260621815908274539177717216558960634352402259213661402570682625252127326508261931594390887107056810059426581977759598476405470150506877860161991123482887182208084053261186866269875324370252302925299754159111155873939775924046838793167587359885347579126642189123012005984759897962585518959637852105197645414247363877812079470453120774771641160644629892026797541025426131717357219150090924396467541;
B[71]<=2560'd202206764794965830364065922196985988822741049198159154150092756144458000176596689666025015955148226635962754718559531934074121838469615693724613709349946388133269805948914810095611413099700030295411951985447935667863957786137383061178307164448082756101720654355074327705859773764625005211181331062864893138736144302005402489077377673485995315752044344990124055283749048976708662501700488355894455378796547503265454981366808997444817294428274440790498591738641286125299475377321873513953105664700722213159898817497734606824844311483359035931637113970793679303304304989650756302421727853149045926736996000397057301022818005199560721035180701003201486994558239583041082794047606442733826038309171067878397988741439555967102743571471083523119700959603928308922468989341619285;
B[72]<=2560'd202206766409134900000736852949157559596268997940169177730321516789285017078057356772879547744522999664338424041156566181750606315378563203174890135855589316169502623942354776470110557124439747029231032841946615177544935417384247159765547409622337786650578184126367666539912491769735608097504232100205440743150441862074065548227775391942665464365841113446420157516581802760573051685759832471599547276263106533858876300647474228150499392908848993791175775679994839592550346756285887203807730699519379283970554984816623452413314380387289288607803315740552518416688847021896505623653061878437530456183780472819338737104181157104294194804765371746382673475033970568552560206282173480510610490566748291532379564063616768736198723248386844127489202545208549812565526705075475797;
B[73]<=2560'd202206764794965830340576670731060913592530898012384997595854637722252134263798912229243451348782273007743352953949952991597205927122738239190780443209914631415371520663885026512818232384731214596912268356844203549601454104840493760690142578705903248975877343219110476383002958128669601217002459327580007554399044847771281909070089652299697884454628119785972284259578382557836844342040921091388330722556529798787014454804556271201582174875708705522073684966124262403566493350903812681116911776731924661709419942092954143496294487745717783764357872891669693965811161776374288637520617616413437409971077681219582099438317025802338249831226849959976730222064280681651633315395058937261049830841197146670673253437050773412786224699320063787817922015403448022980335239509136725;
B[74]<=2560'd202206764794965830340576670731059578383171093584651847395594461016702750544318898403920394065847544434288252144454275005407125911815455186777218800621312801129766795969743310009447397634297796867485895892818419375071845854967012223765671899916582766410164768484734314187881519494650861768808326838641137598777886929124463577911353788133778832283280959450938844854203482353225516980038940154238716764874485921483180919939548630507859024069835907232662419539447884070238099071035387326228097584063533560971544088963008695329515476211271280777846068513308971286621392006261190973929586776212157813027546345060256763047303693671605665555766465466239388783239423337533759884126582309214274437009512440930057748235867568020414801750057738473106893119214751100561510581784630596;
B[75]<=2560'd202206764794965830340576670731060913592530898012384997595854637726367632784312820614950777208689931040768098431370730021813517141137678407427129257416701015567049489594560314940602195357008769499505688877666399956781602239726190182177724978960596776824598294948252383684907746354212328595357336455182983873143707088064259857605198450558665627848730433390436327567374460092388128237625265223048444478623758941202614978535555641397423468272004083276940870778990644566775007826090478788447089352910144511920595850429039890984216489929113870951459911810092491179739589854984821419298934750413541833847079371595589980127817942838661301594038881033954203541958700459720755398789524925332576536753635601669378648313298039524096453534597381573691279433019325533477657349310469461;
B[76]<=2560'd202206764794965830340576670731060913592530896722121294189869816004423232044226069424106195617983435662061550161763143224220827508807754742451471207263673630967657511052127502717626796142721339568677861510901601941809424738919244215865033681322414622243796338765533129999687442865160692289347387842588433199742035457240041980762816154590583170140660463985901787974581616238352054931359944581626323940686630580454730668961101929834655398476529122324784175282637856068708877559381727356790644793750085146586132428366260611431666210941841185573868059489156826896656051896249776399252019108589630159593333612458511118347641263833507561406335862834320951567264358328669647474315456124513304864273859772766176366885811598056994077840161452197155063800169132604223336334744704341;
B[77]<=2560'd202206764794965830342044748947681230794419032385598017474259849268568588290595947563929945307087012941798044703134536723688660720720887558901316893826781357646244489635702713455919197634080780522910084411134053481527985451890952343449652388959139695229065746375247667097025836591603913665993428990325485473301763653901832884671892564221049360743342655774174410482806586224459936749210300766953967252432341982528624108443943227722902716360803373251413130453902095711942768828798212504335868939053147034196353569591573005517599091846530515573117472912411870319969513899035793240441133506283496926039152885678328856093673457609581451380135926747675575963568725171856085880505857580230603114386540954582973812758599783297320133345780554178825590595065010242638931325655274837;
B[78]<=2560'd202206764794965830340576670731060913592530898012384997595854638845491934014285742993883823598941110873652919928175889228139690395345165876462492024844954849986599374493841992265334069287337641133051493811589642337837488755321775295725507969046164759339282438185862760930885139218360625372958346227774978389735729147261443966173478367165206352495444017793718061975529970144491554136660377242291315037044483523859445628983865152080628884787168401090323344814725598233093079568597397364443663921272995621222586239386449578922663679415764646920379508680826070604682951303914085626316855698335697222106686920684515229214046899065688121389534585439422793776153635214772666821943198867399086501183007182616961789608991031893970823791126463864578321356398652415198694072540026197;
B[79]<=2560'd202206764794965830340576670731060913592530898012384997595854637726367633045837232290147021387774268478005619948431922039417856361272436659775403293167635104963370749095715089232749949601042670545470553793861211591909180831063764301770363174378328029794476302067125338780190126096658332790785092952159977162103525012660397794746800403517890843573627633552327613606788925337421748485828940771501141979147225622737574570032665871472173814141648032508154441370369793763241772673963387021908181123986288725752921546609648964172839105539370702430174295708514558470030138135284525441455256740173660959707910904553133673770352528121964540459363378668751307529800725512142890901247581569469814969846881657173290236061368776194931830409274805481805437731296571594270711399979504981;
B[80]<=2560'd202206764794965830342044748947681230794419032461495882663240397374238141333166200706719790326868698720611738576497770095921473829299028031513413006645764871893367863088042429704935927876509725256772224683015953744086483624018218240229256948735736918358525350726093634749105879349689580996615730561013265983968118882800122217030814891178993010049156962528440796376728654965849605731236799163401636189987269175442327764830120518118463557315327093395572056987847487506759620530978933039017791868504568024724032156490737483537627734442145763447259713069972647288251239363324506669653778365535098671857889127229607876920281208440920899008399210680076333257567087534312240429566899362141553633206124846264860428264473369864138045089097321223586946457586211369352727283142772053;
B[81]<=2560'd202206764794965830340576670731060913592530898012384997595854637792198537045190312773154113844896053552007135093365975377327305546189331985775914560053431020455283826852136288516408162972912611055874047011630931259749371162108174465313306023878024121872785284031448883748488676811528153996904984212265859677314945461342700136970364048556581943504526807680477155005047329215258780503459700744403536108741537826235089013875886949707797692222885679785536472316164746859810040947828952011517481886073898611450872581718196224345959708189091408260820053407752203538463837426561328195285892225407998195469255661158906449469101911235961556416445597419697561086433912828263111807936480483727488962079486494112696615030940519353320390568239718954750513158588954476782362095351256405;
B[82]<=2560'd202206764794965830340576670731060913592530898012384997595854655698204428793055853188952968160732771098970021185552956260785102791074728162302233348022058440095128124815143729094862814421376585025085429969764960695283908956631255436595842814162110989788929275920096320359742872375009745318814186560834563940435473962280241370857649443934021647612981697690013974304637164934429330275235045804674926086082143669930657060046354774707008170795037613324934091456490540338310595515453500595993482376127998160652319877602222400136620992154317832219603686973267667136796017821253829238512320601912761390539705665102167141328334178522526146286774284589905013044094857421495268324879424636282155326277891278142200041607587525172909723089809978090455636699267199215931814261393015893;
B[83]<=2560'd202206764794965830340576670731060913592530898012384997595854655698204429053622533007888865662261863778393165313169068052940333381531757860547800474117381209402874357779698554152906462961803491885427853569176016013549535480590632106444907097106125243495314448308765692597680238742245510081167393944664735515892733155303069910672330991777563751065265087311411178005199394506523132768988450622134695256417300239643484676217558298075031569197991131107678463863328994082734779579754029332584006124347797660187670227778029390992115698299389397205547907534133859832729661348510788516840089770480265926665602799324871936752372506631226798210182159517324252700321711177587423215901945617821342000804780714059912009837531588591184691454269955710642972290536359925170371312452195413;
B[84]<=2560'd202206764794965830340576670731060913592530897936487132972361815196491881199985789068025924443017771143103056843417760489205605538637468709623776308902875697069172294899932349868970704689995300187659476920293278382979681672191791229529583459381802211347104778435534355456552437516439892919669350396994934250507920952360107217577969498662461184305435250741050502041072570407947158239490524830467848106324245122420932024157139904765945277288740759706193616593354917873969327401993706385220171401314900825109141105497333337113114212775999778391787625386809618405130793309059199567925346076731200838117246427474121553494951659057523894070065087979565237774269009681104684601921449968561635066522569428718383632560324665460766306103643075923719445671816084440319986484087444548;
B[85]<=2560'd202206764794965830340576670731060913592530898012384997878600801468929541625792308152201288971991041343696397082731022670453743661721557474623393080403659845950761162119162933770507756404435756517923682707053922838257168290093584969126610704753826025165383803420836475416974893197693502366481616117231893486686599147088882958949204751889377565897540305768822254610849962412071499723595447801851602236633372337228309835763999574126579370700137680681078620199303924739842993551719704787005944051171385116376824483058886586909478343198903972064014560730731982934010730846688510634685650027599669845868299186169614150635365711745306553559509102945854899342575211468175934385608214656690316067465251977396241585288436349719348571499958527254582810878057802070985950949077767253;
B[86]<=2560'd202206764794965830340576670731060913592530898012384997595859221659761551779740181583586004108030895607377326779628517216311277106303548711148683231463376492351956102776698963585098283273700317748336446589545448775108312060181745422311428718143816213407922610998283152184914323751334311407109193042307105663891788773393194139001140862088800946465505094440256785988654784053702723022257901510535737765500010623674504938122155222066093672047933858241676983769932263242576416285299589393010971866404081737628915835628545620020793475966479724901531275074012052769392387433873883566486750822535186112290529297194607431067374843927465636880942987514253494521489461674825387027900437845433622439717662251720108197185048105993764167146828516332242715138470145324313949408769360981;
B[87]<=2560'd202206764794965830340576670731060913592530898088282862502162670676648178133443753462056840007227527426644919510674020699198870664914689047836204272473376120800888626465439576212486150279535065103293440355836600010503913938543348549681195122319043883970125373493289453377764997385780734165516053045621091304917292867022012242470490478874061704876871538270154809183301421821197428343975833287667111486919811621706045109781509603754288515315042223176932595356684196427891556536888670203479226400096275241516817877476385847985709018508158597354703048294089569771275296918101645701245100613878144152154055335592058907903910167131137418033443797493007054470789995902336817360380328319208013505110540712369908188466654469960450145656724308028643907279411916112459345216337626197;
B[88]<=2560'd202206764801271178268930936762316680501913105010182726066691368544398003195479530109402487350825684630660239371341385180504179611787483282523056614502123027619720247932146980586007747923718765191111821137203599005543491778306096798423165773893477337173848176261807441799334141584922186629784460976109990923129348547035759139886366675383707884949739100749460081772705465501090728218069681781364638585831806017306197985299861723366611806499790064721487182372391733705242282986998283537249397618436413436247264201390001089548311586937412314297262429349874030722101228556615438964052654108079472821861254114477294640889938257066047170090916685694276974248589129076729018723673603593104465913931070144972085630582321714798144677241013596380147624911198604398099217844759970884;
B[89]<=2560'd202206764794965830340576670731060913592530898012385069978872826584450213428629785370814497431690131340677385492186005028396450865621262608296182911718893481778656433722860693240620575980811605541969278264872839383959189251741328634687347518084482858822189205580774886880851405212591437157909263494370239858756124835905244547047431467144893712234317520125368721068191878721973287128615160971639094014410455341864953156798761041731362647907023117957927852386580453365100877063801391561910118034987184684108453798482913081676047785193863035285442650477296170053949546084291361837265302556209286640976667466781136558592785042685053953898001801809764465135302531056515259715407689342984630567488899782859327514246142714529349835977196566755550317512221633782204452564949550148;
B[90]<=2560'd202206764794965830340576670731060830141945910235651675708407422306564074021230163750085512775189196217252258494722770552093038679978375356664724411529381032865940742001969673098025689740193363736172428825756537044154948370635186637685423765521410925841714473850975463890855336999074571090335847641779777676808391766912301446319076848589525218145941648850658612217907761169973903396741656922099346512179414948648960895116580392397326254657273870028687606086084807502430027768092621749500679952827180659950964283138705874270071025295774225873249421693984308623060342199726091433822923873417714951787582510090023538776191573975879043280764164410747614363178579591354469717970898953088199500168126423016425729950375267850139708104974112148717815707859064839760146746756580420;
B[91]<=2560'd202206764794965830340576670725591896054771962017698253347358797513110318207619419555246234318052091438749856916171836955275211391138086725260615799568793540272687091911854108980143551768175169709590341027420801522925245078553261118595040305882763665716184456483753176108828549657457568607187346422962877129086257348228579551203347706735557072525468862572371012916411569244540324305510825257868966439021367629653922212425917711433129298842553795813862974037065316425021654249097666179509892872714970646146373135990888944996151122459329437568978345340309441831743928981646417702635459437006229177122353285305529652783868193281161936351370990889976283890229867186895715811901031977927579200023329011528533650403431261399161489801301378825287008955847835368386154094692484165;
B[92]<=2560'd202206764794965830339016479208026658399785454440490222142601687528058808453330635950368559662037469210342469952859116835506284878333488997445368663403439173625857639071419154684632338333011226537077498856338182964362303021756003381451572574531042169631934232095190277030513865002918812411049126881832634769992353924451058421874367855507756642743805782022050762102328282748371017566044822957332292865037350543032610622093233218796283833497150659231857475613769769519971741160481355346774372762325631796246155019035969561025086708813070357906382251890452139583921598829673154804436441109860113785283664467530640039246112676050000657955249600617346944390658282356692478392956343168992366875536054836484835064605237582215570598394255912522489666432889718318239587998538941525;
B[93]<=2560'd202206764794965830339016479208368471995895389154246035875271842669561675979679488525283689050874782466219875419232693353452676814611056480659852182768864090696909280891965779335848677306281415999452887309832303128682126101392944356898958692566797113318181257706981688913757874381709186635250654479370703529252423966968159140169273291830042606662609954860235130130535701497575309154518487281678776562119224492992634089774778400333930080161964754703387769597393352220422419749535182939323153980371810381320294598459282703016984990348460565329851510292263746554467675934062848607412300364398518395528166374759278405252953958371800535088814877630945790565104243831144921455623863687592341709564044285657547516992720573823630239481362192300418209711316847408305071014165103701;
B[94]<=2560'd202206764794965830340576289906962706824540759345807011553145211095224259209581517301470426085182507919217441008976879517304841328486843877801125495319024532948352774842583333754280696995584213549246737519049697864041973669861460279934945519795010299105008931598863239710947181867857744509549748361473086484569719591039565725511741887909028695429942038410171826237432392210927692086881238642287438467797621675747180707997237958025854526301636781077477837331748013713326519801216229542614292142144651608600876501307473710571653243744515953440063445779256091857975812952272928433370607755750346561127755476896802020422416093408070007240323511874635444623463096918157810084115962403216156306434166136178588467591065273746232132998933508293080736000550151540317573218904065109;
B[95]<=2560'd203899343741352263072221764351008270114544360126718504178865927068436273559235142245842278714728663140811036145239240287713803579078041342365570022727114574085588796085513999587257153002094976851606412643975974664283753382162980501145578349761069623871941513166309218480655311986944721441953254545691334132463868207098736200797304161844734126011868268899167301430988443551650187916472126258071535154201092490103141346507579563847603929607191644525633307894873083925881000016154412953935068809585340338566482466378722851904955251096241666393129645237169937744168508018059973619856247356329570589478564440217439898112557449768553455429015789185371275118058221841212546888892024628480398395899600115301975569620205348970112864652706152288444977662403786286790927225922536517;
B[96]<=2560'd202206764902130575465669988539525048080671537370330085879916097088269475521809930605250559632088705953930462963837193302357157471924500725711846602266508794480311536234004314500492047320376562061260557833789702991114465513244072790922065787545724500530921891832686534793360738457744468818937939643667519165173895318170997912068676503254196662789029994787620288463071752119037121133351278863530191412402323320500172782291602193229239291750966632844673129749931855553923722709037885336446400827968386478031202671565266084109825509759071482274946502166139739991356840826300126661843977814170177091445084780194288772824854281654423931944456409616753583911046672260755796038102587830854360113115320407239933012168683675139425821939949674990377648188387348928988413240935728196;
B[97]<=2560'd202206764794939564471673461584537890759793757078698644247341000957097508367962944319064029299203453146888311419372215503952844645316541222026074219827012885081059603405766158870581824154233311454678917117446591304245587356159585718265306222134753116040907850565695558581202193725437057920899855867509440466299638753168672297091490914165379752626534739612000127917427998279637398590756547008460090380015070609636894649182015403463308529031770700062440624739085894667067988778327375488687794541250999336116643958529717259818105941580152184505526995441154244912277251202288063867253769089590084258540924059690874387693275479285333933202031218102772407191789632347122249783325771547190992950937161788043139267588550601041569779681074851564075787757734066559124739284760020036;
B[98]<=2560'd202206764794965830340576670731060913592530898012384997595854655627984798120915398368914754059672542473744149221693957551767302839864577607833536788818574816965839387167301586597938325230579037692354095786206011033353561952696509672303846310745681846050141218965206493273912993822028983194186555884693879090800604762661898787785876157992165104427582930357461203134698473216445905341442579042739468016099309129683806460426459316195539828519697690679735822151951609536370228020507533378900939817060538966189884691004726062839702929547721005850699552703049822489313121489285233663575719067721927077059492014551144016270339894333319143229995612766807080844745050593532238131166287106438382052485238108573394631991587159916945073057802318229890042040560822656772542946808710212;
B[99]<=2560'd202199739931174675712540056306077967941486419826974267524295755979782113472810276544349651623582024024389181838621985849164315662585394003875553537854797876059452404313972673356813803710685407044629450749202143551140953949485657162345536673458971073368124930704732912953820791390265320640317419400913151724435589319863580941190238760512171888063472519605678206765134912289413136209839765753986578517463183200012667606465467042334346451985959557703821317774928447324296372611794029495816152214779819510055784538321718192560827195425146598777044736669066691012870060683506661878340644593178473246832047960890670926270186625700482907396343421837879249977316434524024825339577645445895498437680120160264876538941608430683449761928050198206566415031472124346295117036262802500;
B[100]<=2560'd202199739931174675712540056306077967941486419746332786080197510479828886251506830040526317467541238089454557133634960923331958848785975402087783780610534247542886236866993421673027416386309254063077926771884591143770308191455050854157725479749314591865925641748941978606499572361004048762419915692435423131200383019082038577804667114739702958649789682067144289779769554671692751370413817660182355541137844561197050760833154926662187118837097323509309954589897420020247113655444864325262932743448115432475820000177346196279744642936251442516048032698696922227846571970023815467298758940760109078674345774185334214659333989193496758960720397556562602504988768415400755205604687809869030477638761387231723404210968688070424986952453190405416531150021167762049092987572732996;
B[101]<=2560'd175125501652782906634249438043865255522107626785343644700119907208430641369966504948532731022855657542688312717140404161575249566483868244511417282323034242844312799407921441442351256483835966830757441210239248785379278567890066690038908453050651602538293920893389661233745470611360893901558852543223074953106020752180902944740285714911038952814517637273811390226596516131372225489434211502097361033156241123324599728406175864011039065691358128266977779619212756982025076750857882109473569399724465259685633616703589267596530246600715595051514895338308002059551777231472976885275296126652936334391078695630623981849551938144760634881602909980665334024577946772954825858246592365134033747459699051496577423242122516565320738608575234271021254450252728428875223421306618948;
B[102]<=2560'd202206764794965830340576670731060913592530917442238413610637443497844801359684540215483627553652845517043624649839008395154394273246671942269912695857391818587623945308127898773125246357098525102613562482910956543505538790812567559089530175651631780406437486130054937818602164469708830489809756033715047400617523256792397036448438471087799365000995741980704407285172704694463678529486151417538660915985841410961387514174477335777716236879080269130762667595102842375185870039854852752538222781956972758187366576260228755807371989511684145121611107677926805278454054406682309378120057048425580657748188028293908008777058273257005824812318797688609835703584717947454667936382713765225056758453006196805783960977018013400873089152850656536713271890917355968948972322180842564;
B[103]<=2560'd202206764788660476398974029422644074153240366049033787368730864220654613847216434482823260611575771796182070809092122032312918948013597162711700715414819892588296203415592039814367397457480263287174859670390777920190982704556749769293974430440915256727887346249302329205495452802887045778427742633608183197170645084245926954977243981291963986749973290624984933977030517494129321040547827678299590576052686510787214707342634667001421521834378411118612498816671298688154294439471148570056935854865275034732428283735678855148316973678921958606239047723444894997633021699197208085486566564082200506343258831258306233362312034417031663227364255075545277210833651704904133404675777958035650898244060720305427259999892000996893527312678197650580833181081235358730459603284542532;
B[104]<=2560'd202206764794939660683647466013646033700573012795278047364282823522244966119141856923032498465193704699800913241733543053481870619535907662523072646853065825567596734511220692078595445487949394048398958682984071541986737829900180665249623673538445274003049912167742627209496455028641026619397922676890163663336268753278177917496536296515900426632575498837030656341933315464470848299174319384737461559367739146169726704201614155252287880825116983996131018340811209274217003219864473829463375895754110208735887063288955839670298516195063499422038231322125099645589773003989486722202338470809812821344052266295419724547774739777651126185689183837896251922035523071678125733939021283596195216120432957729056233737262802275621481866133844565264023211838197594142117829105960004;
B[105]<=2560'd202206764794965830340576670731060913614257515540979060588785616053402267156764594366870351912319402093463128333234556962720344142346608205233058974317650422503794430372832060886989962813391971714973859139451229070581096197048399597740182836709623386214464272722832389032406601269497884471481152405593896848048169749255255876934318490669158450006701229195172356541184613614273930381525879333434943615359536407970568702255865223869901796468553095572834187188979566157894957377054275875928870585712727784715360108525012001934035115361669088606174488716874269458936085123352416087627693924267957291081623256106092779935383018158160211413604432249680946252223607353886946697723790932524088155607822735470596818681550525979986249358715633369469975662027428446860918544450995268;
B[106]<=2560'd202206764794965830340576670731060913592610482691976917240517388624189772780638517362897100563845810483779150960035245292650159065318203698532369005930498524339653585970367381843400871589553653355259772763129872951785559190069895719075038720775549186498193910072490263815406234776491468675482021658265209216306489266061003296092472313842628480214947686017767472960833938193132556280008901408660991788367349501021981352444948278178905843256252253942230890629417000928627708449885945780395283986175509324696852863866176344391175613209202520410365176560982836674899757978144410139864272683278372217442860710232212462118237283061632982049711236980214560748551618140801558637742845062554968197187980214482054578741099211455619491508253167431899929282310651332121563798039708740;
B[107]<=2560'd202206764794965830340484915842522143767413221131189477728684063063878826320874941562260425074083700142981326533581392082888843874010923008457328817716963607242766776267970011202373341107310564060296907113871883410293428616051950105042093218849495184856531658558203243891131085198251417008836993927686201525171155341455996927430431057669268764063704784739988796688321989182278078499838890598942665995057758215797761814429080337764573388989162398961620352831770525221979078147322244720064641390663159389775182739102037362059975665851012647945262347868375335049932295903590109361590572185257125720076445921419562274291216503287127747800376944448494372678477988708025595056713104398299424153937189752572270616066751630668161996123132020535716655399625518736329672744096777284;
B[108]<=2560'd202206764794965830340576670736188117535453276025371735421865823450585829665443754361464027045777998716415728395250713974030539064396598163478362147480860475792964911251595735664444911317857889134643316312256769061147357468458240704910474362684871001217791938533634407233770110571649804322727108694340620193072354676825428352549267868086277397666054788908225164239252404232148484876909076765678296246798195330071045717362639790841948455420074520820079016349133477111328033117339483895925786706071515918047467200251283775770171139602034659623190609212834478523108340369937215137681268626056807031801006625973611712055999295199371686700496686653413025535965066230194885966151536059378986393146927178787342018463104681698303490291063896182510780017389878659260919692059231300;
B[109]<=2560'd202206764788660482412222404704933769286095405837559805098592183491809490189028236701848300896126836671669747348638254727931379379872464655788261237051560332057101812643292840366609746078085052944208712731879805017179095504636583684604682109617499829526585115094989145330616559977091550977659334126656800393715644173226458854616894950351025286478688511265204206675212130802553379676914035182442404260404498322573963967342127906832315951733404926613420117781015588167886801570657050544007832141592976829066989421997887870436509705109817229841072733901189272997430505041253924308895415229681172035995803280745937231477278350982810927875688496577291263466065891598735463661982920863891572561200766932647057788682664852743309497496385780657593813632452248327588570870352987204;
B[110]<=2560'd202206764794965830340576670731060913592615767612402544189211038986557324464889377499643471155655223985232345405834233866276738073264782901724452957440954182476432989623489570383859280695827288233405912566611018362131713440679944327167689499450363155007219980173886742440974039346572044291462742451373942755343866134641538664640798698810191909530947442691225269896843849103533945156120716486725945881587159149142682854125518053392159054882093860895436838035025642565157630917114391073891681944193059147558821172277890863129566896318759202229487068025647589981077609390215220347111939004490453438613031217215152893931624769572669337958845787466815511984985040111176989809967942859680204728297378521199598756859484095590617322142376001507173877087837196953812600645218485316;
B[111]<=2560'd202206764794965830340576670731060913614262821181225330904680839282458587896329593061362364304126094005050455586261423677979979942372363929931768625765591074334895770175248388713913963837812734854579936018049553826710393194811978799651334138457926069751336862351071255708973795694079711419927314223683463168721673227881223109404562857200982267566519827301315416465715639464267114373995460847344055116414007019757268707930930678948887973778518266870592286659148108166029968697211479529637142463147863895878678583282213210659691679731042475443780035471351010060215668122245313699594191292878524171782460088263846582862069614260329274275298435380433253173993374279135166474567543622631820163721362747107817107210646826637448505964713457907232523714823541292557636711506789444;
B[112]<=2560'd202206764794965824327328295454583473818134855148208843861417797286039665294172956497470163624253976182937086736170997724216245079745241468367143941087693861997037985959805045191221641319321699826943139889442799751882024922370192648791405741207176436970659609728142450215619080271622860746895719991276440569646106068465328047374227893651979952908154813102535604543512764647150002964191314870034883310323987150883504142282568172979796132138344857655113819856164627632577773903466594156095992637149910941703493218099972059923837641737216667047876395110598387085480309303470193121710774722268543421605799235288972360130159086623365638898578163513757736212900975906711481761670905629875988626896700188076775251033082914774400452068580001633878666496660353461290470617244779588;
B[113]<=2560'd202206764794965830340576670731060913614262801756115531465313222043362502268480838274623210820961801949630154334846564959949802259666540341430978887394902253512480789749306407446708515324497231098282774448437246375091916194765915222544825080273447146178834598522439327434537804041744488484155331744000389778798953549925237395271153676413486214859919656919172423663325255478202802368938056789714346527014650577078117527729185927182153398637077820494089264284772475170869592096341845287105878985551842986944011243335236401463204702545088351658818157053662240868148029975260681107419525548107708175672415702785434263256499720512739426472587583101711985966424506379156145103539778943020863596682070008537479378132065583395720784560019636210086461280815107135541361456581985348;
B[114]<=2560'd202206764794965830317087419265137257023623453916878145472449734705315829271463294912353371407709098253557324416111136614802362516891564747503310106380026464605561562783584477910891413449411096850628447188172431805128200193918419537911541290721185100025187954521835307083652006022884100497874357457913173517355758699122240535458617232817423443992056362552960412720230685800952137610036353426551896367630076347842676894765340516279548575104826485375240806583938897052359737508206152711667562067436731501269858654839296094506383254072760758698362984335642137797287541505255375367215704210147083782931927095094684991870150758167710466658206861772382995542710204683853172018644775971715763742949389830218261324953705663478271950949772203286931373095845937556860102682192659524;
B[115]<=2560'd202206764794965830317087419265137257043992177279788495524329255051020186749320974312857088352281870541030914749533913272767171387019936590028576953390253970500522294718050430972382633384675105674708701734946433362749975320419115307805729027202033296871546715598356093686908838955208964868884285642640213087401763727581629660712699557749806162346413650648247974841769706926981310104193459105005421053647981631482628436128596870071243640538238193103919247988127135806874781563267676161113406678281100932361340162787645483888317424572845470531110412699529702804217613135551071471865102442410072541018356594246397729969876197353283500029203046175571840351188354415407971876705531893057357847942480519965360634016455365357564314157008411667907610789137732102737654904942511172;
B[116]<=2560'd231086393067684338824277196213890658679329704966183045558806936150022843396048172425392151143559047750400996672090792883321346378304879083076228629869227568261068147231016615363257653640316748966648145532918157840582866426730107987793221248582280667436439824589944731744128789907964944018909298529171302664767531412945173610183636350908175991268884877674891155994910320132590470982648911057121507233770517720135228460938594988542922957040671403087896859539334595352471770025626542200230961276138372830309981161947474284469667496730548809890616684480590778504157928050187582706928328966236950279782904076913688672574345000188516717422212596268017383488015478016565830230143551734536112308084119174651557395226989331750732218967914881754662871476497442892334076257003390021;
B[117]<=2560'd229288028038034320900572159918712024722313901691156584013686590980392806895628196861397220743475981022301422325356159372278078513497889796242965915366842163740115020242966835178470980962309380422210646242891659756648273733705121615469597676403496700741300541747029775984086828673738541468957232588599655312815498357775141119837083042342902951713986247798447043653933354170332172789381181327519730053652661736354620409134132498898372975811197611601229612676578610759191050719779254331805040294094943541721703309778036171163693164180753537044328600356246855652637442719543187559410795378743627139615468441719450397632166527040576446234895015178130357765820317106031046097093628433965867131418108344861754524568320879517697467820049498215659532656849096874782596740700980292;
B[118]<=2560'd202206766510020466852937031232994114113680415319146342058743371660349955918399213733006719379526936955853404695512845237806607831299570315569672819916137334316312674200571582610573441880236400140824948171267818719228425160350476453409487454746236477271539571975464541695440623963317444516885116369999499838623315507966540528685076421730883833384080682354284840922762166175134857006327050614846348193429839190356255837694535229772425987481951073182760962030194781202937227736853221560968307984678867837120126210830583379941307724941204855785940956162156633582421784981953005714281198256032996811369997869405565742814173000004295436809411093438162388121804338630115493239826840922144602011765442567216543165340430287270607363687873147551300420298747822600415710602932274244;
B[119]<=2560'd202319162616043018900035513183366184372176188285575388987605479389755792348615697396260602049074580871240226282378716853102453661742596058542582573610284961758306756140153809811505644117713639538337779334878449298805872771553347066254308879285800580128495332218245549847593436553345574893015987127177039540646339211273525760984827778950201891192745683763903318766371573123571608169962371709899669906609079970157622802590339594094189212692102102084577145643225578926072042459343968752376058173602416247237295072098666868200710482626301005233568466983844906027720186015048771566196958743514841859005194058151790352073076714836915917536696674093310367399522625595387292896681499589193554515363222059282337459879026301672002591591761547798057471126362152362414344530714444868;
B[120]<=2560'd202206766510020466876426282791892487485872063175143557733085721258593969019847109956077072555407729876722627378878710693315807591124462253073512891979647950788780181582879940422416556735904868851894263882506791857182017192608347983657514642995987776415026732362856693368844715138152926618335607845357987927541090772384527810373368058992445889758069998946707696034841582520250397297348425043257968546016498016771824166423568255130738581589241334253470325454963064584315972038435651552634480771248297244230822895875828511713290743100371737682769244224312241679209859180186500335957826247599844111428445208112806791378494393694289190098364858536425223626370308307590786167001984967782882849506742308120284897646228264183023358598379301303856915134050902703358904026750272580;
B[121]<=2560'd231086394782738975338197389826451963417613115178895993555052266922179401634466028608874508236513314155117172951486386023759971165587087349455480542164770533668901741906368945371729115291198588651544590082383152331612615300088785342137715602326766842734887891274304239668160982166643357898103022721483709939444449134416281086228700353753130794189228189534360676013877483264210241398716295739299425914479173615750669601128782795164508676085525012278439606617448744443962684166579859738797530717002486993098008015894555934711664851194624589029551053372068209584140824983245757098187303740017323946923804606042290975097000147786052686430242196326840409580661256463573371482175623103333873388101177541740597529249232215452122602292750890871587740495043029520566675925161493572;
B[122]<=2560'd231086393175295507510310898288104047779141058704535216436222878583140824010026811446391847355864126111033640517762922009755861481273174725269307896857799760231463757241917129603032548838731364593424640435965794312852529133911001331925441539707206621101639949288889049626503701739113830645739743934116264808769118988601667678724258294030680759598023540862697366913370903794674167558753903538819353313197955414462747145530701106606572575917768509835183215986028415079819168628943886856379732164037644509834171856174315294309743201743102402080655811183118297884743962614584030382219527018989899761063054833227995414692442043130803760896786253758952365130725364484744919795701046350720441573386584895716722318339028325850197852358469648789278091693996190532613925829364433988;
B[123]<=2560'd202319575950517408323360766403667552522472544017166111354454291289442527168463126335066849368055958269920479223561568874525718932727001604708446819578002545987936846410704862202404467069976760487048827341424846639331610401964488468232232078757593703623890014111693238849119827022921546104259473315249817523825493764970224033237075015397194879836150173859977321956021725016532844414450084630664049682472817368783935998204754298947594379679965715629373212175968591371224690613633899742239098100738798252764449949048685957971187252666102610139885741688969949220321595609531229071964307946523910685817829148215318912405249176354556662634385908116754962408790546435845145120812713604705553652883054832333578804470796628487684539309258682238712289620983568947261595328721470532;
B[124]<=2560'd204012182337778025254331819483900659668427953421422443043757911105776322406571123387326258878299337136898582329861796625770056436684855117243489143165986553135209290247355600072261023504311670476446608978137281609289482276996819301936276544713843150470332007819304110493423613153184525655284886195171212663937968525122467407021810138351019499731585844897850449626738184033429792095990778887931778344675464243880036475082254501913266137813214375482375389884056227205855480399525075981196363363147088858446588482190116248203833155716796745052800713339447179549789972996526313626403747739389736346908421859504446093226268469276757478881549711390545131049529470835823051272383654963690752839967350661672997274912172383443455942277154161690757207024677518193988528806692144196;
B[125]<=2560'd231093445479960948960659052264069615880753136563475016810091384945074129662697942470485194130403685528927679711826238416191460782623660492179434630645152334038503527639494624991376154131685710409122233915826862476893753057375073097415782086816092357933591280256992913827923125032797824279949685254219723707774839895151792120159003887368023107310581656274813317056485671403754381908178573158600454174091460191021579564843225657930360489016009157094235310206659115906934217694442629573601036669628131900449560261370572116386366610762079820195397671647358585742806266801825492047742719929616620594477137747130407943910235874548702504993897142514423737164295626702551637163270490720645458929533411633387165478136304727516670339767566074328203709899044869421308495722522625092;
B[126]<=2560'd231093445479960948960659052264411434692524651229060716709448940866424040803493380939371417673893569642127142228954286174467607344434464665205102779488619397475185137728170416814715613210279604075383662419193031680845027917722604478967564776028604578938215903539546969229000702920105982380856586821082817185019435102519842274333504444417835331881607301236057090726006697745889014667182304723146661001518183326583194357462063569900958190250649196298986287861323046433782981442821532069447472109187034207366435314359906270912192977501083572820911742635454512132470992580349284617135589945927561823374369823560223363891046388013341089170520365973872462940079882514207878252396281712856143493264450262121659712950606488130002385914397551785581036743048389203709585899525522500;
B[127]<=2560'd231093445479960948960659052258942416808418474569875877734098229817627350825640948460940348124831669638473860314303829260606340092757759494983414345379631084928415382536254288055303113457892003178479053759285609448831022174069540938262598391751486957553197199142909752553748589121249306250484961180878438934967700222637491210717301935330866087054684936243356416719324352537869517264390763379841158594959397996297162303557053895561606409737318604556639363727884780089066157838638997674181057864698645446378411669658572715738169862964575817636272271559553505052942594794059884691991129770562083029443944090981407480676180242486796234189800840463585684249112191775887440229732978620946058142313789887684125813567181555090538700668513154788458674634132388225851130008509367364;
B[128]<=2560'd258174708622143872668454363261200791536959537583456522181027942787084062188777254891896497535669429113574804430638266301748606041029172437542453989302472389385018581237579841565641807414206625599047023816234554551850020354996964747005258918829067461398507936536662490023688288666449946908170498955908422997898937894820760932671422790019293594542837528233130665218520548006179370234696006448891831064567283571008344703035410342208332446936582814021346267417246324426481769965110285703707311922951884611834976980323075923444603977280236052130534080501408490912704457548225689921301102820756582520946683988622027264607556683762240195117032481018835125067982512818517174224539287334525464805213467379321970048171179686288447596013759671269003110309737628730359997547849991236;
B[129]<=2560'd231100496177182922584674811638740000307407044082658022540316033277909814932133586013201142388306546002740699750864097460324611406771946055022092718860270262980351184090252131481702266129369676704094084066383981078635495694310896806094537318243106965099677083674384346341700849197818185086914756375931764587484745319744240028230889177207684692749717818392555542649310457902438047260025932319844080847981210935941993530409503784735773454185227748063323555999422082295803311129022166254193137486842835398268098335146382977290756297709933865393462605556583911361781743311054186645462302803554748305597630182336854125703226599827855520750033165986420944726514794371495445301162441051842493917919648687187453567682243889486800358266405342440279295976630572160392742846576477252;
B[130]<=2560'd231206284076386711141203181275407976151574390504770143562668098936577289361837003245375866856386120392244208567815469272660499607696027360741564100323172462785259153711387178163990171094867719521735829324390140664880856901378435846017490262284928470551105892270669838941037590705608031900709521272512555315705085831950304551258786156094745024858596794299762765588365902317069185860955294087301808437748985143932237210346349225314841830202460819889159754324664746707582116159242489245456317812076629256950373105479641001811763070267140797158360521508925126838892147923826322604969572157630863054912232480015799321017990722291597252219120502028266186166905646888221479767280819750563053206213144126325612028012120185569921339092063154523834853201495163161211064672676234308;
B[131]<=2560'd259980126164956067579175866011385552119373573178312884776618091139451296512242817726436728471695424265072914316600719448958874793868186053452550786616474891670712628460096205628211107755225906018475468323998677113658584896160384973028343336722418238927874135834085708351907535744285251262006847703999532921130130343252810132272047810234915516898863203648898876848134105604284696276300864815125976391580717318570039981545746570557733390869555680483368568602134745785125864863908758962667464894134129354831692033494289199107847495717886214660478503040455938917347690849715162134313884471440059563644272625831545043611057275881526951610167483149007704918167242774470523886094279266200859713621338014228023583106783271360770653188176054395377560438312211957129605955017000004;
B[132]<=2560'd259980100439136519895336026273207424934186286741139678349359620902005624919491385028715332418332110428036705276030615589236880796143422724291280152749927952995816419986343113697100440502767672870875297301586608699747077627601077246680085787532845849612814723122959106448243551077603975878705034932828164417860574896529171059319187563409289952178295382373457413668666842557610312904557810575001880125276802038472607648022041737465088162321504787680359044887062801405505560648275416149128185711778218707123318508831284273723655479114363028637521330547205521204596432872927097363204872981431428032521712076063685119196358618328413317283584534851995939467282818062395900874743897116925151102109207856172534435052981891695610368527823962428014564513041617177770917815895999556;
B[133]<=2560'd261785103039585973388517356996529198139529199916141566720812637190013834239014287562690534827351607798468015391591748693935495686741702611586544057786700363014373082513202375005516824038263877858097653748333141882540106437108793592095832626603053652323330433688925904141660137781597314166353632374823381753404520374900969926521536131761554503112738478835631339003072468153569018783362168042882265274668246373616093946280622383062749721903997158729605827396869618225635903384121114940144842580447561419512324565164743345633388678772356076755029319150969306464640441072473781912202516565017229579901311282602325253311175426580254539484737899956707485517717487093444226497446965860713942109055652214283360510435484026662425052030110261747138887348772312720685352232899855428;
B[134]<=2560'd261785517874337443498511679118168114465612038118963650705002689526320897010525254100433615721794965737272311649783359369079278377276930820110919393440690313026138279757837597726197435348021742140873712940214145214526831334733959129713154026366480015759128496981690123919970739828825872323449365020318776147323588823933818931591003225609846833925652073575664906966063300744358415788835284046089498579139974776746984515982044633607360207297302963626000425229222564757416396312864473514810897597270712627982530439796029994878229501793106047113036256044486977523463429481214706366150645396645881403705050015740721236197798184003123638801093798433504956576394168701567855553498203610082341958336519842083335677920460043491770515482173090730664327648769150819166466952399176772;
B[135]<=2560'd259980127880431060621652628369359032429184194769396325124805854537805047158525742161268043990474207438424179095789668820797559275100495404124439456497279663276563131308818517652900640309137904779085723407887910730615607091900577197216750809154727300777992983928277310197556715905926695743028946305245358516213725977182842236995760256675526791982469041886205171966021304853017263805591312806169112247143816266205580006983727595856241854417252116610788563927177616554120292127165216573170507730401474728592455243361575433434646952452965568519614746322807201025694785255058975955514512592784163717816957532840231229773929030743205689909521526567352075549575671997502566312551355082231731592412440601860570137397741143404557996792823935361553188891702747577788562779060585540;
B[136]<=2560'd287061416855204096657401432588891892790243330480824807083203673050849225369293592001423585544542623815338529400230919827664842558358386970398614298899225494128541858572619275779908718084752670429645444714210786753128820536411863750685724216052835914764325328734610369110249066075022435339232156789064585820663550933990281724829299335069404305864011072637079587791885770993143997071033956340511875478536685894576872041010593001290308828669940981647699084781558375198616551569802356992122164416907739519169484924728787437660923654236543804569720856476800884574822870160370386764711689859978202455854637466571096487683268903654081487181072419197943990781129013862625544107926630827065455633677125648685923574634960464131632362089952174270790432224868889944380717583527330884;
B[137]<=2560'd287068441618530028157216591942312906255340128845130840377365442162651510817281739877147384422907943298762522336640392676580213942949859830521149215016010755404260927681212118795854241522830648172067463787757459788305762665574244168219010668222375143164529039549210756463387767823566012780219950725972290377183786230498887445328751112713672768823491537316268506547436609311060019222935082092861206649183151889784136310608339893013562601876280174213037131592843011925834658968190998216480586081956596372420201990126373485040056925636898503758458061502035549641740430999585406168334649062422609900068025014505011712397647216908973800730057692396352381880176342606880294286028348126065316881313057197151114326746186520330431369105210833936971667032162473347295818004562199620;
B[138]<=2560'd259987178476347110861986931236063832181504812519506235015580238160866353878942202988207514032108519531411116948017913631132596389304902931689384196047002435766404908506551845786953555457418097569805117438874423373264730440353847568124171896913363287614458290056873492367070435743460629224059724063687444223280345908999629870243780912906777147460089343964010082508555256023929150089477835892067205375843038111867423419932345758573545435991904924943917227449451406471149720613537298198565492409013485586408105579212805826906617885957799764473437645642382181362414207235552197397180905071201140444991153506766690826127384728831941685992278722104044107778789205253378556323370199956516518755859575141032109529122187901826581563776568224719993496577905278919039913970907759684;
B[139]<=2560'd259980153612161872011917428050462774049506365558621064423128853801869253523363350297014480138089806621996169797203363665524471993887054260561508591790480777947882428869591177786615146597640915549899032879511326374812649933704315872637504963554212241762345817716649791785893376335299332637750072767091991403407529324610496869601108644717671848131906165304530143066346297848850220648208444704992787526557161213576750662279444808964082715093421935936280345769178291278734387394908547750319412729940649249713784814923431184529575702040665058928423435329311570318384505806931677718100489374301165934522105670151408328659600511683500693555578275365793387486701186042482808230690195090432101944179340991532508140118236307439154788181642978607763511605177445453856358860681659460;
B[140]<=2560'd287061391028919331880511839719103132604223263806420906471353049728689558398395404260948301201712390775858606834605739995597456812229259065079433749044915410317112568245453552498973813998483169887338858584353314634701428591365715160978736003931467257176016908122089672026106267281212701594490354229876872554985633282105309947284241979957803878099783793774846196883429754826951045940809333599998115974596947062826866670652947127504187474854427723250026143923274842675142792455273609581530646772636816235718074282832200651800957597326342475655107554123314286765439748571887923893333820661952248522126658581849745457032824846552684859436429655011270733070497358885057017626644800479994702409194612559528947051111372941271164068413779994027873759988537048707312699111459013700;
B[141]<=2560'd260092525707394882598592749094480976447470788662984165781832793530026782027571985535011570224144194191599050882982958399889401312330818728340741138040252789032000767131611199624328446937270880484818878957212950269764002790262736725523633162545099378523721681341643397649779153367660036822389569559344494056649135052006656766456900294594874815438958762571936685735387963346165211365717078004165916763523637244723731743748970287853927488619923733073476055776306672786535613788112868713266693103881872702616766830753774749347176648262729344027259935049118433865243685728546483986089379915150912904136631473205761790454068360921347566286092894542741737903556952180543630520411115568287653455884679134832512342024337148405951924993505563638203561980646592379393605749411431492;
B[142]<=2560'd287173788843272458376571808853978276179731857093802827670182831998900968651111002260546749402262081977242630349798431349030220507157417802584168259888602315513912892482273467942565512630029219321573348645906459980660987040171401549210570967886557933478243421981468950726983554917860628165390647178856128241078590530722466564639257178010749898295615145001365881285373315270939073552085371303082090808164415025319641244665676471912984120714174115240131912732053761158297111531511272225072253069281812972589158331381831361356107117874147321940654587618849718152086519206627465380710596095387373327845573670903993351394111867052292206381578309947697522842968382509969585841931261990319089088400794160065490543021703415556519708947297562522406483844269552140424665934592230468;
B[143]<=2560'd287061390921728321262344074142857326994928616960924069430865418273694102195319973591087557799960308452098233804197850211970789407908596238893202315297664630855085675946602725979548550428189709947881350309486865834788289887759235175298078792573392750378744173732730554965414286924693126147088223508547105127860832229015768926812544694075842983692135779936776383582967391670941792221929115555294133888172788268191839949362392927331514585048472501147400171435930549523516093840332288537264622339116158112320134484894585208923268282661073943442364048329933483382126862872476604638130441166978059896725453078686610268238492815298480389742964728808764318805907846257368352546298261597741338968735072663711180812651320549450581867967504416175407847940164889117616629519401370692;
B[144]<=2560'd259980126272148624356964380452613585894698170878839134890101542188257481570563840234491530462125206398790466363588229128508376867665327020036137338911099931792400430692520537433524514425787450610875379757434858505500420345705932054611616005222031352462361392099015864985503890556258005567692257808755844884962226321155816281635531053227486519707644859663244113093101332766205605869468252565664306330361752109490407635930201844090463949276090573731117559389931324339041381018587851125649225312106932938388150146923182454416303370125751424447186432882546648662094629861673794901504159638974453524877593806923095793475898797668381618990306164509628067892943237623980373710949035171905488422151148915860425151575211029682812941169352371466883011676079281288687320865572148548;
B[145]<=2560'd259980126265843276452099007469749539645896728492517073900607709638599451537337914714631216536097406040889351596641739462116611171514915560060787834785757043006464795282605159264445405141305610244463496871093737012504758853550033324671330686226989334973496226769642684471914104483052501434188824140146576682603811266075196576221691496821302893807815732148193315141517245940257951750892666885114444504225713591256078275213519088746137742659779456668699305786720308192179091806561663771874996373300781232441534374876194657639887491759574392621641013596175972968929901639196688627207304573628145134364163809698333036393484449545033204100451275696219500273712209231096121469839991892413736645257664236257892566239787878735263258164199687827097854620186156089314287320217961796;
B[146]<=2560'd259980126164956073994872675674818833886792570768916260222837396721187379350623494133824421308960765240747373588035855065590135607542905550314568065323527069380083288715373202278835758756884807817920138083581122806830263034068343276577877762173612466705946817905897993611090282193244660230840082178960371468861629172327017526042520310116002282203592524219650990610570905715437476897245504532268178229177986990586815135708827385400667382579857600572469252231924731565212194216617987106881968296830786769766281967843348806761392883878077793133084311887001377502712955154261099623234144008925083739921209094308693920519553064950186489993786462178426148331784211967464947930134776111532526447879693637697133114627302925464405297054116049742802246485762648321095972116526023748;
B[147]<=2560'd259874338366637845877887080723112614413890308934386674754478033709363556416856322623716047019715499712508261079545755147003151433690595969508986771828278478960268837189390817742587837096140728061887963499817965687266441716232942746088264780200884659208002323762821019958931898066367838089399929690814521663174495877815251779589069597501556984777891883779565463209214220902829385476217871560162749439383624680539557669588090961190198678152998252900407701629345901125298493583389102325134661546608932138554439068469260865744374712618706419773700778855115052453452540987204909058963885601602862911224955050441198267388936259949834484557506276092495607760083346181073303148868366332056648548153521686760844942879150752867786727404371574875346858595835028562781297885874242629;
B[148]<=2560'd259980126164956067582301290703766329651480216768090942824715571697438831733394791437367857154058102708772754109000297202469800508964413625357489338324428601981701853144285161051549086402222040734812126404804653485385570372887161286930883398622802973512270991284234434466259004952782770513791609224499780351256914828938930978429266577561597265959745663882885108561044641457773059635862313986722094310974839010631202322164742195163550838087325526151437571692620669479025629502684387288712306857798649585126400956113248297223578776985084440622622029148279869423459995251052773255393275375983763593352965459351938594940734813870188037227566012713136756284707407338994071561474594033698579317071624229854429191003442031061089873204704662456862574350983671681896512818712495173;
B[149]<=2560'd259980126158650719652387191659961597237105491790405659429022208802335262944039319533136930897362512625118502350603787738300067188682241385784630467636911958633716828080036274592203716825335103339833761172570867799732297382529774304299993843160679072729562480571331262691097035669269604031885711896405966303261712937596411054963076934192376952619106471721117566385073417448267853497230641750708163003372685422322368902243112038544106130788292755008965697722653650675479349206504357268677296978602426083451809278784598572964718467808036248471277336879177146600573189236178966204582525835875256866047047732183207662269384801177827502368584498614185170294060289012563258458038820689578511180657354500197442676612551895923456282756091699406534083598592983503212121165642679365;
B[150]<=2560'd258174708622170144950021118199695519713927916187244008983524714844065013505233553951714388220503958511084608056146799340085923997213162668522661890152970358453778390585648364187511682223426867604965488258532701439477015757826361467130014014256049623781794893018807355756109163778273822225444603434692963141626943440661465328437696492188406986158134882314527526615493627251729608589693805263304911950748809259169949751187806426880805915434943078596167112246162316291048999334364938519873839663342827364973187752253405130859464347358447309086289400620522964884934225221547922585097257810970807431625258677932962529234284596245381225910056088479147222240568254423093517655479311992886837124971342157819469004490890584883007144704612348886844773108214310462428992530002822212;
B[151]<=2560'd258174708622170042348970691232675380671787523541776671414264421696984608343731671853021996890288639052427079659314026640997316501420686603693888201947388426389730302637885900481808021267801488134125721663262558176810215200451873672905135509585625685214055601986402081680386783470004666130100322236345492507654962569876329569411697220401200151343527307530492189249015471340295219011471404646390708779849004367920807527599164697373108422419040906884156359304690846422622068144667026979450542798314176503490838382774061646072842032938200003928911438841627190142246313232986070496322255819011799478815886130580848591411632744141745831605305798428166311368188725813860901173023472189223113426777110089429928191489517483260440320574076714561088544591176000087991668177673409604;
B[152]<=2560'd231093445486266393126042524288450115909240141933374170793957431628438635185375402780015313565933279309492646613976902686203188318111648991450768899805521461764420346621476312908139338815592890999757468109067095001283799755051202575058672427725879415358239130023876469088510268813900340718631634016421508823223922700574788914166426554507926830231898443596639710442022943450767849328586350632971480972085667476629962285144588348373707001934990107915029632448370482440634174091745129330898897477276465379892764535681012858947338163740857823398662502247976576020447753353037062283459150048923179595035978886118322742350245788324827626203670339391854244543114984694116059535154921173239251944440525281771302701614588936222024087917836546971389193934371631665882807625907000661;
B[153]<=2560'd231093445479960948984154420722563942086205711379180687255077232915947715675317099938376386260844100209795899203511461101891972252941401107108099785721353949085360683539535843721894570717776293326560641187111912211377290757399698733955793414210354789200521219007236622257587191388672584696949310931443037037928164538067809702255723933792706588682144264783448551030113128543497703804445148215702517138787726554457358710446093000919263870284951288834607049134342727402398608674103220292349440084710005080976966877964084525248555705175442032336588142224215364961619880770361115144244913813596013000156777703527845477273296027516355776923521274066964971156290933386470338780342794242583051255418900686909779657268450797765292962099446397791500461986355217009035904421916398660;
B[154]<=2560'd231093445379075382106991178075649746245943257482380751350947235367856467324626677827632520246790517267069349961030075328033810116606086542333844867255636692911596509564816473031289762101840348451220889680554196220489491645267692443842707069581222416768920191407545499332212869574089794733983211206954857731286734883954199965027686827959618361707953753885337633183190959024154668269344331570016662826271357185714439306879221887501544182543074892579106925398143147624858410835392803243323748183818634943696074130277182469115775842502168391000731535584880122882237960294247901348741049288932545430893600570136614805223579710629363159404257375389250778721343441208869446468421791592851465703447489947721959282778611652760826885597164659925649639152506332888863784384639358276;
B[155]<=2560'd231093032246373768407126185749375898989322909050022103407978373577886040093297546766988601857626576011298084919628429112917414959851352427114854377224542155950648720095392688280270834651972440196693964630100170559264491253045730116331632942531904856126803424163253921774463813952811979364027708544667026209834499060063162669132132524863913823261143158390009753202684119388370673992018572834370316600858932149821542735584789354856280617509011977582366776715123318507345401833524591532479684609192615362690664345509374062305074318273272003833645644388529852992868146957378007424016157933792370464313586416645135304534373881357823271566446542575930027718709037084121044214022272258476278498068349119611176740574852521498269280365759654027240471360160339743547356327381914965;
B[156]<=2560'd231086420609470362158746030186711036248990207031256369550028166403822757724820330142826154151778953564350078846742303074063015043411753683659803852270704770296177490993725164629421271405546054983717114300804323152607572885957657408562425603586087686550050745744600196706214544888120921018755156403883044750934318088742244862665365375566648312283768889939919005119902871818223817680200678572974708667105114388160980825202482234183014078153209775849606409704636900534789537120998713648130808371249598885073047780760941099346917105009093556933021046173369803361720631233276553873126746018224620238185435065403580235914431780634704774719477811559212885975321322710417851646850145981403937361233764275267582305749894749273283934504539207469337105883735405676951514619637486933;
B[157]<=2560'd231093032145488201529968653888856418583621269922350012844018871892275489125470728225850012407562360972956678124124488372360397364932676287033317314492592524772932236915163246634041974484616511219765841883327981701098528726533414497010140970365046357513824250809789829431471031642476940317076350791267136404606592525959200546961161992904866627549895004085670150595374555803391746067691473543444328063669991105834490053319478832864918670110199314118343753965424668150365316219243119268988673799129388904024235164899812678332924239999020737262597850854069484258676750262124621259616320965000314236156097485367871670591015215968874570062514805859171804969997635693834563527839014349015493401921356615218381440045537631628849125922345604474422456319411377909214741499473122645;
B[158]<=2560'd204005155758907597436024060601092282099995229093256095281359347897471581186378038629636723589106737007612409009616327691705025366887207108726267877292837062505989600577175180622691690372842416823891414332562906603732203417953351056477115307249961465070447997610471170457779039065888692938817567410728625518888494240854125568340711201363296040125424338930045201703848282167213888264954570979108056697913955935974392085466420356158771818247906157421307718991415584096615744886976984855700741050515636625657588010715884312746233303879719180288403038168731552440922564735243958162290899855142710648568312847995390365593834238274008661157401084561053945706146465883653572625303028190397882305907188301367854609455758828765764205073865407395640691471688554764453342730427651412;
B[159]<=2560'd231086420609444192500348747246842220448286212547682031861375549175913763493666281389324725570743847492978046120475118866192311467493283521978761691203214750357606079899560829138871682083376038156423723964454080553795410042624888034245659516154591273451752053819385293674925658390581062055611373754413404419401814659029457672486622020922201924154565559365774535974942387050669068141347440563953546196506310419955029218687125220002257567765657544091352895115212408693742158378243658464134833387302716855052045047906843269405837972179769244895427994248136668724741039706736962646527500920601618759943042641930207758857791486478537858113408546534247849183611581431030718361639804121759291537014212257469256316092537397159810870443683503961929157131902333250712042141170095445;
B[160]<=2560'd231093006419248303753535392169235801223970200415968911707512963942306570666408524184209936850976219818237261049543098908689062223071092294189196170128172047299113934439181497094432878674402921668306722535774058138019775089028104764131336087913599942222035513609191376924498360182371407562036996424138711674062129594114459013263208196215566456087622927303892985168619323150440042261358533863019080332940555000491436958200876340225759749520144246178945618071701112250423616727031156806394968565776563015620740930727239362675910191793917488147911468841662725623823247196848903466857702953894603557229450094189043295455384356601727473731294704511782695507735543432877614014345758655915916993917118386470538278100661106963520876310873701455312103621205480550362902547964187989;
B[161]<=2560'd204012154789292576160026423358413057498915540655738089530575258585660961489704757200453283848314746330446796490160488180039206620010527063816623541353382358349136598851130904895704902438175289528865409307168332694153229601203820264853013819831792374656770326703695054597897892243043538994683595994555138828434126863638195579827228874427523825649424737755812819593187932185461657969197583025653378486265052072789090834798507357316865003436668617116911066176859547670830920485337779901871476650245541821353354859321773620778655410849424108177411357433216074142922908562372388309847722786576688539422920920380508081955491393126317165547244673929566018863612605228399256694391935238854086833731812015433946129299163705135039337074193205395329228182064915379682749105204188501;
B[162]<=2560'd202319575843300227673903089141252489974460714311146939962430908176120128393784599257861181650423306959535593001152743704727771515753825194125088596106109685374049535566397966351880234311970525676297096780362146254963201892339553507960879955117249466800961575048649154975535014740150791261210881285972823241187730489895926222375880997568488398454093922406051414906270691187110237988493698616560694215295096884881086802899407019718482091491988610600976861621306449102331786432000813646642832025443552301121101037732830559510993677044241592339687646236301577704540389501949431851265749164918356165077520028445318511172471504428694614456635228139556773936630654115241218513132339362236203894849763128751409597855117449166475014838667690234849313406907743100851190341760800085;
B[163]<=2560'd229294639681267711357368503479596289788917138323781661056907854972223647482476618928250349452152109612550769890593079790032675939013147891929689968600806730716313798877535588440380893097131731440698181576704571319891952088946899529154307109285846362624287104174979963406825146183517772223174986449524695116541459017704312285205246070367473581677636941158242008787236773254550503923680672296627345997438355538586119074693241015946021217865912090260726175688863631136850839343590535936469643355227331404641198686532728078783113446134531305654447166736497286389150060851256711316055979204623734611156154491526515645045263865175694684599530280877122511251580496095522499913609719783342559133111353183891263416578979924597268722502326434160808749716851401847437461353022182724;
B[164]<=2560'd229288028038454677028245886056513491186047260841816845959775659174474491155253241395049846761528679387069517747759210278648432013597318421671170723855764334798342502900990924012980016077831628024761228503223427439620646356547005836103887315947249079011804049855490644166499418963703032995662095556318162639664996734510083787082177544386189689435475972744043220738543020391253512559590634682938742378368642854670390535435693475756481890502527013074466090145746027951240038831884341546574586561622020029849450857745467454584068433091223792840489328520872253521093903577439511730715127016175006939102957628433798036130210956300497474822034569126990300764302458007624183123179178844823719568286907206925370924879318415070336522788787932442590128184194579448203047650364577092;
B[165]<=2560'd229295052801360265178448360533930584056580189850438400410513529700037394486742326249030750532125898490406146154845861746389974443262786792394023512949960356749995769425336642408270495539285062708454722990917164414080802956354366214121575045160002462786174120602926295174229339647104110302372869171394309043364566840544260228865962991965512699171092115696287169671010981166899860302217186411603883848645263165875689893004794728193222620142529289872770175814408933947612083904365181797708293406846744526109316986225524846668888507358198113240288259333600424927853595315947913388767821480346747016231589076993743997162961187126936857238941574869610536573018504307964590749061221428458887708978214414530833889915997661511878843983296117609762336038872790538127191417917101380;
B[166]<=2560'd202213815485880916619604627906558872079663623278646930155399220419448701997387949725761355385419449133603388076505384434125285028317541567714220613093559587660162167850511508416740730455888302335443864193673344797832109048854727073099041144843919410792473661019095303896743798279530432965189053412829792653486292193782055656733610201236696498033986248258773233200581303766011197148082496075809381860505470893856764556202332598472631405545345151996169309400798851505741020631504283991787031760248847496970342037061272130352766868968265394415724740441393159123362241741179317249875964636862387552191405383035029748161336565238476954667774735907252983690462150115477969699090252236127185687343143260265519459098205126416921678432244380755094544448431105777482526836433179988;
B[167]<=2560'd229295078728924674313204580081775326906661853341544142142789100985555397197149698026858219826187179828892149952494704072935382444123159284203518725449112732593245504108768778716383585806579829770251559307226604680015415586285168576553120876423198120351829017843507102816577386578467481180083815984527357786481838094664014172582301734935844232850612727135782806409886597959649212886669265291151095419573221800068597431844868590823878079000373765866672182864553048505291999274221470226558917139051379477657888839495254635818517146506340824975422345555348481219572441347959235918113155631085491724882736947415382351806228586650185788552925413639767407793207115869618364754110684258002969764214823090970054271294152267813311760700371769955462237453822442458785544324718613844;
B[168]<=2560'd204005131646862938950248660925251077798403324041593296192609332811564018150838678913566825595399964116836556909715541458515235569212514191750655957344842325271637031430366714543932303655377154123347836294336575281208365873934835037032465392886100316971122273369932907060356598840167210082697675463147733353547105911894086236450923115232065854239002724946928667042119758103487515043007954852149810233681221625654190578067223640992567890497591882705286540072059542872582721653900416973770201800375249201596503726949085161948630037875916062339882684593509512091503583271859512228680496419365984075915046185091123793308504470061572440910690525083341975638720915136225760480777080242322113794815378478812169049995328904162035566172636733841784073625751044323204881196720149572;
B[169]<=2560'd204012180615997684660888265430101834648599028215049972427965307213678254102643189961334378091195194526037623462667330206424467315151873394876426159380685623841334068470535108598613238652663228077402975682762137404899438704201533833504333200839729825557514244668564445414648028382124171095863239967203495421111337961139406794641100921879633871236942544697751337933984976294628666285698880204545835312363065148350581140108196860671963706576470107381758451068028685840108068234462637301081936268384192700597599297623390011340678082640718202610686153273785346424360304399464447479934789907991784051803192366185388430436338517275411280167014020762895932026355543593183788895783008688039057381990658638503109361953362342397768564585293774964657846455838051546624410008153314628;
B[170]<=2560'd203906394431874702272089629394832350959578873029663443282255214919409125864416460737021532813126728757282682741389046894501673742635206142761407950299040144733240850050115038230324001297702061127560174048898674857519299774410698497599485545029705908568181716794415045445609528667620968198666373614102438669573506912369676457953932635695126130655914360087368664575307674568843073781386689205340563488512637347650255037302353715183296943243227395948570729802254234629477074984786508926146710617926101536422419532872188525762739877937813426085159141788209276381182577516544680997613530270187738064081441139878577030946336132123128655081100085501566141782895500834883426188986379849882416517963653880594907231103683386087471649729950600988174865265999090851376711538324030533;
B[171]<=2560'd229288441171156188502888140171820960621670018868972247372223703998761363201495464537855320645469461203983283157311820410740272761221641659050507280080171700029880321123211751724543254448947906053844739767876089782835603543543195760163694095611512528901985593802299674857238013804073295105421817997383370678981004245799928017084769679094465626710518590317742217787640231579044337017812689228193009880275510484073634368381946728664485073927033276751547800347099292665113677239497968827239935772904507465139241147308692519772065898225499843634192033496623375960290484979024611829834794391821683445144228754383917567913486119574594223837100196851400901580508658279183983930805499411545434189198076515361476033970782547182799551986264226288009333037110150778023470665766880324;
B[172]<=2560'd229288441271647671111034255044959667831004694847297155226592520416017893323272231084011713468823555516968615830573767644616351548093770861428868218147058375792111022390056719790295208386779706293726152632315582800814410802438590250554773908754819483196874572272752438357284853424013626091111013367201764354672471411360921162934906033433650086698723281806026916456033373382938280485563689807427249900015429077918051248495490682633745214478458771075590354085004345399229876234542491421581520461638913418157029236461559082151763566780003707841672182927867983086350765343713401674343904609391678465142656438386337656776179926102976718786671343823965757141581704920654788098474814069244544591811085954189713848398863496227144109766860555158021639342043449546685812608773477444;
B[173]<=2560'd202207203949838344734325239087857724517619770967131578848353508908116324990527042726427776921623077412619650237427015522432933512601198155223870733609656883595927074611856620386770200851263534616308693717834719552190158178637763588703241096048737647493221820381840500871159900496617264101863317484693391556302059796931489886752671459760100890616633777319733256701695089178046530636396115968984291588385413585295533022692378110108128543042800968749139403613983023999687886486871832745374828684352777425399432727457743546813419288176261036858814854498998390021297788298471025886516898222797810992504972767307314721064188087458894418279061906795437957052221988903822868022452092158989252251540149732782379140395293026186184017274090429164219193860235610850964975044206613828;
B[174]<=2560'd204012180723188605456159163238609525978060722333482085419500018779946675248705412331746682320259134895389396180391526969224671210239248234158717470605524989825040294221837496467448413711046347419223425229358534411627301126422751550073465017323023681564452021458508055105737160979343032853370309120582093433508118790517383335333478255109655283564899496111120311380453014911421383867243230804679720220238206296835849118489721086104250113581298936130031191350976565722117229068067596524759846480712248317109771428880081833280033646123223595684489477441228254521146134011915327834141536189696906089225847096015365922681621203509931886635730218947118642822052405437135016798384261333884333894636125012910609325165115703096740948385114038036274391599089251171731693616462386516;
B[175]<=2560'd204005155859399086431680624108465004758243909345781709238261153380122067882238798154142358482610003434051779268922557122696613722133857271370084197260520027620491745304958789902219510676460745684988940012430070211607565095246307446781893723622514773707181599770585492513726573612628914154785489580056456446441220402755148998845656813562482425693164897604413222220721652290530497333910643897926892442643771980108405056373078958991491487258522790987463590426175095245321762023071869864935826070634613004708435602757659963364956983325487273786435416170187133807655452848295432083640984017600895308341620462339128103880287662051338479536237001316676543824401016322588285487846670892372781730579976787712469793593141329874538204894174721557300385844236020332133194509204145237;
B[176]<=2560'd202206792242145464691919084493683485604134991503026590533149267839165011993375495863734624521592314341368664553791305841300752924662060917812686672898534626929165048064288278375344275684374442227285706745570562853155958962975152428390891444953978885945185661942235602991257108330496154003779819970210025996737157427202437853559381208235397293106555055739107419944744729138700334853331095888691164780515312289037984041470131452813833534204304214839965491430080468492093567006396943973438363335742544451732993338045796006830527123738326872166908980944883285031520028802527648974233958935502344013455581870165281067885230000063247134040858602703165137903605780613236240646184497730387134997394841197176671897060969455996278626318824535038563775385903276804342293320405701701;
B[177]<=2560'd203899343747657617389652787630201983486567463038163758606927486331640787550287914722830173139967864032664390289105698408951405554383175166374943124567204033182983390331994087123899628678642117638766986999448408064154362184768998135374106930802784943819878800650417743383064202050598678759221265793615912567063358966265122650754146939222900309526777620443170818258463833616640741916052991775850317498184171818680639429323340684408804012845823147262740859889671188165426284357362606534867024221022807893145905745852493598872328320351438718396764837236837799445222689386291114328375556187646259938898184256511939550192313228684533999341031044772954940161102591453711205458494083285148997729957412380216754010251151493294746739267408225381908126612036390819444665638802773333;
B[178]<=2560'd231086394688552847070971191269254245942904791780026747027870077453794436114624368044094205509272725064374093293443819884111957328842521220959957052239850965555558310946735754769025911596232550093639962830471264650425834026553570468925223645152955172345968444327180983835080663129466133371399140339169606020624330478358169149128020622841241673466875357884385374730175091783847503380170730715176506645029544057258235529102036688875725691920024467554936711479544766418290949637441197962021378582105383666797028636848970257247672220834791877149454234639499288352712056361159112484589228818412329270622053132512894786718695826244743181180528203825731622244890134495735095142989071429594319601669787087805831977544705071182090708729507165138424203822026942664428516093795325269;
B[179]<=2560'd204005157467681522697940939114803044857820652799427711030475962856484107502182786352411361912397702809899606738210514812367829310336980462555694302595795299095119161508192861977961414822878392529415552103602389885088292381821638046619863163009991634643836684213088180994988231872305597520882376851284342474036438644777106434972735536041368260357164960173028223854786200114878572865040469503302691572067693343133107459308191960712346649703396612923333022528971737402766963516281510760991720720938282103514921043938405346361863413341113001463734091796281394179003726947806975335590761512429235030100526619702228228371730701006690155240552098172592704465807492046821948389714540217459866395602295615586844607509728491707493227889738057181135016811930949027318814398261581141;
B[180]<=2560'd204012182230587110470841218828563783643104136616849517406134776960094829013695663626532229783445402437641132122188823400878668352625308241428239795812365640555235267140004643557308795705430889577245716819988651727391602172326360935075387284437232824742562263700431536007705272290284912631874005691334736639241403938806648841911510726575438963346777407611495905356759887136083183344093132047316814985795452245897026605888242486115330183792906814610526341299358183270196915290786638753085523999247201592700854965327038938723951058600487724192964324027742285712767214155673553490663396253771648884599632904091495761217216649525329815993877358371422712818167014684374370092386977612651778693337127547086497196884269503415008394043684658280830904636768317308568961919338501461;
B[181]<=2560'd204012182236892458400565692688738152134290838513328052847322557997202108113243857546196014052352059248702007731655049115923833295918930858110329236800829591310913148788111096792117548170864206292894961387696655146788104910257437023824604790965819374871901190081823402639313240031318116274046243445120689672832101845220893024379844844091479651651493737209827845266858982398054297158748293700489737700047571869736153054339070204944422024998268123423228731938506764848688244297899900110805380204938209844512563690988654805929620384351687506411330957111520740803586789069926036334914482545012450659229650631598933628249776971744576866445277912093252791355074129267674464212715939133171515432253311870414788675900192313006252743771172030891834591552368053451920369181424702805;
B[182]<=2560'd202319603290506025669017752615956701451031318071651291335463600531560195020227301216754526755671694136420828907192981835835398713832165169829276281112654789128265017578877300711504213615018225065233465295069623226086240203447495844128024278553311457124980883027076312151525269242135013691391408619882223012946484375544122639629665469439022048048831138368529209442833426290039295364016301965207810777434515521612931844380759816903876325142059541858040829052867416271644057035448768366656270380771806757682513949201677847909389754833068516848933739391691962955692720193955710276043257091149459266465717384390875920712954523162291233355919251706283771262648205133118494589331440546616611369434419422705494733443916282006193866293791220887253769519504284522649342170358961493;
B[183]<=2560'd202206792343425116191992707545525509637253871138459865520885564683096329742258182385945962268783544339208591168133695709657823650393984986107462656223107924547475001390410438439496363215232280597974601669136944159576092176707894670587410340068783597708882435729431035547857700813810657600976252106068281554247985219491622946562173138851324102314713104094048187666287410521202007060964586593390587908257870320720891702476214332513060919632287694384668316210913292980944291096423533702456495255312328259869961703980617105595752082959328978546421866772746415703327665936326986139674835600069495623223065530556235031935242548395597619391880513762287357154673293947002344835848424012645209850891375808645234309806072711863627576062272815218127566901981306626286058415125321045;
B[184]<=2560'd202213817207242440453469275314972981622396236295701371164441063911520131673201084317815815769170032886201655413063677829399098684388769962949011107718637096562415614193698458471947377393125741140679428304426649767105688587501992339488684695777108097819050742023662243512347583431373808965832784018285271849887994540384822252615562335909633806077485200091256251575464916504704135553079530320219267973717621787358704067707014064007778020923099071533499985688058745885123669091302603388372881773719665994184361899709135857532249922819058318702656067340086946672577712915728018258148856920040307580766327125206380975238041624543359130911452739428150312627396991995699240375726211565688144583729417012083247036512519631921621817253186456059938272058258005973077444328919749973;
B[185]<=2560'd231093445479960948960659052264069526542095629097925303103829162582666042702565092374677295022478505297210687648746155497755920751920079141952836221126230829329243762039410338893429924501636590644685703155094843368190394008104632488549542849510154795381325102936525729927083518831111636633668837289315355747520897661731071389115704390474505736761672824367934824868609668465153427744911803794043727165566658689835377087574819991560682865128413038869548364653256536962837030050021619263473912494196160419692729662310085985914059480753758845532289268133202186000265121610066334632119940990447218819873839707301755361923348535277439997707608194936985498281921568817595786767260908920840046931261995243161049355411761588010804687570874487843063874212094013949605489271306016085;
B[186]<=2560'd231093445580846515814327308764161797092211252020983865527240908263289742304002972782585757079272058413132502992745774652562778564912653038350971905278903564075840542873203152641722790750096078601396602894013218107178985456542487326075110580073634871567947564810027839662616074280312347165174652160690323577669945824881331302787576537028397800692393100150692702066048432043216435279353470271829441613064853165449463318806357672317665560005344650485318032798511618996662291008227394861699358041377186877089981333824357633398031487821875798510203921457647751830721999382548948826579510713169846325011808398783909915136553379784927368057808719818099684765005915696072942220642978668172424663743148540645550427434349458323674227884248556727196942958070107622816210619639092565;
B[187]<=2560'd231093445580846515814327308763820072487053360769108718688623712578016000007204839846303735333882843903749197390456465427033236712370223393101219737228886657105439511744689511379153566964207427902725174592270916541936136012722593463809134406900216932096096751933272228890702392322893363682712709510483283116765684068975588607919690886855253254248775620645032238214715310150541336373474563540919602347006802945420087835718031310064774711835725308193828044653087328190093173333035443927897884084333894732602762716045996419898544988924252951073696562007499058785710031422429169455840306147244657308010653644595013109131506324702016696801357503436236673237096950033288080168195619135184278740137113922555255043228262963688591732307698812638089604984523753929197405022530655573;
B[188]<=2560'd258174708622143872666986284950923460007365983196207485620461322783193176972719014845787027202845195668528917523666892030254966492999944649378929836450597124499254639124176113356440670662814331184027927719105119068882836140838020342871480773881408443869714044053924702564490999873814844543925842354274989176350500612177562953233055887383075563446662474823579729348820519345886091711036318966611306926827096443722552015726644336276283090882771351504751011321179009871976787995986309659602029576589261641628023927635271321114009267536194043050130141460454594695142633203026519101655451904805145916026515239304279405333731939803733357866382235441614681471142504998762630192878424910151929583766280260595962872047547156796512248104814609790729644231560592106028865438984000853;
B[189]<=2560'd231093884533974065781840545383045929529469521716111776839424268314853153918447622526947557851493012790777955130927641667791618502179268417303713773985655968532955280611835971411148869758435432473552324117847653609642025563507892430604861010167411417041231132627436040041314810370953002646068607073453115047809205955824143771667955551778497234418187494543155426857504722979429955076416838047340835424546533171543280992536052879446519366798253672580660034303966730747560673474191153472440367350610850984689535408443928682503515264886591560478662969606896978074232407282904380538767984687399137636267609343474920283060380799495800449549073234996034322984101311706857444820426099482427815202623830238122343980708778788200285247593166523272884440161216508984094653315923924309;
B[190]<=2560'd231093886148141596048948578518791971278851376299661133959111083948498666869811669109495222692690861221798641756323864768619258979279904876306826468164707575156101419150469367626500118870090283431613053577807861494284342750143111786032960741952941746280365948418545292684329272615622202579517642594671878846025015784520334347608681730177384383508516040877650726020600337539760143246371759343852476053783080709985322844769562302880832244993022920938584811006422755889213016469441087243062530099994663984869988482647972213299087776195005294225142319586586662242021924310231548566299694115715544953052829502967162274034828031592628296373352076912205041105057202539036884729750769855396853150396269746892740656892383976791729962806485098232784467500907397884900641704571655509;
B[191]<=2560'd259973073752679457445827655963519677475377092639220148323701751918222085479367868052017441496065238148452689512621578598880483357328343018115077382680027416268553927407117160037116041640775158385944775855010324327658614804595301008106810271830512566667461049855013598283606334928189627967068486301226788916855944344942571115070706471488292804464298065585089625469314677116358723771562777051165411786784276629081458327913889708017917640244110852836587579709472106122015013622260956578973377142576160374825546282004374486679065741295171132050491487908837948959256916455737805533386705569551853325227169621956857654287718964387164924124410347898841959924314853816691792464628856969635499596966265843171646292430843715152279174266292044483702017323987155183696356985657447765;
B[192]<=2560'd259979685389188785460465944470829881251033567446823222641193030391338596905849906426165817340056798564659926024115606990065087675140418621059920547563856732221260095854362408488011835433524179357552371018206268320990577465685935519256813958346716293237095602948881705585139549002564334763394784958295877470633007843120718281826078371490815575014188417025608803929451407680455485781209676463347201261877109850540597810674232174119887751190583045971142348901276349963368843404178069967481590829956946147217991929599633121521185737855847936648699512499022167437068307022824069255022917270469797920517007918390074804587386035095132864204008609158225427920926727227267627043602643423181099936342657659176705251235357115410550046793741113624307001803528834959293964561092531541;
B[193]<=2560'd258287106442802353104648515970185636909137197009596511266601284505061462866756043543414069350054084050126161629167320455628365574249596699078782953634400132352074467540817923671307378425004715739852885011802251500193922337972881648259705831655520479745073293209384172756902351747929833691335159979816864253626835870551302851275602270082325147178150509003482435258718068595280742476545158153144853621527547227204100740681679538101405285328962876353044987137958481893727509028809007260668002780328803088251467968885782586090195441098784217624828886086366402103113261689800169714950461432621127188672371590501153155874055575861454397906499089818373159381429593064965038207847294854010519706942837027042777308287657975602086999994946115707308699793356695350371703184906605909;
B[194]<=2560'd258287106442802347092959973804359083687640467220601009073327065326845475626394445539600563585555040323008596319458301129903318498194030206856091979426716540384625195106513894410182753334308710607218273949566339394749793208510508154779006313436799035623025910993687568525442822484934825794760277443543952012127868781764234873969977301211360279927813129226827514185195780445299492355316188180835669732524666638201582576066274528109418728315411457329710730224336326677376695036545236327634892113544114241907842798408034470352934856915986108866396908286519249720169261493440159463880080113513023826392245072728803989310534128161867300855686288756886355108226001734984108560260170358037506435618266849859917340077821704957061555633647971332991191254417071723295251675785549141;
B[195]<=2560'd258181320258653194671404109596873521986587470764132601274133609325462630827126687821089832159064473320056280550127378223504774198442872022470294174447568387561472023038045122767087036544823792132611904809364207782793361937851668199140986077252361682032764015155691550543794696271108778147863416677861616715541118739182269272851259827632214307126451372149597538785135601259805048461342880180416582454674734774718502918110458006823110626656412332272267420248609589454965934622688474554287639914163327240798726075191973055927944487341280256981549281106798034349216415802477483327847453062295522728924261127844762191789641857135901060329217467971044432154803375788767765076999388709226434841763541753552093511175604245174858836015293403905851623148670418157835335890237740373;
B[196]<=2560'd231093445486660483361323408907305418868567076442482128452815906386632134958442105404111689040411425722662186234352272490219805697340870619165045251549003167520049291350940752458518924051592747049797826643309254769074816385405321966080865407748735900997772487813619131705889776919860707296194903978186353022871313286554947489925847636651578283126572053282729549530915544437269473829033362998371265302112535034814184804477228603084402285584372260049554570444440527813193554387535431201908877953491767001626492979168151067885483375616975686578862492680359130384228064695203326150130168679634556518262331922018919047962420482359565968614893770749102905324090413552297333149439043443338912377978533436198479189220253433925757993053878234748808259011984575741726509610428618069;
B[197]<=2560'd258280494812598475267173996459587417690300315723127788138539678053347877603257977512590516085036657767246050518593975174897650388608703943824954639211815733562599369495248878340129981438664666918954382401783194470650753165811961514039500194204581429909353656817307384976005672249192400932691941566557197094195248434263181020385614099604104502261876462651470078503059509438790367439777990104516856939345503033373432915602979517081177683313583793313237737571766523464737418804610773310629505434503571277919268997634988396684729919014844298640565487429587832622672369369945782499523197356238742176856260961514477290148499511145920192264012533110478631820770332918796275284174951188973312539907491955382750824055214424442890970557205756223197432088158927650774446749041120597;
B[198]<=2560'd259979712930950166503092892632425040089291559025261300485193886471615729424100191793072430631581059391653504185977102655344500137951262154708447329188569284663730776951683772121517133612259725573701038117912890291199788501386819611396515611367599635822733761871927868865622779327266473789628655582294091296282387618603366691082751724257720513113956663640150743747774709936385973915488170274891552806914568948832631926425442824555219691523029215313723489722840635581281833790799563890951546189762671807145863932270066179501957573698271989349661564801967975293210272320968308163627762183577880205689099859450844762853288116197520130642011025999305688596957195189071211054842234466653309433572317874989191210210675389600626128186366498307898892889183490266788831502835995989;
B[199]<=2560'd259980127772819789334666012802296397538061819072247983763413673389767414601292390416745377655103722312110495504047717834711412764023051359911741956702512948636862647858976351132981254032174688194364143711071080590741820050827925818042183247336868008414416117948762720935981948571923932268999919537821164229588608290124169704226283892093887364025716796193960389306933391587251092585550864200320730318169756084841289657175959269931942020168627753213156073011117916725274250862343081879946283590625979756323734224512223723301972372247645120158052968430438985534750376241428384874944493370836899986430177133498396244369945026727415611453339954229182621010888340681257067680376682690526420481636035395005170749334976845427837578061487547189564420078804732133571085997897504085;
B[200]<=2560'd259980126272146982763647181253543161900733419197463580281873068431241415111530978691414741208516491512519267083863018017232791167123513018469653607592648977166631525703508174532820577648609687312475323389661296189693850264107467841967395396333183561508889657604384544057584395781436388491489599992291009406882277276681537246060517581765537465266734455367331176273740833186978097880549416088673327242889442010122186952519309338807181684791450943630188527868479433781973619449657555096435433494214151455341054290357418361003859602148373051511094320658736853072652529533108850171764993458082022599646512558000255783143714443248745698896022388156573331946793079603587534343912187294828144447929650310720991109083387715455605779478036085094190395357239199022357697586517071189;
B[201]<=2560'd259980126171681772037652650891592752749243251510398602825393040470329483131730834746157949127703716791592374447343334013299633312441018741165196967807012883381207120711528831215692229211409338738435861770660791400557755981963024287575553750454815429643452118582572794411024981121997467934411025395171554578443022108514241903540274966667185630095970874627718075153056486524748646009994773428972178390510837866521366108990713421679167299642088139587070323517955804214975064529266436791969585375525616010873178611582457229529519894843249886299281894059484792029545973576528936674376284872041396946154443663008854315127084361957266523359336617504014231337500385069688068743627499219672203498978228651353590123079178741824271017064255729682523696467510650826742649005748344166;
B[202]<=2560'd260092964660497802300766944965579649220423760328681902547901152265724909774748694845540659911515519657591280354180290840887413383578734995647263063262261250122154131952050794893235665578284854830256355229730834889179374987480007018665965213250189368128116178622736060137168851882274595091999261105690377672658928611058704194762615470955884938146202996985780860805650582971623918495987449836972590122689113083905738590788302238800480831085795472335294757658266426026664481481521290036238382042657623629466445267746449057528990090440873988064666794169769543214104317182087316057295359997152857562230487890184630634201286054677890889033146122579711259046338743320741197495264299984764085732480694178979533252549850839204704663090383945769466706556682332673222615156921816405;
B[203]<=2560'd288866806849951186600238962038583420167180865226211456200228340452686447674645293307380886145096012935149995709219763281223247647130002731165852719570368344036352923692505860485913073375177790107814886393867175989426075888632022594704669622288666097759427772676282731704933309193834700152559176352806281196980927999296091501775457702733753552779271774636313853669597613163031506443786585975670571768422044267896760577374223341613186983951469157148872927802640875109748960633975208618970842224186245424793479853686855247830184859526748919573946602410360612787379693324820061618891427694736875635005749122825843843114709737234720903953037426919696639416759189937121674070395644184578152257553052669818611090164881971037029807725517357940412108953312182016119649867762390357;
B[204]<=2560'd288866806856650618775583446513344500044000000538997212252276535365081895784780608878867104731789378591831995874442097696956408009124004058832771355105374232412206275449086736207799689019181983451765596492108702817960191189782542915618894494177746615119496332626774388437835940155273703540808316959186591702252610603796992883076159925577920206106352318494685813057726754879116556612723029732148600667386847807454258669661862119608574323772729537007769433751450457651165387971210731382329891064143708073916255349167125213239831697435993030545112283531930172442467210886203162754079803990475991162180987440101328234334246441575213276060404832718104254649417350875276903831103939063522663509335801537170040086849436115674508098602903760360809411055649078054051269627795035477;
B[205]<=2560'd288866806856676890657735030936709480369657514989024951186898409798406408095087937088400401916713173314221632562771981635168039152223989305773671834137393653740661635271682733352214533025647238442362744224464978974839330044551608979196696921396050132928578076495466523007690643050790518153435852199056627438086555920010449017951126735358216343779528275942631553999604143657737718152056858516189745959447696477409594726247563318284119140654792818177134893176824552497426143720235402854994271575482052369339702546762629278561604900895600130942529626755754670326344957899952009873379264470398311657584413385570464070563003729250402268377878792308653409873340212798920440911183511352915504561432580736210052503109457186010285942917855179004519290092613845702511804280907060565;
B[206]<=2560'd288866806856676890657735032430093170787908991064330105707877798154434324320729625532675356647882755162054774547836133280664155019744255242535077418500462561072109461855633692295957705004850618438938077978394181928150207436747476227907511088296932626290888222160138389456272771633323418061728949832051294372289018141940621273094283985936319247222420380608983382189000974312118337561353989277125341811702820765322887707661965466121418696091877330242415622796587308735870068303225090084582718502814634033614941106617068584034852879518294733970514966788417964149300865343929116098845736481896754223868001616713757526766984595462123695766433061990979437369348217368646373979766635264205483738860598955664195484215006572043058493432954332600078639140252851395810557652515505493;
B[207]<=2560'd288979645446376948782250787053676613573433970721619354671151236981127051155654612681091900152609337817320080245804243963583288008309633358573434220063891169298141863684777260365975544591404126846064038574524684742344288065639713769712327454256125468121935992062892012478387913762972926729387975737975775954233864052808523962969962344275342987173326325801570471792593649340780186341307466677798721929001691901382249471881441685078509511901353222297058098983987093897491484985632311806567497859270474067493335383736774573947539285663039324757288071509907615008838494445848423801214831629486613994209088103787706270610527904408867756731932689532141450702485910174304095160167322050247526283544163523739885913465126188332584490755289035805230987262744864354186352061435958613;
B[208]<=2560'd317753487534946311211450673811336501178740668142000749471325906007583308668155569843060116207753066410580689844617308627063740443956541971191833205583084608508930536666632353460091601069110986544617238798933080515543521383874085912558385283006525077725229907907675670080648486685870647332687802115549480522615283633691680576580666535154119034186527521918711209114429612342808605626755323719154670405583934994304083592927233365588730171978363413149896513531804687293115598979982103536584115421528209954503091971352490760725248911078625146299030530164184103037062147926967081882775801678030478855948317420054906627471870285507141280959414207980072205211840668995424824289466773470267149748951763634776134929783075639173801574481080239429104468419088705498630764478638413141;
B[209]<=2560'd317753487534946311209982595594716183976852533692889864687860067747810280704524917586462861309326762004703813195715582899459322543244993610742587592176739796376817150292471483796645886801345314022984208880948044525734244852516731849382292867069807211703841372496672064443053106779724022099382643704214074653582774347487029384915337669806806377318259512341097019152848102889169611476893738795429127660186103397267830220438939977432135537300877211515693239872610501046820911807037360737081966391703985368372292311428392883313958123031360346989741680362587410878397308362842847216456392174471038596810101102828181715001501406469531565628472308199654837966091751573165320898268550198159350394348181886876070378347783586605867500014936808409792979079209227556416457151297705301;
B[210]<=2560'd317753487534946304820906196863095721359691411162635445832818251135002682591219075400115264831622535140738190654121764484758236878841507698454855227054542408534774081095729097755631209910170316665560443438341029837154093533502535486691687926421622309502085328409574856191293180093272565569145469402183897939233998661858531309315645378843836159112545565242390278046872565031236307580437001803271609446122915152055490891568849581598716441889662448898359550545549636085044844580717417834426529280577824212738516982485089583031098199140716891728239765400834157344587201616879087485422191274297596562876522295967009632411438891097924162909891482179326198848644058195195818004930539379618556827579420599151859427806376441581523205484543765763288701319477878415393508529089631573;
B[211]<=2560'd317753487534946304820906220664260045686581172212007233377605044567919655095232610825752140666375270787058827220199340651108750139254471911028184933166696195649675789263286456676502212875145979102898219523924572521050334449094524428018419035532860247058653738701806150498558323116079668317865634879295570375916493363616688418522804095330959660455159086578899042140192752593670844125193121953032203406860716186036366445805106850741311332137903203490282357573101049119809124305750436150061336943369553884578436641323087842626250353607659267172752088525894238640839842181566961173129212514072607683037148997530118171540552597793181497792163520923177584089490668253712853829950506727806425496633632186695944747278430865923236241638204599730044911970595658857301786039143454037;
B[212]<=2560'd317753487534946304820906220664260045708312784502877904963354642874947490554836252843386770692744085491694874768517753901972865991619148624032181610235341486892060822392004691867298208151617104896210370391647846473919098822231475410435862679853341438281443853705467653491569992914567349669771492699747504412023112460360477523634902761612372843261253637354609188199166421747741948485795122558692683568783857652637450164263496253705758408166404820298688202809236807812493043802665378332636012939259469742303044739178864601335868193119264720972195590990561845927914557877338119839895674439177387077381564111170760317772541364399178174838837410822417107166227556969926465171634987017753874125380129716224751060816739579654904102660347239061654401342614652295661731470093145429;
B[213]<=2560'd317753487534946304844395089911488860701948910505839135531854074237262826465370810543843036022416109970361866605461582573962712924814271881684174045776611385924293830595331525657709007616393128147947770855880367852678853519140424961698500837061819335830840499020121043063404430259692638858884993290827005561124040341560053389342556181789480008259896073672471504696733239393693570720733817030399124434725310755423014180733197871515470086986551680138109395478358582772942297890468293767197678273983520194819649371091235199354911162065911217279975074978802495140700087949364259812697226013284987067922222016434046368640902959074457673110328236513497804023520497761890981511763175658880408604848924617523260721078430739531722108270930198061374312722455772210091685221787587925;
B[214]<=2560'd317753487528639321288993855542493329567894748470228013670436266589678419718534776473588637085289086982827995142077738900464698257640735745864555664780197548410393441233719560548993367631896476572559860120015579144487220626654717440702619225588949504570612655437231576996069497307528746824121177753348617126175180475093622912002720540758889327887859298131238284725783129240897720589582731239077295012938809831243027289808539520482194689388102331730517421580862278371915275120737713039722634653376812491855065870283411785482486923701505951466897098566378117731547153663876874002259683605613209240576439344145203708377333146425621626435351753167698286840467583118457800879582810726546080172668968534694646296782764009071457654749000831601335490309380737385472162991246234965;
B[215]<=2560'd317746435123088415608060873056233879647461691594630337918283153718068934005903215028873022541615844149216952068049476716587426842962640428744350090481921638557382243245852302310963186418855755890611586293023093860030391246335499133785978351685811734957196247375624818223345779058840459532067440259048802537476309521670914823340292631873092909862537441637579339507179979432541831889870716291661151057797961914512582649888485704887167419443189100884436636996870847891364823714420627974020418091490907525768538968346615324558706727767108419018223597642283775328512879705486623158028553623892065845886229068766285591452783632060055481028810873774258102137017673605114927235681335448517553684362437245033977397067714873397627887467163411531560990797812734669039782221053252949;
B[216]<=2560'd317746460949374809223695876718010647302645154426264453457498676725077972171348150998760707991291382951926540229882765458957271869987473630411777349444189417592718688631130869171533272935608604091185271952661239965566016053903248008326799016497767422341688876153923060034723397936967055761088766569055616624068649572910264616710797805077058394490828205768111883708195897138309442352967198269487801135511481987125824614877821062807851596971053250436490292132220458169261683630819471232205847607245067925189972294180455266234339856954185308135978222301066193834460216153551367576958486929428375572664872411093944829925973614913665671991175542678444245790043218795649964707002090949715097302200398622509751741799287302688136240907306231079390883804167748815285318085974971733;
B[217]<=2560'd317753487433640381438687106292655936377567726233049000725506697465330629285878245126730620841494811414987087637511811607461268417208125988862885696425782239821821339591102645794263777361205721240886932623527820421352164417639600600343241601409693702861732114672273603901328443822033740786285724392140325304030657348741942762412951256455345466168671937793711974333871216886367167972520423687009153808437821687974344719501276438244029382615199411344529106100076171099875400346631171755639177054285560841481429864287045065966801765768755266913524395965147375429639496408147168129729752716509544760128189497221791959925264534780801831810662012826704559048564320886642832565449897664577829247529093851259619992986527836379915941570236682779700292343894037444351750785325090133;
B[218]<=2560'd317753513361231062855010033258337593438400965091796374155645766186621910720505916099077251538865969733214346337012529509896737253669670955995792394299429917999217482767858669240911993472913157882052081684758776850220384655758754416259700741826598343460467106735188346002794115347354772178941812509621888203163242546677844173682098876684885345349012894666613329537630682102205734086808859855112356286987800078289985584342811021261167501777318977183328376033385372616179234558604905615528944639287157273211380385046266016261340030658635128244445482934907154778273816681029832032360335455667923357779719831706082305162206047042220723675498769441957126891310511083421532497164413549169273997823664233137665336300088760415285282393769243290670084618986787510809559636485817669;
B[219]<=2560'd317753900762203500791669405650300090499659171021887104730574228384353512586878366574029379147478782401654763411407986549920248501722363883466245803280078716703975684723812193587500809552776888396699485518073685469831444462346690059224996138197052731743673534470150148741722829448508426892653026251991798708380288505841335885996695992426582456469786400390297575850254764594208748954283229266311869195689826721405445461583018094255999341326331120193345774475696456225325555599517034524532907794035335404731128157283639130796688592795673435810319417834517169274234011027696634268527984861965018048909981961167283839433829327691839906592430258759757630146628099444753981954277272854616833972483905170063857543714782550548882912449842546143590155603221573964650682754318808405;
B[220]<=2560'd317753487534946304820906196956433620670857168425789794063270040846701652017769724453531738360291821491403685266793418234590373798842274890490015354196256493107038258628659750616329340587569398035916452406042317049750221389987875068870100122949188143992959802954019316534425107481668094507862735770599496940651878257344216767077520218264412520175262643907821597121546985174592520021836645682781160147905668402386747707610678889779520297790370737753240801623899821176466294142174757372550380526360018383350074593270641778213969426009836965700437136585156210392040961546371579196663565023611412529536877007032027653023579145894702389516287875532139891005487527527824744174475087977430962469893889769421305476778537248442376956757905328759546295387790426703248345191960429653;
B[221]<=2560'd344834750784320143710133060200862682141366950018189261976008896771490081605139322872044652538720941162129714263788340078943467626347391695668831841211004199228198216831955914674358447746275440463255261211047362541588134527965947295551169565742335177695787439158755400462799924022112292708231943344335545714512355047647639471190950235256766375101058015504387725290253517347390662815506416684021938844047397836738691788534263153717096240700517256892493128747581199666686256004603612469174259508045160409655966280175149346438835701936177423549190826629448620328692904368063135690240578403165317901872247691089434340458225927495765552830538915274704522461198120841639534762736470946170102737575450104511751138927469074366444866775596008975460328799874473170538745330556879701;
B[222]<=2560'd344947148605397338284308736871898818975764855390588230041483256077008911515121434374652215549535348699199024953969072804776178656964560633807509520476628144408208333719801872054585330453133932006885499837695410812427906788607256882258803195622893723792404335917607507716413041289873817644217983563942139753152203139629965185863875789171864983078479424693776054757184351965773829856618360700512605402943880402454187042556135668288932856405258659997100765163023000170747541700462992643717980153048861330760523430919156979918419827977178219436868061097298798823242388467161903232954801872060832649954698848537176104114590267906541114817429290539390020086223747798168093138909071335917359784505434248787928905274670269334474018498246793235544841651578372087874144026260492869;
B[223]<=2560'd317866298684192534876895883411111818309883010885907212717722667510842571941640277807161912600611137615071003936691053438512831634053375969953628531153461021878711957807163459323787615638592705684153971978463942886727180866335555453240287829797885937860176202281633575810962797570613106683708835554045326041083337132049319297208796994610532663370773026755959248854373683675944124401359492165331430455556684125161137047296212644510339895518308131724201405152306382436223818445098638417151597499745417268823367808207740728760565373156480130093314226234524386228135497618540423910759058182622294513152629926407095093451519631769830063428141612550814345227556453703874474461668772654815618436522417062733110011342193302617245203036884820270140890872142473394088955152114606901;
B[224]<=2560'd319558491749591100255814464918723839484564017355805357056730105981304556636412406966110438320042409095602766051221902135651701573072300300676005514654836507094204436978614204553154734719452631864329058275691203531673634832694856435778229140342350659555657954825280259620029808996689203565480743974315960103560310958796605413327916804998743531760317326893091246558438831718951158834574808803183707927088417022584829031553061192006043594857828634286459305138938379590640540768600905460654591017811463325143050013479926059468205787662404959884833735397012956970437195444609425961142861116928240036087407692721388760946485150761366693058899277891207422355242479491710383574364138321560506683069534973472967757586435990458569459573408675252119298538427618552561039459298333462;
B[225]<=2560'd319551880213967345106624731377263718891089371975152602183421110093948483774549082444430329020965382200792441636413191199689953789754433649128276574779808146189069199143072707462127380622230812914204221272597237136273578392728236113088957573260373179460942503897884219791461611010605492366137801602465655111031207508662039668389607548490269096322830217151792359350057613163865986212293403145582662353719396725449475190528530245135328632729798389768259172799320899408722323959919794416336681523430951365470618654760803972621075361086475287262561076271897435161512365716041557695852323553038046322540157248305844604063344869462803922242897923418933714425277298687666746255458696530717318317787601393548511607098601322898417941419964019716720909410973256521783597792383747109;
B[226]<=2560'd346640168219941423464477829955346034493020660772893565874061069997431982315691149280420370861846522151625845347123132853513944221517901208313429728005304722751265541952525663160756734001249940883927525913628241082094896861488891034830449874208485141000083846758760318865525908114811112509104950383241285712759577523580980489736443604398594081380813979248523129217675697091452837900881193273730553394309811283549261731141612089594893120304256774098313897586276121011462980191697559437179342197584019266330425212601301551996810527034323784775537056304523536864599271749640025215667488907766388799420949977732540009354478580223127313575439400028074433077175545052656926622879692650614322103684918693320233944249643506176712265836373877502741411118641971921943015401711748130;
B[227]<=2560'd346640140779067239244690912482129374509895551909489349523181250312541859976647720316090396308476776598563861433690269136018792627657727806734290383381061697943618874538505130320524471102850133194499444014313683238254146923703419649339128372561794051425893031272286800934026824450934277881741943526257143748193489505873318041827436443404171261916844712045195380131287349617290490416463390171695930950077739754977104289558349209216843282312384222685462912662100294322794051185199166827154828600208466690398626991445927630529156398997834876693874224899372054696169182213736166416470556859612302066626673864347984080062714731409128633670780323002002672663959764440771390990547890765887583820718115452770188656303304513232378036036210199525820524347802381959296103859323487009;
B[228]<=2560'd346640166605773995400577120175475351950240313698031666749471488739164795146366890767761068194522842541184046489410612626116054951748253519243129502205524781668783827490051340218437546688243042096719044542295920287582176722628571168992069516020655067868310742575843102444994260653411768095490577146796054307292569135322466209195070355796160993104790493615971755233870860345334836450059729129028596344464864065703262903411110766133458975679825616625319163213211766117152372555870826453938377130587122135579858418383319684296272277614564436502295722400168273569049397036852418947649362112787964783762193286858382413160409145459935379642945320283221377843823072602886502861014253282097173515758402236062488109953926212004440233157504179902816894205775963801181838184362164771;
B[229]<=2560'd346640581447224898058807793793072740507155726240344191738180217225941747177515652468349893351572172027521720550372284966593755404032109702131296086973305866797806934349559891642626190863114213543624547008952028738337542644164981248017768791913635724190550754190924978359727518731785572448039835051222694186272329942844251884613774661347598793205527710217811338463657724079442122321614682480345060505354948254166888973664307283888568679531064221514440762800554996073395370143653562556427412395651992980450795368639280192223022271444890352826801552586935644935197097797481528444391983912687346511206172644303682317668160105226032724571558421151765278821077628517298984466990380633467491105892351307131022080188625976048616053671916553717757331995905945036363101806966161955;
B[230]<=2560'd346746367631374050104535634545757098546493336573428238019009521758790159691176133945053408406139428924666421182125905512590384017277091603052695089134101520721689842267219940752740056286863479084275863744886598139197619916206297373613741972468308882747849330101309682794038826351451687196154868943617089792159743671404954984048050657856635876613420881642674347451842623231369989432504175004485631456545839564919794100041038250816920468758408474070121998194954039794772801852411863744161331447353024731098128933284535626046423404230969529607262219214399710955686145490004050603495939798160056168126411679929086836376459981076084538034527800523958384359154379013495161776647682393284471119698471368736628416779251418700280941747112521557885704434018090969799426140479439395;
B[231]<=2560'd348438560798050727214549818494268200602129020593151545603816495688678818942391565334955496041169708739326811574299255193776599156366353518892181859037612668069204103306547781247382186367387092528428296334747811452979639673957241733765491541039296591991520604922075717760850493551896591202388124473018852335316079313814206597687291070585322006442470566795636383242393378423810607267432671200411762530544290369329023551146946872261681136461372073066045980664797981020611260332399400079240966698653544616028508649454495264258699102308411181713960945850883443351549830849818210172062295574155895478487469560834508374324837169333016557512568009695271038187898685806414224362130837083656766272852025948170427899872506517875952676168420762014448390178763272299702945810184684578;
B[232]<=2560'd346746395173158431446363877493715713824764440913228823546006740621325900786032161230622558371788813326266536091235484637729409306425495493839010914757911587768214489993476875436272171477685123029214958415003379387980359829128234653650461901524404419139857941372375209024945350696093749786507121452861102796641256510494364716345817334460163458165320476066657741905229417802945178248391575008747601202842085296469830207398580562325691900322178075997058584810469053768899192277974733009602949375963454379542437533194218048429740864885162846077088655957087816711317988928435263064261016056718376972620325327411759137029058115285726819266262466423095006940207359834312585729916982967070090879025570186673776499064201535404490630261660533058534676849673169462511906554414195217;
B[233]<=2560'd375526848904936542061070959929113125243271667737286424106587184340816897287884321018682404583038688497474496600670968909641825473591671096277592919903791576646957258051225206793961829304774546844670120019493760386984052185708891484277362100407589682637653277717346496146810548544009824612270058248286372098989818877841497087570824039293966533758001788895373380840000353724977572619037934065362357427638447253421253658753731621358400572408364987610715172669099995748533554132734088022356704118114523695010730775159108430492949097120704774204569264780213042785462255677950249991769570534624251839000571528975950912203019908855245059323381839549820257636986015484887620478753041468212510139495200920463923975296883195987739186756469209095346691412697819916325456925506569474;
B[234]<=2560'd375526848904936542061070959929113125243271667737286424106587183217577097276830811409139238257516951203291836064484757142687559043215647500987580016606826223074385296081427298989594665763744279236783027958726943990402912178642325174589532731208525984819564109345152335012335878394360226019080044297850670145358207469182218174440562903255075764007569151464676304564970463757146673245500652823688967332522762833562655129110319034005267381757097741286180593749127498713123369124302337052545942414450924643879649283965274951085153889757604229128833714867817210069011448216889001148191084272576286519495915764844516352728058836625466942866043382304633793982580544540505187417160108750159532144584169608083703995976705410992343453129944346456269637545599960543138908589530302242;
B[235]<=2560'd375526848904936542061070959929113125243271667737286424106587166364608517810373892650432926272866024106750870103817540589983406331161243904371592544153885203362254178399033415398741013035459189054297657797071113162856239639124156268141609397695753260015939463661983524486981713203845592121057715876933663972241280925511187378916563770147155631379817585754988556812014989252272252655773197743984844620412475057748193472091797636094259717386247891300557827244828006293541380756025014660577372947972120992726507117743228521027438555951966555828850890500126186803637324429652710848663494882406763292734255124596271882108047191485457219589401028333542609753799829499042212989946071086947336727731420291073602387718125204162892796394846400439265576559996272283867269545747154273;
B[236]<=2560'd375526848904936542061070959929113125243271667737286424106587184340817968492832258886869673310431100258640998040429416015997903057993074754280482346248922696337973779821212970557860488402507349841757119310624957708119858621097214295903699702266843323291668067703625866008239076434578836714428849002314881897016297375674406521832111652826269318714133765465357524619520004863246920096353775303352978116474151411073838229168623502355668871801861853778853879917754565443318732874302237248606364074868640440437391894170010232245528501382430270194484291125693713961352356234866533908844761976061245276713073864109834761974279956871385728780356650982452811926552159169609177036279348983214491867954869500779488148941792958295716782705573386637481986143034129943946947096034349426;
B[237]<=2560'd375526848904936542061070959923644107705512731742303203823232049672469254136235936305915870408881441797364496215658123751459240287415337224147228511381156317510458263156382430335043416499600032328796514562688409386773118000187241906447279308219007635879059696510540250491020928841366234131277684148590469514739011458788449435271516909298095720567715508399966967826171071772121370420137597293145710387137432676231215976827986551157178045497404293598957515410928540181044170042767376950664001223214396101324404114478547168935944303722705205364757155664475383831758931719874228078907702730019990059568603086398582176786257646519023734965396344817625094540880840239711761682456860503125656536071314824241783066228392963407920817223610077560527725055278096461150975991519326788;
B[238]<=2560'd375526848904936542061065225155606153640862795991279131701118668999103513027127945150200232793292397927528232038559664546697083024715379447025610833725195491180412960697295406806542588213746075533204453409409289416994395075410361372166369086339266880301548227257275540919535136028230867464189756934782589101822709985485632424413213420652174975715815845539446486876661475292543572927512279327793077888241347237409218980310167769905459517662979893027429860390277394660564310217187923862229494771793989755901938163516799975844653310305844076760150781352546058475151102564731028546353355423401661733428628892044592273682879724453322148975736695956987686856026379378924062950071669979999805597867409874475930830492311653601957653538311886358197324473101043739270403823819183139;
B[239]<=2560'd375526848904936542037483836582080028866268975550228436299778143311619006558016560733946595097244295695416156657526104402214709960678569788449602372304373203126333876510934196553254711838007589491830867943358748854804954613856315752791597049006922004796781796669782237813716727368077278028832102545794743000001630000549333573315327361710252013912280721171458629306392416220604064234680630423037612808281985670038805103337069915463406462060173759553405885143820089126510373891156857038473137758536670074976556576094943061442034994280127504671619922439288081782851013128771167609395306862821696563868110113981168567389617052184183384375925360760197876921696784544971066848403709079032532802376980676143411379482208188612990335652455712739134067247236761346319464843621532706;
B[240]<=2560'd375526848904936542036015758365459711664380839805793990750324498497261492383932042403718780954331924348499398207725062316205806947845091146586758844827770456663936173677946673000297634828208998078025408202130556652138790226120548222543092999005849299534105518538254891891506103792761431433715839547615838998417869557273573012899169746383219983638363838790302774489161716313421525830713629022209992975503409723281290193676886105811699150673185171942895590379946744255356390829115594837123396886576833946252029788336239589330068406050250345470855792060279546281128700179951127996245069234916702187968585913441026860739964247079499391001733990364986967246608137925792689987753620678465189856828226377012420656518527727303538154520726069405516664144942866714236635253182649667;
B[241]<=2560'd375414037856996234986423279732991204290631047314142076851835903593959168892061348054767653219263854623092258318270815478844302380713898963758472236421186900519131395017076807677827932339621186557555041191414956319132589406271856179910708165228087578225461237246339849303415168704156143722981745160492301932475570833299141840480114631584124005958843565516990106423094263180850202069909591222872260967278060832913837534585473662290470843665226108173731370990224456827208800063007842871614343144617037560009490882510986016918077278331468463692462692265157034250034796927931413452162318204950757069705689309585123637256186341201046642149014697652737719134256730789705575260690623609243395531005385165469875703239261259749307805061870048713350524727889289896274518525566138418;
B[242]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614622124380461241603259487782026270908880245333760961523792132117959449857122259533857685058446761548919465169024989514712398533613874737171230756027686782001497455119413036999171814375630130917216007485386761298368565355964560149939384333140213185399858955652518080017576109400628748841091811875007553059424405750788299137498186145298696496119261213504572170792061612076173465158938218688011945827998939961827694843302689917888204100760676165003058633850918635557221192133479277743977019789042122989486603468771707245588399053983992643521599186490576843575486245128928077853974945123793535955357398998895981375000083298873077323319236299178965065714700789191681360555543257841747359176685987636;
B[243]<=2560'd346640168219941423440988578396104423301481539449802853021465093237677057481490341770169542899668185228165494510238214200130854131177838460475687306015035367302581079600765322852436566792766418560816994918393087691534223884020803199982925848298410194537915174998667607576025243539516726217358353394702121031339709976418577233019387387754705472310054085902973301808985870190293251893555346474593976776471973363285817903726620716917291433392816112257225333535405205742913322119456706253779968928693446902432705976891389746890320014454358571740892989342883845176236738217605792043928921910107960537427927507355999103058618143259751981595087276179784125322939923224811091800526526701827325696151978347535134670112836714329435787295946799484590760200082760292482796657516414546;
B[244]<=2560'd346640168219941423440988578396104423301481539449802853021465093237677057481494084737407752145437816989657727544201946775909660888584263196277420567322311011164378463993401962793826185909111462371734585381543380586674414099616499268701791345407287040475115265389760129862581422728466415151001055006297904993898482580698615278852753778953155158565306449599997916693967888872718978869601499333011149074474462848517136848327086498175332635657178277184185926054068223441740061943164970404985659234664811224060035235407884093120669914400469176896686048796862162218333022573761748118679281927866087477757562120067971689717400136283079203129708795272770957051368405849783996172385493499443533996399232137170389875884623401692458420412347154575679708126450816654680846838996861764;
B[245]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678120577262328507216558830889170960411062017429977315742325748140102296565952025269758298173451307609662457239316892253008357956010901981309524699231321763160493566363708552960276293053628135015390752986947499590559639591865261317392409283085498302946279738693600482909909014733131751870608170753874164531192886354650925846202453215730970720880816365767058057208832481392587033977868236681830004619803987516130463255629144290971988899528505084492175998247173591925748425906291541246246537153417582279824737649211701654168663196856271375622283284900307861262616414624800744047840508403763636941038741012085097204283949016927637999181065601336773443197801845846422576969705874674899962128059176266771014258;
B[246]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678120577202207092384122363244393354859957961174077426843592624528780686369552787049578794974109402036775105773813043744821634662209189267653718553731705964654562810821678943016508606357582083799046190438258552788687994192528359560124341806109868253723116081168981557012534267056869958271286763882624228395069932824276320587478336458435507674037621177037922400765509738578327790640205147240564064760742051369749899853093504070928023980478872049194337506716815986629614127046609084361477134512647139247143281478726708708526709682444494101306766994214382029972433547034246192811757956345122580340894204768552474729142511448521547327932311959783838528145699737517886535736074524467092041118187737513842794836;
B[247]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124761592792981936654258000149534298776743685578558186338270770453701531871653285071117251617746249766163187269480896490586979654411262479207146885212629187275377841838186899014085678872432916561406082151351011127897300916067600298782581716155711781773442425357061993699730005819895246546540230040069242322016611521857823063205158710768559288486147679000433080183290778126588907468705880405432679969570449514825594351140806768544565409836541008650073912939803704373779495978359642365401635024435202619793467931369448540726229480339158340161416992241526471061102377705669596167963251846797833454293875148428708187126114683746125798973339741540211452282505542159291193131949783683228303140262381098267685;
B[248]<=2560'd346640168213217361001767036793235861318926445428962888816742912050459026503596158548661284612785513517658078154462401016708088993077968046411266986956965313678782596179367223357261760837883817230148473737526577354354743838206805649231495288192107985194109683551779313713705952014269452336639905635892902974325001472710644921094990975472671831186968987508984941394431507230352258339580537987167578559388963728515609109121530752819159798696653834481098075808016215481114257534582292881365225694067015105343296202985360047266946053144374333989776715723144399881758059459757203514541696045641122191967643190563229681845406141858857695773397535983016582884540270138649386227094908362691808163081220957957641102438555463493320057647940461784835440956155123457887021429509395237;
B[249]<=2560'd317865885463189880523142295052122792400353607825920095277807794088524890073498937879676361192741804417124751480357271885740877786854255052162998501851799253588048610746728661866679453653984884113869048128385741261357074654699847841474589412644917014621635965867621651735990231193162707951876754619903434759833510070972851448402769311070411860655383490812714056193507150743070206046779788576981057465177208805553131077071978249225101122490774824372612953534868699475504184235115574103416361100293055480002342096773155242824749515577167341346870056575324036419616303014831786156586847748494267308821857434824969540656850248368245074767964419968040720609617301883729823062171760849264716019318076014323593265190843998433326073592875845126272191313593155176582894269085725250;
B[250]<=2560'd317753487541645736996250682737925379915482126612520921702187059209468758938248417646943767798981289366275724915521607092738893091407762582841677087600349068637708941448363728032058593069849282667554713097397839024174385243574972749767967322915827814580037218434005264284499344805618023991698059656713722655580511533035262379220135660027206763635511278973449569830753544691880832617924223734101092984451980751853594031348135803783683398989287785262397149703889607122002552548057907917048136242297733413647380709598243816151939255466621034393092976393908450998351766358886070394775018926117589332485335411631798336973967400577474954101953246418092901350284258409832572612322357762011704778116906836894055832246007914936478010205042723776554707441251789568355167622805136225;
B[251]<=2560'd317753487534946304820906196863095726923063743680768170062177437513702521606788544526213491805190418630894751109832841492482971257229186401292355738089994048471958939027254271005835556542869894541819889533395090256047242675813776787367718528410176160352136365820006748993607147186763980934980563035201831054132241731035430427953385944381740832085875699300926530189590820302802000955886418866472215723545216231572953335201088492093484381420480812231475664550452355884427481139358841575577066775600237689167817697673959422699419535835257323794456566939321174234799516207027228709591738490910447454826794140234328855197904935627019353291709774301103545727481240476779353674050571802207564572669125573222134027393505903564031147703407567893556013033388408832381712875025076486;
B[252]<=2560'd317753487534946304820906196863095721359696716807625409912653852119802880690799373662587476914451193911069090657235558802773175249536716861414030401232827051479331585043098328861983708387681547237162220619851243703499833848121001588698698574868815668521482947101516986040194711235476494607223389168897026312520117188451888660080942948598964476933847193012112477514110831317449827631881228070828024826140830603853786552729259967072351974694874307182301665652172643862167597573106044820819081941609452060278399706047989360874155534905970288641783805043858337945112575578335276244935972738192142270713437006592724408859899041340073713947213202372323753906831222748318179649938582446356837646786443572317099552213125468266466614686873166380263841452438106302684835788971139347;
B[253]<=2560'd317753487534946304820906196863437534955801364096919006860475322615284882130558772921061936531771964149498239087358683892985132801107621303565988932806907136315936699173659033249280240823133525981680933232940087509041547891055566455797844807416673505779392854715116470402391888025124742937549293780750202619379214148375914424589305097817440426180105730277795738536672105675963274704670683133631785658504056761466813609111437977329606558397407504527625875440324752505175979994586506902159899648295210591727643951373277279131092923532911878583671566720316863038683151208494081778475430661521035477474626301803758113383321636796426274786243456071670228526147787698173306613334872531942941227998871941547141404359749675999598734249090804297051970714035999596172368411639247872;
B[254]<=2560'd317753487534946304820906196863095721359611826482727362593271270814581373189530612006778407786640614623524036636879491731074137701951110001840110117449331969682376377265516321349822966292909452521695326789777601448257490522176055609980226556020868266577542436346567130628362255274296430370478115686313391509930761546868923177347200566064993635668563510257159380220150220888228154967782892758668736001409444437172794759340885018100168542483996487137043827867253232471291193409661721204373021540176521652893145623328210484829265326091996391503420564858043004714527430875472783061079327571449836737602205183568074671635355206976406741071551942751740347445908107920231573313804134206260225859575715318793706065700426868426779395989941618764418820403795334320840927449453692210;
B[255]<=2560'd317753487434060641755263935933895307868796531313059089930187144231763934164371817129561989796683938614790182166885878142471101065892971203068214657749223324431057810301013757059473716911923396574019963457614687666403249228370821482309789919522480709426397511804535509392089910967023842643245027209655869606386647736993820500381010236694956629021739611745064116360280182854979087744184978902509717441961488198015972670143276177261186774049359643195815100197226968018953729722957974679415620587972239133221594889776149852659779830205547207992227827872720124388949037416627106204230733155117632335097877434432192115065154479196743758535169274916679600063717368394324642621971564207604498073565344585229463518056587762707153876834736600178658413332786480041350741906269995795;
B[256]<=2560'd317753487534946202194898462619753233703360157226781801623213405266558199262983318982201916308312192467711884515274402954650849681600911788892671269558688947624160616311952300110787878275071936145524861655826653338256357640526119665185905788969294804522962848504610132575852147097616828638513821089138756932435131808761503298783044285502605188652555261599433508543090052083526733211585715261997246010881563831466811632626534942983262638043171104321295821273786910741196323249555350930986435395696934440547358885790853404719436966776449326313505140214513603159410946704190837071379559624151715991949353300647868849262584847548222386471275484133997817493437191740264518537299440681985551917497087308838049904723684748564328596292818141858676524833300023960721209169011613745;
B[257]<=2560'd315948069992134110306566171017952653200152872582352403335571963721639733422862072878105258022466719086022385607464785338101195530181815128585024054453450441709179915046548598042130341875904147094789919676476551520221686997657480973017669973429498865264785104111077684962399937920984427541982556652191421250309980204428879478003039184523832463844681795149441292882822751509662997531687372923241746954110908086029894591913370972622391570348866833074468104983018145722738572916322284374505950245374984185596212384689758108775964041093343165108415183998789318664379023217707120727705831129591313633122753354258571277059399344698016746526281015759229346405459611425321474695111043085386159041137295227812197289231133170963473805805481745413634068853962932749350753881127321715;
B[258]<=2560'd317640648938520543038119868084517517824557377420521907459635320501792548689885034053218025983056347544922876349951534495809463591875530969732852019603696663676028638305090009942927721402839944540731652706185809235227954561496081439588167072894643005750060354482095381311666890724525911088253798137661423101224216584636558871415788346058860322578747677624665432740880874587317731115799805246107256898797239582087323195967300578620997892272686846148027904891071193806772707979665270658617882956121089172954114990722200913647528594459238256269123052089577235850820278227095273675754221120869562235214321509549110168294967485052841179022246610653234673433979258832471549347132598639596593591711753683698953013598060624580883802102663538416720078741371317471182282849666605329;
B[259]<=2560'd317640648938520542638894370453404480048226440710511727196753897772337056549868125820559187826078180402939622526852819024378787780626670746720939668131716435308219781089605299173362043784022211890016275587635441865529936667090792723012192292540975421048673083144242408062303625554727345328194392727825270849929470542516724228321016288569852987190144505166444184223698476351320207893434286676576029036582667034321539991612328771221669418452915945744339424574316928277517662466884599393089299676198424297263580925506721499577278522839304187310615640230434718070432569993248133075022646706327015975422298499301802563301249948009389834180965739156232430267195176485274148743223822997859446598549161936338222599939804669292153057222965737361192387898302173394937701629474189329;
B[260]<=2560'd317640648938520542640362450157960744466411970214354718679991686109502669626095932683589427949689659253161371866911967538513882402716763941640675223694047219217752622437587855730411486761041105534912382521920247227322858488637361059342928780987344905929949643532059647168841269967307293714084409164966271752363475307778117107273646096179561744738958536682847222736869622733477339246749182134750883775996060587482986141409333594593836986849399331973222119788354941298463563690817123122948339654369826681736307203212505559414996842750401362289975679469082904844484324245074694362590931238748717255318162830402690066461153946404708471841232424932969141694696776648696993766201985573709599443256928337424998845944083537381391737262923463468468544309961916108539040237814284544;
B[261]<=2560'd317746435122669694684622212694024785303861446098327880176112366031032375778795317006913245828696099607160884624684899505231830267737235391468697234972848144148376248303854337497334648950681380644977968991447831884273811966555673463470213911254298498898607490126233912958956281381448451966960286257250506777727700329534336249118534417358775988563595062324776791249004042743676828993382016718337845579639882584018324163237636701085447851822498230420984829515945017806981288636609039660075112267526224750022982793358392158758896496890434669480302512039108785664283379328646956192580730984644776827127231742798101815903825897296764273129140273876442461833290667925479076168577594154596146024518992188020476071223495883978467591851379352872619392464056390611460882734107619586;
B[262]<=2560'd317753459986460849312560956725472569092506888800918249883062862634991083163969174093271217195096721335843334880969806623357156754529479641609411789761931153319318258634991674486683656301903345059137721112144552962039608367829453151261823566700707603283610218172830254166446365316343256110070804933214335255735180100948571636889518731204288686673401071910766731876641707256784688532844218416892718204366223312698731384503266573817377934971120121651026536422691090361723874596825748083791703571581706664109805182918569269998851316754917591363772215336432033750764649842442778637998101423852697728143810485193524996717534378924091172027051314314037948615651712901313980372391334116459344051555583171207093818831445929087759148091396139735624100005849230490243760530354444051;
B[263]<=2560'd317753459986460849312560956637990987047485562195439779218219900017315703987777361350898064867256965483236729602048058731730113008879076056412011633032633159317246611694014461795018754136283181353071922724564729801050891401036120747041598603959548158197031179645510987879763193018873934680232688260078707380685442739611357615812234783566352598227142944687225602343081362019965457761602687409365228438689952964482789351474279392916411941546689405777274795728180230226493357274175921571096872690886895724867278274697298143545555459123539941351034703310452349979329371413816018465127876979546135543276598703749636433085014000399067050595629629498253150843820459708698959814318972002007879906422816845123001066793849315102733820571602562998696870892886219671496049095098058002;
B[264]<=2560'd317753487534525948292349245794709938068249858466808087292372734227895761474912745898135216077055611002415837104828962115118744433188610474897626997064593823169306585898925531106887730188413709353089954064780979547499877691830050619940766871684166005525451645815778197329614794542465214946200545434754086186804680848326934576591804295242590237633243085912725574550973414825586983666680314280941971427209708624020303831655522382098316003232308610572729801830508922321858975062638718133613990481557864091301345777251531235502677349347441056339887165860646970423341797032257295623400782526491743440368301474768895949899530094990803500107915295633829514968362260614996947320577959015037480947063301858386023620820950218843253767139988907850271204377897525890533205784333202740;
B[265]<=2560'd317753487534920032537871387421663423500086247618536283839222068791894257653588148754663485809209020426233263820413083636101253994494812841258117961721460968507375335185209177797297582487991533302604905080050048954147067143934727940374627895903327492794619976395927464580170065104162939639647166888377222210324001161791925879851943714501209422854799571734830576928994329481439722313358953279883620668263759864751925410072612236653919443632103550715041939527270090426247205519427290971393015052946631228718079090989357874748899874564172709199758086362016020705753618783663600545403099882025371061945747425299286598980535824904037597675220417023634567597174654758557892878775610590983892911129561561724585958486328216339641475859017441964374170031467526155432170630492197431;
B[266]<=2560'd288979645446376941970361744943200146659999522019908206910638247492810100740838637370338268729188677087330656798637929021678140513235706014973759812029069409711592971367387808465447127931092489062694752313907268847624446285830897836673711123412120858947424263569100658654720867866223042708730378420998022025886042342827829266536545814963746888725749657401356415135536908967296217174234150112036986982377506376055219300730793233487905288182591325081499201897511315084913665882300485795404385126621583990756757442604016050773297334317389311892891185523089636851253787250434144163863594734439724758391586784324082065864951633260840872781368521044988165509227081054367259524566157964207550846326122444771054311393266226796502154398073457186355259705058960307448737094792917042;
B[267]<=2560'd288866806849977458483858624771883918446695681130237286540045596898709761482966975056288394160891480090463410409086245711880041422386743170415642274764497860817481281934374654262979126551741319786079972786087461784827060591061555919407263787168624956202032353540836595922501943326864180680812892046297314875485101782194377708813559786924305820215019302064383659118277112541453371223870974811430694782263009645931578054737766669351204783408077398910111070025336646132854594513644192341321596899725812023994952536759426757880512940663279683269103973959881976107062402834231850989340730088228753566455499011588223840785467330130803614928891858566154689988718303982543739709501644119916953332507308292813562535153268176764505705964703579565786456984762365349713187736209735716;
B[268]<=2560'd259980153713441625715192280146656348164599996474616019081929490646689327162569073469254301450525005956137870729411630231637117791948567878911898097014100217303164312660183367662770444908517390735257569010134985375858887701452046385940321416884065362629415008839259709034441916730449783723495757426038261345414938305972166297891714063625337560104529502103077235048308413264933588794635382190455526839960285941561047521964503493359339134252897595031067565389238109288238061959544920929130552000621764200942041974164213060858468643680010600114769383766807301647142889889749141744196470552291391395156710290472892205266391979829791626220269219128371265744056151951135535021869627987875042621422236707872206990578404854879850276257464329644252135538732357382213209350640705797;
B[269]<=2560'd259980126165376424109298767177864280144426185042439714215724752053711918711988823038828305599271269428203579734470458331702872858297478260082661441469393474001022944051984282568755502114514424877434360622529178520147997265948503179578801000242269185647900833540530496935316692594342910704381353868339700113648456034013296122846261891163609185128360983732719290222590732732034518092691645467336981095706128021511501684116217290369715576768741842489727430546313228250995454058457376275811547416137805894951257033811375145942491109039678145012796083697984210322382375139216451295066371340874240892476979712690171855283720542377430455113272753899181136870431210907312957287213714770287424056501166239955759907038936249981807910134786166907755905325898890386463450800963797250;
B[270]<=2560'd259980126164957709598431109480528522976581204176389254795563441565035817826931338618664392124133212584026236796659287452535988878703415654806503388700145241893115554280579567241610919995639880050880533018289753551938009545481786074441487136754248314826441005100224360756490886516135237018309122745417541907373350104384107151558505299980478149840639637932774267077888347627602619225000516347931746651514380885766413942714056239855867581978066393645868107720602045309979725091924103037777334902050907727053230517849335300209771384900260755633586873452307201383378908629571156007042400264727321811007717921802697677062364663611311791221079466341826934190509663112343475663606406262768955543112831184362644061140789609442469517421745580827622514659047338976529262277619389504;
B[271]<=2560'd259980126164956073994873034185690092983248946030463350693357838691612958441051328836841788657584786490717533226424112379133972763299860838236471488563311602748525007094227840998225382360134904686832881951917914218928921105396264308487979163139330391234804749014820699397178295344247931241375194128524285002533464311945704956164570845518108774451041485041521502278809590394652696540763488351274870783678694094638057351489442253662710132478479909460480940092961719020665735037888569948675613912553446728536087715234553449405550707007616147573529552668926317208690969704580749901333468381438995044340830171103888578751762598381230771214355500123035737177945579983684425360911232045763835852849839293650369188560679649517775921833579231682390608486110676164272680513841399040;
B[272]<=2560'd259980126164956170206853155514029587934616895873898364354811990626711331131052158964428370481388318118433893937909464498084430128493210363925700169671043284880409469945546266981927970355232722267633814682093530345175088222956725425070080053102197143530536911884143515275885117814778746794288566984716609681977036415366544049584639499912232977079908192658236882276823779475116632324622804080515745266285632906102107835313600530665198290214207875279265614574548262579609050088834101638240256282449951713585759625074581131759121074555666050081375154969642094753964309147820516092190827397422419081805083885543824632329594255286559081241735107460869610613246075412111206895106144123120398153836890024427982054374857713175343229929211028183829895158830908138897431325842215168;
B[273]<=2560'd259980126164956170206847420833495914820547020348726212822807264190675175790277465847679504984811791608511635586367190170538005986887603135161843274936980744967375952952811934737040793123090617924864697109154202775334160105094866109057623423245899205076014033209887130099440038993547330200651981277390392011003698660313532290335662449425160422174927987867143233078352148700015593246361599502434452505176110994569943935026678591133299570392566331304397463230727819952324471741948623895868231711027849080736289100359004653004971874584088514509659247554124557408227207096999122460822418533156645384463832742229979110533875833289820056073191083859285111728730501124557114737070950907868702654518018594025959195205189395068927861719310226246090722157368044346014003549101786145;
B[274]<=2560'd259980126164956073994873057986854417310138396197753029943385654956091821258853425432927861803567324959089846284047238692576625762355076965363395941799757801441000556862999797809798332948017222410245954266706392639349847287536744708707424059534442254094393925472518897140452094254843546396706035045936606743483131214071976138645393211654038033832309685666658284099464272615730616878656040156316842743987393563797137053066878354723191324374228050421362004497692511962645905681133348885065674352659008558387894693821421757169367405243615877179504899796006939714462879696877513864892965299435563702955857377201895019899316261486579178868542895594956631654298511974677254538949590963192738541366698740056296359643063334483713074700118707810056979806222507544511480369298893200;
B[275]<=2560'd259980126164956073994873416404387771879767763498718924179914044435435987811082233252787376235672593533905217409665704182379635889975193385881660184778961904201236497117048295849963621683012689289001650374302272993790314408452973477108800311365676977124138639756634974475658162082882831194582290826543350078866779119748773379729963895509337107858220418148910064768124673551453655771469722842197174123350614446760074602544962956868046742936030777878724529283508038782522081835110364142254400939947536724199300900174003416925636660085603311705747561638615276102241990832909705989888482768560489242641806488624259988982696347174304625108810565325963803065977313443483578508925750354462286665657974234363351518834031484115238495159842920763462020177577588735245247520168940640;
B[276]<=2560'd260092937219622078712983056172480110885186913041830297681687066764691229103699959871019440887329543248914928482219920815768014839993730613984524231882602500999002176630061301599508263083264832035420612470232752178719246358447538173955741754644179749881805646035317515385595994129567459588997629609675735605719760809339727556967298606639016686475332434340848694267788558734796399658256602763689593520352686616360053575218160633148515422605056178229304628365737131147591930703833569390760988130318311765313381578621119616941072396096185716775973963205532529764377991477183491318306794406359498705484141385698811022591500306290786083472248040540403907976443507030219044038212880948207541810496768453077173724811684252375412359319497936531847067698776776491085801510757470992;
B[277]<=2560'd288866806849951192614955415625360895613953233336898727562182412852525714902641054814026216516182792430517548265082125751717977624662277627134866922233445631902652942438028721398396469397680305840634534063190102589324432893493971521678501311218259204737815714120416390766169667264423916495622795667440620097600644174156529830698699829192951861421083069171036135894500643493472441482527676445204179873011320839893279535241723020218658947537864390061216447922077560537233217256034702925533784409385610453851222328474719633429250322030001598186275948718496421190549544599180562743635293539142949259443858219814224267701276883866290616324145945197259226061592327182494089441745685263294733160963809515421883585583989681051941582603098518813463646743535331749283544521391895376;
B[278]<=2560'd290672224392763381114578964175901481970939881190232139603399573560716973981338106464013211231137045496969994212207718179939639427800762007124333830448024633465594859214291636750237158104767421702597488431095694200327268323291451430664192274714090397666774983786449859332873228551605795513522552920007431513144197577004177773230600410105317843667617322417382930946415512105102705249204953355019820447634385979299096925306482739288523027092590782233354964768123091616844851086388976997347857899850440910475554232879589132402481644664803882275039678846180647008043835420217106147127160923039953232452806577566371501296284157612253274300852718498827585410781853707847076865990300784423193085047646391237994430722281010246461581049831895674162333474757556846988297704876194821;
B[279]<=2560'd317753487534946304820906196868929340066634276223634716905255145780776909679364960328608483517924459312074692188690964088776759290567131318327241465722876867435289462235418244624663542824719625723186667995182527045578898192552483143875733410173386853694083345118223364375487126753002149545584957962460846518977647399780734397124486382466318801168342874725174148487729458336743059851932152689271354019035519211200985445126126795974848775888861274846207330344212246224079499206530504147475114072391443252499250506356955771189448149264900794352331059558122771834987866048417287040277781078595559936933790130428293050658776020921083302548041185128218769032860031200110193334163851968339581509856762525229612601069310853293049767745787239286735436361939832114215075882812466688;
B[280]<=2560'd317753487534946304820906196868929340066634276223634716905255145780776909679364960328608483517924459312074692188690964088776759290567131318327241465722876867435289462235418244624663542824719625723186667971607344862000944512445037011847498094451764098803773510197305647386493805548129811935976402306517843613858446966056512719615342716959063443849667882784004123509082125042560032105097063045991356934863950369224972217543291943724398280603727004471444282188510069315834591044476322860867923554433690568529845116034788217711182793553707210338115266248778565344585613440524906265116284862774295606351355259534913167143613561720931857597570820524295245773872195401729103333775850295514418466259932738014075809025682897743954216714780321089653617535768852791131743749906243699;
B[281]<=2560'd317753928310713586540298462664295929299889208391024408555736939218561786004688350639338032633197773579088244755610302098701786443849174148961725784110667209816716310082271999654957951291618028835850553883881281945489965153134911362793105091560098096585570933053488678905742460211877363664200921839936662449056414479612522335570650244605896409881376619519704251701637747599877015012010653918531827489460329719059094566710859879384070221752965437194010537774639525451328462781394785862521023684554514929210866229068041954890539580685776240107831884727121461998238280586761465913532107640023868510748285574274412231685823938048737738506330585770436244823700569518588081474943538075466763073390081475988291307621926083554650328098870878084306002697017373620777302517774360875;
B[282]<=2560'd346640168219941423439422628391713984263886703685131535420443822611832605293037333574037244518787172703775968942732286651639363198996520056094789732631319330240838777887360463577840927552306084478136068263117900069369054983563132136956737393934329106134026571688066644906031380335181623018587968642600533409945063710476427440871124385707217012377501075567700001674975824023294806620316769763374931925913939898111832312189827625966718240063741537905418750462320996426506588565801821599782695274859803299925202479424087227951494752831457677702004270028094034319995835677308599377152937671078686950196256527157081787937237864013624703552937319638923724680287671928776348631462499712500464842366294963062226971376517690816888673834349004819565948713418750840367049745461834499;
B[283]<=2560'd346640168219941423440982461496531257694782913037625399236413697344452265115959338427353673822990720667709456007610797439275785516251183123645926678225799734802090037117328540162575567999985994372592813821206334863640163545790481358472597148663889714342565014457780067275451999339793385267121747458811582603295044260782181902415610072144762570657968365571780525325371920205391114688339355854183464382774139458752720667987704886010151594880972095853417055978717421171840798207933968909058328585340225752424783033958217829955301581159019745085788702299214308135291925634520081350589080965249423159753203710218961853293558970649706675185664760586643848738128852348622239625686007798795845351828997686766735321610103824074697369307187195090153892031344163369114513382953993568;
B[284]<=2560'd346640168219941423440988578395762609705371605950116401753755397320906330115331328812468852386497868685624766778922666786709881353568246333605622878032792873659343429094883184064956013034323219323755819050201102844867563707125677432883157647597667742964348484450226273075338668700261586353095426271219128986149406158602143599030554098052790764813931780368753178803596221189551130616536499591693990183518732567007962233470986668899580553109853273854755830141732373906956832042161917561388007397070944211277769507639723699826875282710183835788746902162017531213276422055838519602482695190468681112507180757064229433149017720913792438233894689142236943709788602881604920477548709989357791542016399599173856094942447415064997504468497554059086003157489412683246773099425903623;
B[285]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197362591554881626737867273962924929099675963525137915904091778949339104316394217713016843603161012374287360889466219408083750848241898797769930648045743045688749525373783608158308119784151720703111636031376670383939478583652322970557734487404089330385032090814126635783115460588062314504985543649541832471850787751101818687191248752137759357245262119242621515800739553994723763745103453538351256988045755637990575285824607511439477695053408861658072710610089665782839379731294171936184197313158421152689964330077542462004594933484066689598894281021960037161728;
B[286]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197019365148533380923415399582536168996432636888872647018924890449265517180842278172079195175177564219023604688307968133883547182986598235390410962638849613276383369464554996690600726690625958888063621426488205360857307952727879295589043663636094335509557576978151328542804877480804550043287128126456463886364415909023073166305848453548668900837022857861510841706481633672438188901520231856076096795305886257304483700498980040395647403812559147564816865900422282628884677909332841620615173837260693822715099451849768151191986993463027117038308062628083869484883;
B[287]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197019365148533380923396865922779648780827158177900795221967848453454095044652718310837480068906341835080797981119534969397998097201822062436691818130815719659428946912125200058318188757318161271213497263277666818431513922056198384100998589627928675559298921429490833833759859091091051251378766873333807556879764034746324119223566778838556125330665271742425432059204353359740318031927021163245927668891323102168336762730048359012805140679763234696372874268439444158818622254779211647364262039251705589127138790164461383717334120704462470224538983381369794081331;
B[288]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197341145121396147756073074618384712962353541362160115379758921011107620259795752909733521878946468545593690074329803821600848644772588571801200460873054173121945272103438669735448550600063702905837710934898054218254626575664706038185238229638692723675359721813658874286310746074688566395670291757670390136084846292270415057288177384623039544356628270953596698030985450138460918215067271619280992308508283332513552427057875712527701897800954437199123569818050044029174134720165811193804399082423322595795507514201293442967115911505054663821496187703989896762195;
B[289]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567115068384724008197341145140575417786714599088588459881198745802674115218212809520185255283991666562891630378244191811411741567859792796487826428493357602975774110696588719541770283403971034353807790413525065197270707038601780639559522928281651864165047083526968260332548569147714273205664037512803235394055129903564287178607991381183247203955755344790264580523563587829939980397009125105844560961057896178527173737017601890941056727495665530046658263942385482003104244962821572437168296781581575772921736363793776659038763412294922391915056753446105094139528264159425735053890;
B[290]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567090432925311266873429198564184566096113238979985496340959643469194952133656835746548316138577005497995757447624029654308311456576051934771169379826663669214958456134421510898623358404159205096585273386580881643479678445821050156363553394595049845864962427699643404045756369353647048344760331500762640750764696974867641798887922823301646396518837505786188359727360267637473236231269425144112677475650330472705062792495713522731141693158638161778052446667317006607003796799194948026066385698883875399815766067624520126243241569723175041437100823052760626742620624981840818713891;
B[291]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719361317906850676857186335228829570195375771814607004827685064761220419558855611127487821085602613746027010565808752893009244212356400015098187109763188538122064581577551681723477911437147567632007399946644908171260143712932904086865109060750256954187389964669495484615346655876665070728800098965185522993397113894827930072338236235353101005280220356432262028282837607759869857393558032689049195665062376136702228990564420366385418878855914905129624062963932643900283869960324640033615991511364553062140433911668266562788207455870012469273645617613168373360154839089381743201;
B[292]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355655711332078306453572195590646943291720107179993066068724984637541280959265064180088169580435896105017360440926786073362041534912615781448683346753256480856693681614299552195914362667828769168502589819044592880369407939574046603673720852225995410400087173038068091334293110258998506772447658063812953951482907861254841026745130712090255280097099269561971040529673781860699776711770747820339146312390095103883599887263345545596249258848963859255882948085046190661897272141970501529732208812963913353872487086947399099769424727190003754996787563425912929704816280863136336;
B[293]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988033723812451869009156094733522140718190100808646514905608457038366627437579074121054161720255725945152036117306675986884068016537369799582071908641823013201065431465822537161864492778441632426042511114336149725287116921658572547479176607075403372981756554799675872465308436121353182783497684392828491159133464155090449407436781484079974408751881368376933452404756439532623068281376398274312218228645143655777014419888014808480585474863871632472053983025309489201045201841507930735300784585636028045445723305539480368582042644124394833211744;
B[294]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988033723811342844742784020489969899972921540445613474233240690772195962718896772977547046863523033584789382928892767766850314628785929674404824344692635015135388053920364090043372953508031962942816478692681817232488391462858236316093160488243009646956388004164317028083265596224514403745006759953642476230649539774109110401360154605175670079745003529510390024660111326181405694828715331843304246953556836217601954457558701481908031807775139288973839231070076954169808451972976994233086393583915905330987382181445076540217655618851711720169620;
B[295]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361567113522630407914624097528568898781818282409608550189385854914226322757036883144472999169736565565374177767311700895881826058055960241032737565718070602840518511249993430048883288844839401628995704996137111100247093717804718233705301091297772828572763196710172702223807710480668597771342115070222664303155947597686049990045383630627416672344578057258956178768399132881870867357832493131160636666325617778399339587073950719366133781685719814827886831011076685539247335550845226580094999253625183532842163693926507287183272171426947915689750088375673994486014372961287273117253667;
B[296]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988033723811342844676938225318322563983949762419353146375418041336479980914823331964498796548988979695926205626186669190805361543770292055247912831334056263807916268903556286990403116539378021661026464664009037191133942514672152337519459981276439366477255760944102021711328593899538394494688879996985840973108105023157249274400680990752629129135406146194466736650374459305348691251333539133824365787067414565893370582197011984981960840092054784787244686465907604014855246959090931463279634185814240356352333344738461102165609590011684071834640;
B[297]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361560783658706004732103664600641902542363614354181395244446888154755421268355708871753778087647534500447196635385152543943035721006511517283719605503739652108695175426456644964600192817048457967132518885274252790795059133437497404314402144815968255137856776960644583898048330473462768708341178880132399706986127033702672026717383626829536338836730706681906828056711754067859792134772375719104831641593604527677338648424059723702534308676709374591345222354276153144228513180428613578634103679665966716600404504119831680819700580213870619223729593097227321127126893659670989200661760;
B[298]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122895352988032565457608061109689092121611278952783333352473830933268703877854987356195931216772786368020973601662204468982178485966163616183979992319212899039155925833747184486191129662370762517315788495734495413869557281528970448298193524963297280141848922494511046853993819237012027091717187763381776133755902794296058154620576389927442176484306688650685329487365172965461599922277689867759264837684299890746672735226613137922952041454279315886419437134296518293426067735129401650991652067058662147872596444867510887932290943267169333678927932688720;
B[299]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361472119191134877369619651720082072433661069698730235089954246520197486904000888303912417684165433164939353047149554433814553218754744984168673558277585283658366058778479369824793097472888332731472498722030014843811773032285889152482778224747501862128377284143164753762102419962396509620922735359843059256863829530129003807696518372266492201905732425800551317227598747286244718275662569052835658093432627271170267666524052995797656137074628056069543277033179598341376199038918974621865930559742851191644909924419812137541568310578926706107394255951904747761296545865782473961718306;
B[300]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361471748210099014912036036603426930469372213584700595561729178296067989915979080709075952327491666053434314810378149440013610511648122733910035992161340201941985899453457009173919721915735540252066399711494932561126142789474638477854623892319304822078569855136602618896228721631340144792659520190588165540119635389958662017085643689623762598112441871940883288245529036757506501907548011656460587503326307349929911813209373791173597276108298757602273733522362329300510952158097014037008769942295789883759166206031767110784886821633631361545302678783865084581152832364396967673283873;
B[301]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361566719355279804053441506467122815751525225115196377771817401757367386462545557131520677961447685129326677368151404776737059354397667643404877592809114649074442525575662981111239553066246250667941330975492914250537080996991535703616572387840285703802376212346012914613614871649680147836618826303580533098789011768007865678018960087464709126163338629517337402105292457125661347685383970824961738856426907963052918389158077549250887826069631673437388002077992143102017026415460631640531025746767244374721140549838208072983249781327026641768185848005457776935065685418940179073798400;
B[302]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361560783658706004732103664516866771136115692876234950417220619484370766225027487859616341239196425107187235702540821783357248581152717226859686311092110525413330905466511127920764159586261121626658642267230488709245235769380713499800405692267002702624978601424893633491566048866366946632190767071902917533615222837409809014404031244738303137786889182164041928233566223157298924763596218499336322892198803931583956625910957610352571773929706381150873364744087426744276789308405299256463760729518138411942769218244801587630204408060972203892236380767852932963066947678973560565795680;
B[303]<=2560'd346640168219941423440988578396104423301481539449802853021465093237678124762614623098873599494763007500281967296513687335419392088496674814376081848979566742051237292981728892641329721887516361560783658706004732103664516866771136044244596062906033682082908235903977857626100058876769565067129089828776698737264805814103992565373953941406450368175156327099048422447861590507062070007094951789836402892901584933122724462002760073283123522461521082138350714332404817085686391090032895411750075728280729315343797166470717099819676995435337186377414803993606541870382109135525092997983299438821011816694689345685553718008582662630045507702317602302293455912535560669663963950188088557173207995071106210038776706453322280845856794167114858295096250550409360056836327586137275204;
B[304]<=2560'd346640168219941423440988578396104423301476545977474942047666673634590095409136184463660586387126194780246636445516679603967610207560672873785916196666363008166769277468239815958546324920157064463275809525456367551085255673218288991056542706930780358153998691145864962239433537024176590794849114601394414961273582518788590237812900424314098644045747216037911053795972470637489915993458715780659665630785427358729580861737549040016196529181562310921552268696969699109413161167436128314880793760352994910246707195645703683596781662600625463578807210441384367489617548974468450550442831253184846810568135322109935191202192455973168279487299908313444567416785681821096634127638719451873323647619915869679719377414140818878546460044048181075329917483535130146821221300943950610;
B[305]<=2560'd346640168219941423440988578396104423301476233885454447611804272409397093574543782048959773067898893985244428267329366620751873840002172752499030843396787774798990026498646748665872362609697108394310587915809637182933929957618467092833318931116999413025187535756542447361583603182505421850593618100447626069436848537699991238859553453831410777508602466224608986322508470091390438126348238345385454579123149626474140860377789584109506605560713862235206204321695876113495570544903790791668233674975232706640862444146310011791439300757361247731279911049936261890847625214414467133763594149182408613276852780566012572806772566744882426227183614488692786453661177173973285397070344533017113730068274113416568398449667460472563848779849779093252784573659508191823754930306756786;
B[306]<=2560'd346640168219941423440988578396104423301476233885435917859629898776014542718662163974169951624181541902443423122670810929418712654957331650611398627065077062109327828315163968085058295367362701852356089860355057936862836421467850794459404923637988904120142502179043904925562410103945598319055838918758832398484075849311363765447621933487090547458033587801087019561886842998657534468881291716551304032785450875424149455326032636318754532593244841867509788394047640801814037676885238700905014253004490561843540767312913261196403048715014390758612535070888179909687563317568074997505683259729600054116549454076079042161881904177564144635418742264181085577238797739929362888863756746530018196927307834257500477520716457309882706192850308354758797682640146319985894696085915009;
B[307]<=2560'd346640168219941423440988578396104423301396649205842767723611819493854373822104010099445408180586885318458673093912730785476923093888963435168478451464348059109250797993301760824542428419595475719635686892365812945570017049961590265590113907814250719162107828945168729983219896928275918865678453227043657955167915547766764008851622427610672695766838077293918661834882596097545269939075241638473624495834837327353782998189253733416445362776014840040409657280523120832101861294012136795788102552296927645442299989202470473220308011547427936921082815015417259376541485657631717544431264029585063961338938012248319030149533980867092568572025203086483922197027632716756050283571843052944623886907587211775828858597193390174764954094570158513252629581885068038837731820733417813;
B[308]<=2560'd346640168219521066937486828891007452419661995294553834554343263970979204877566674004431222817267624088614193523866229107771663641699394886204303022911086858950399054712054270089686697782401570888860626141158726520363299680170394762978744419816718018015001165756910607262824732429972149902450198250171800200014175124136079597461831284781144630295994464889957238368783941544453523730119382841824038158361924595730736008150092369387180990529346588532695512372743940126513769814368385484476568819446594881925453656551491373048405033971786398038037997909650582708964284268563605654954235633954412824979880320429115776126638843442952534865062259994922665147855130375855545648564344791459991383354597568599291195092333588936944019885105690579152263627351293967984240166440338582;
B[309]<=2560'd346640168219521066937486828891007452418388640421083120239808296147893560470781439972598720736711895770266461054962436559098567128784388792957115218916868022914584338409332822952081567126488360933246101423450628970136321734326417988318303924012248881206349120721810242987680869224453238912744365321040200173257657219119724292562757546930784219863923073256901427597502804326738259990325304481012616531941412011285328414314945647997709497822282622642225351572402245977239553920265804666312994735933515254255226025815063241848740171809139791627720176815900253831562519585030031663187902627786264022839372931490296015568546813453032069037144739634440164924197116078659885798235476829678300766501674613732633074355049957095153283083700975344959111715589913177854266913977282582;
B[310]<=2560'd317753487534946304820906198356137509167880937792738419593881201049396137117862720919147420191031579819409021540807078298533830516174747661319350035741409823384720883255311605077732380988068437898163912476905733304362515587890645904925545223720790208117626145173187623913257168279933671294615311818488909499210010628059676860892876562935188343120114350507574542375921393833294115763255887512631391548840967592061515132680664244251878024378059526057127979086134092900220300458009127724495933017554948327459848559708036638209322549717168723799846284202733384793972992338026841891089028540998026089451479590274826368750761483326274079006919876176619199968688913526013572140337049006550727648883355720123273484335652539079434955602469271767161666939988813481459189495696527372;
B[311]<=2560'd317753487534946304820906198356137509167880937792738496499590909143089375243973557712914858414797008282643303056300045936901180062108771660033239134295520925397067246320131267745424130705747144599464653005281406660103303061045290446519820935260452357789498917292113822318721080400050271306597000641473773371163937411352194984604356667400243160120382429751157688449000563948601019205122257552488917679900184739614387216320151486782036256450958072279758167237786282164835457085714945120569891996443424862045189357233463786242213928123178938561524193897057293130924222723343745317016627432715997557978914459928547613061948937138241886078200471695577042861232179904104655219973099623832156619450996476547942577577030662221669056628038625048884059189664621453489213157420826627;
B[312]<=2560'd317753487534946304820906196863095721359691411162319286742949858890394108415278665140259409260106879799984137078447975278439948296524640158416172979440692254031328790661889818655007572683860927852732375037564532471543210805175835612471763013879223981972852844224093731834187908419199124840675928042190371093873093955829231759013865622220231390316553063246586072572632076109782875322950556360640175304206736804738280649748461258378292685769326486379794835388458186562256841334116822001424405107961019924785649011228442693928859575484544730607603120409537597555371535865130116860820266473150794798353785340275557927665112191698261147642067436238357436872083243642464398095078085938959850548104331890483011730484033441664584836481294942064620606714242349358945444857336173568;
B[313]<=2560'd317753487534946304820906196863095721359691411162319281936343002134539352237345174649307257866305351539473040538043324838102283940237970873673350236521254975182907198340719861905024505141583602191998927495188960745296500184896814224479192746182807573720570999867471351345819229151793616133602142352266560162741710522090871864461361893599945972495612391118775145150600010395578104227115147124579472082297329600022727007264975243275867219672370899508013852532960136623344368301784355534784749752485083610190169137750665217206882264331929146038706620361299772920517777869574430441028973422974499279743176224748427359718370426660230703108045230082564920563829105284004609622256231068040411935356495170723835665469070658470733821220975874714999193653004233958915747406194034816;
B[314]<=2560'd317753487534946304820906196863095721359691411162337811688586404473928929542049364674719962046925866062158345006912361807641648590285380535046300098290214365926248933854634450555042143128561353092978839462262967514988185461265498750412136506452484447112214135921674747613618810241039407254269078290079356060492190081029745766475895672509489061099490009755608968162364479604338848350450854769016463970423429195475607311625164058241276971137425773463121142629779542429871510756299682900166080740450785772396549146815276246630498436315854967833664395030073367782636732801220697269259626326081553557998490413133437110275707224057795117065128104156963238009614616466354160336556357598468899431551061706564337111764749713210116900346682734515825351248387607637901868895878273458;
B[315]<=2560'd317753487534946304820906196863095721359691411162319281936343002134554353030447196958756435477478828486417709489131245412842725395571445905669536450740998830845736507297197974926460774460928955251915402986280433702067083623286281857393283127465235485095425444191669856949079435817375733724230390758181737212437707425345895827536777267516136526689573209512901528558898563274774638833951658753781327015979237195649101754637897823033244784146827017595628758774540169649159292335450769911375954819272772565484031576809597547646997359305222515924789216583270394897640268937320141245155046284646104783484542554551072454524778964494221601556185132399464351944863347002218041354305113417749262251600112517024135292271693814632790984354746038446572392031309828083541734907922360161;
B[316]<=2560'd317753487534946304820906196863095721359691411162319359143570385691210437903831214442527082243226087252498428349983738811388816586924090578385145421950890884966004658377752863935981211471875025795196975970614364721968920466944714308844910251445802152123788797315528107047314002956132053142252846998952384352254595868999514823982215432998528034886796556398493057563935606114992810880478978986721056386920585268134442673600755084459524516371885240598266175748821240348588256393691803201048456646508230365008829234858411733580549702744322512491481422783441624726380463432665906122722253602585196646162220338994134187928818026318785430261533059529388663747569241525029138040719490393222294425777153941781211982198054657176257243836465378591911063212214068660119689021334029120;
B[317]<=2560'd346753005094586844653826697597391563598151235904907097363227980012941001124239606847938592268058878585857298796588960848610858188262093228490339484436098246439993522127358126573679451880958743945236707966628198317736393925715119433229087070690455613259520652125038012279235135046519542372751722698394883380935759048457509059258936530600204160388863753251521673012673035543347755619200069027790754867524427095642595881731575449198279609805323406555085842961747819686733575940879581236162129204546000106314606061181132407296386832039677308617446461854833135049224521873186429364532436798849807396335268766101386354142019638613092042423102397705834342871677256695787541784686847663460432509073133545950645320756967017491735412967158404386144245824332613406530428735353520131;
B[318]<=2560'd231093417931475595679102140442529344206006919365358596121294925400655587452840865083241317940322326643560833456576617428573562604815717013082492163434828768933257771512959445468244907764672998020647676366064855139036956061209739604127717276590098190872806053396042847365389542237537014132301271253675135907570995359627716883754346863108231834853893087650665672643048073514670476473218115450728627211397923809324511902873912530364138328534989805052991437794499170327543490783452689064711873596384016786069482858035837052764690456642728814753295582311589579063668653120855720238416095535743693112657851658939952865129897836411342967866165926524163588927378295696781029848993968938264082842617840761895250253170361098707596782358432303792701318048335949542774656188308205654;
B[319]<=2560'd259867287669442144511845552963585485560224362507544774272171196301984889656281358443266020446113497104946470155168342713810890102580836042027392181678883752798239196244989427099856354622506742720630149461627251811174181763413536364312057294706728530473344857952822686207977227976742682745185750752370103068627543993351278004238705767307367112014278329689949902565759825164472980466475446707523990584859027697715545148617954537456357365883623261557780814922193240270928055176932746976885752211491439276768536697567324855579550205610353666070333754718544885245443215474514537665961354933871925121228916415756813398496787171403460265799014880994583896716431548379883848409705362721607757381661917802188636239736412742001918974871258472713376593439418801258727437192520610384;
B[320]<=2560'd346640166498161082471717000794529672579508242939218004648311389288871180857044501804912631419446898317683142923536394151754308368700594813111993903628412523313298937902475599875639539400037587553728189659831804345794205813256671187704070980709845529374464181289282214844282313168508345851166126124449666918887809110938630931405865326718106316713081553555226872013642030241590359134486128736610088889755999675371800901366124169582526307232320216864439000934652196394459599436164080264816582759124433673427924522057408388292074967572893962292733507391388616930360267162528931578432167715713536184161924383371362030800325784290232097629697130675907374833473728643560722868932542966880927391591891018988367711670475739340368612014281047820778029429160379192554515271019733089;
B[321]<=2560'd316060906873505235576900002012374009654430029806836164883902325789641940985008568936362585226680291753146872962659636110852745830064426494560500201557492681022745045154315160785093182122340253665297814780498118716342831275220917123028994443684648727648013241632433607816491306545058813873955303001371719493524387239996243188426609986533047580977422264228971841332203427495894102902690901417039223209369178959623979959565663701148852856905648029554108233503159644719963444088012215932159724698459327359918179601534322497576069628594841179853790855927457462793739536367279855691393845301540576007967702761172173433240203613442483894395099924469696756024437412882578832276748823326753811714765341561983751008288231307474615719104083696467727955852686269682513806805342712584;
B[322]<=2560'd317753487534946202194800592138713702222860203769311019687932674225898274078150484777729149509836634348723979210629667441997355725378176949974953394673786798620188803274780146425670198966079184939429622090877987097928098654682177166796675779968343636688225185417417679737038879733532477427084830566429105681811199386440000306637485434141472092235197150054350452323880977991935128985880944152604401767722419764498252102098517347109985558518166989303087189791917424550564042704434891158923052275812690285012824759395986059632126390624197766270893545670627387223915077487756093525614558710573311041310009338831952220740670441431925926296381276246635087045930130344914996311809580193313251475412709730100724377445742612913969499498112883168162111603630806737202952365322313737;
B[323]<=2560'd317753487534946304820906196863095721359691411162299521692808698211844142165704747327457866260690525845810512854482285598332150893651466575461643165168172885286936290018955742748673360289773612238662816795482986251570056681338626225112436041683696748586560996323398173213980754654131109469608322263194036421471714857992264883696199827736077584647230694943935602065082677920414269004224011506288520373136358211018373051566981685740102726013533998078133903967200845683957712467523460760274895362811617300800482784686039508470279269298607503083335351305728667756925090581870290040554969397116458318812889261403833184964849126772799017647821679259113615400538754894219984063576437592157644365606336008712669414183973265117876186446013741874234745248986592897276820096355009024;
B[324]<=2560'd317753487534946304820906196863095721359606520837421234616955818919699407821542277576063890415250723739267907519043404134341220388916003493072607520587931836604232604177612489074669217564535600554636319881252071484653095007028167871902083870222809484691467307977868176561134659228640019569619750494415553674664427354701901757438189369495563301037831879437070554808386395170878399913291132339651349404153406958721516768505442505403114255194832200593686136949343709852599331368687082682835048920764731512081786809471123209327446216437040282757044412512599277710718263986035704258077598509334796523677323722737955957494944471257784321917338108529286638409433032290944981820850836365228025334584260737032230318635751072422169796877493419815936519839361963449839869614638040354;
B[325]<=2560'd317753487534946304819340246765367383011010734416601004832727433169148998644722141255619196684211293433400999317532303199999766015281105126695530202733684075604115973730634790684988330577008530827521005762088171090838800041863350391726772437668961367661179723107836496469381390502396553409723935971996408197474005114412782897669721324891968886899801130785323508315943329596306950583767950411954719353217819911428214703289767205738633659555041695742506199557723362650573131204367405898751719957145069622968527146211586051184908412924522510745702019323828125881311750515017693837336308901320933907636166818089362515812601031407589794891845102932586661521980216518751927380206215904172313921016471389310749843881248442845718095645789788374556521166570136986076397933609421251;
B[326]<=2560'd317753487534946304820906196770099635644715503680958773701458687331100384401745602052369610171522703377693847481147548436363462179474006518011806371627714621130231804135740790535951467124870270722179543340259139781983623606815201358724096997680135722110395925179107302603812335473348090824301464679160714904018122806219084184394485341915287490049031400994358928505045094433581712438733620094603853987436240301877771714530526859688315749652949641890493580554656236636513258626921757602522692543284974864587717523993535531781104199262621905011434025885646081254092578822037767957184834389121040445504707660432684527689567188388550389024994303275434959421903445599305151923154217787890208509749489203910345987660969135760053652600777615369548080874967302829355271617498843044;
B[327]<=2560'd346640168213215821585127764456826877489414210721824209849586109835455313546501680703169052663209646119895333878137546346647805130801090475564189204803553430591592770859444654007306586213979687320490848680657460830051961619505754115776634389734804572056413714584981072644570540096402927243219089231375709581330985531285024095629726941650346124815461439308016201634835203295236228335999987742160408286635219706831373254442746404763337087919048592636696238581748503195464988928799870322422455601539012408003692190037668616756043208441296550463861958725893004081296028396150006920022106381606193361149505399911636334636142738456530639149309998517601228763258806680894748368684095808679751501729342892752839245907391145452562297632952389415109202359956706419712781976850177108;
B[328]<=2560'd231086420723781065643201911444655533564470654863477574985537838353957045725937738658815310599045626852227729000917899369618059868742479373791775602494602042549365542783211048644963533242978644570001898606588875098410875919024959967876170108530263189830985331062482995470278099260064878453689358331020383903370718493350084909021430433360782889284327605992687442152758372753164985907766558214216717151736738239377564326244172719722795245731407247186217024528052245010418215613686013774220768494468823165246551929606780416759157697285795025531993053385468394198428751548421432149195825437196989457406198233141188495868498889967772329010402968689815094527663799861982587024677517758661834606785164574481966609348952991557979146462090932278689759734196489440984693910712390976;
B[329]<=2560'd288753527585369407195769726124550542439999628249837264713404757724042527558586706768271305316842535069601800923827830416680784834497829935771821498716589242418749937517994671403256840367607801817666072335039899222612685502614376622259733996024803498871005444980781016893382399007732680595998303526918734340398862378337657355294608028786069605754784878000065825838688187583780231826917819133792872176149976490813075819631801953464574298462537503633542404212466917452539642780070099739929840249503509620229742596917118676798445895951380023858024245724596780562475915550111835209735783443793531985601698439941046518619089603478077626900350635510654402463832926344451534092960369246236660752507851890122306905407633280080761837284178593611145203193946774499134517004481070144;
B[330]<=2560'd290679275083259650281787114505612290569079038576859906521698813939167426988689902381115682157174849164641686544129393642409252505831402999812323476107178095174356122171327338987297624107374689130460143520532470060292729398485002904308385374948057648354832199930145654005082662896407661949336112879995697324829711196087299696578036371095397789367998718526161235233636342052956600819473080793123411461500724917050292567957791222865861992292536503240327724027824081962632793393419746881111905316450656715525190935835543805143658383279102634537342898150572585538373760624913728138688566223528519978775296599018911771069379178593321256163949736848961321276085379968133797340411773074922794773282301320896982013556600597870488488164223709451870384718677038523219045811080421655;
B[331]<=2560'd204125461810830363726467229145894952856291385198917209030715662464308586860361016220423983644386079737760982832182884909367068519391258345758515773239287004638903498382513387070655136805792909986483480584047668137786569324431281254677473187128846801129585781064321840686623334238687451964253646245654002265388099908430659705981110332494215593869230522306436173031853358777886860999313545491784475581434391495480523531495759163700555373121047737555108731877922983745457192493349792671704247672055009652889831518162440118341704061761172716244183070608131867491965149265273823812128440286080211305995428465954437625351013242433359043711946445385335657879516522080749484654106553674196279977219909919407926058919896818272980607899888049773481181169691106252811139356918710594;
B[332]<=2560'd258174710451561757228305814672544198989774941598061420117678239462066502414607223486599620771967923930413876905895402524554887156195295200326142642401596048847949608112538986346481743393889050781301588506241138393747020705603305134340800792523040053959644601255270111541157082677092446628386074039595328771320738954870438928716115877395761678493696043980644613473604071597469062933351462180261651878361541728731437204470043610894402118980988020430991327147830422078917148579206807938175472698064960586593802032020859443331964286768630876179310305149996772648881318590005706429155240444957656519342323773171022201873251437176346845991085872542928589920948592116783428077502155855119929614292115911206579389936150766650782780228327728411413260511180719224737608827121186596;
B[333]<=2560'd231093445473657249464126085919728956506363447855719606176333774641554059281114916530009899827836766136798505119197077930797165863243874384568634479812999564012073947603803268357140926305631703427008953523111049889578600862721304953738722077059467403261324465282835658903743632398906498163549640938361575997140841938363654292388287211523022730255751517309139185679543290740200883595038780077087071037193357396731867893299324685231370554156966950663458292771740226981877539945576587708124402100343823487458642302642242029728309907380876077662282152065372209933053324835337495368030928896948508800293913933293553306592182809782980485838945751333751587208232297061183807701350833344534182066375780488988790859732895406533165464100555137682534310723207484940002228222931661671;
B[334]<=2560'd231206282354606370198558490021580844954873209302937098685159385930698115721620017818407014904027675990207051251359470369028149957125090745648965183314068125917614895248559831148161557151802170792522951555414181014093840975291480260955720343222586739693990438463636586295002152525651743314816019547801712992793531194880980550102150600068105323640593539811218472379283904992479149836931458661326488448931736041778292620382657004672656164425286999112045027151643116854701894575539477340334439674354347141137900413472049134866698809486790366011412996570313949132144728597437789932640529113382263959358735150489901901665105661010802350663526074165571009305494317274034463843023224037894299453368824347865329955755883624226824962672611201359421297373039930626178851329284846178;
B[335]<=2560'd287061389300832008156039550176997572852029856850443528706494468340284052229061628375803826150440325514823949974968303905408899783413429293201898188948312288894467045836633529166220819949818312212828509139507614842392237194046171396995178698476395546568556709118294546890667837257125305805491290435972112048409259574632429935451392186819478473106728857896016300933253609603401829309347727461793922430099412886284420765696448361488988005943913628635704078989717579712368108002662117687388541834420933159058379430220765506474030497618022134284438142130954570830433927495778215155929595646516035248162271961297045617398607573726483589745920533699372426100406164262950803928928392282403134614447555362181129074478848926910803164656537067649980449974655080584166420538231235876;
B[336]<=2560'd288860193491661523228792500288233408531859295598040101771935743480078500731298220010234134712626200507078291221330804695817930480722579336286960533229644454512855191480032166828956304796839829419011604325408541914203170265521258291323367681810620223558691029023745730650373487350414559021943493059827476161571920309448700915870550510853540648872187235140618514367124057832583857129939130966549710306875792895546578098514032882134844945170926315191497801394766141186308273344192830589191756863684379147096343700448855446940972154735286273019687022981395739763280257545197666118543730133475113027498376553772834001774407774390488252606407208755573763284495473576838891846092036804843341999319217363672838853839634009751968582252496915010221559411562965858346160659439625824;
B[337]<=2560'd317634035580204607383632505276021373275503309057204659250797128361278518186462414132590675455649182145726199538026822892249212744534931761680608654339046049709261824511863654422703208161488961350544137247339564207730506356811197106741052064552707392541901493556156544839607043972844148061559936533616144258588594861087647837197029912031324334845401049699076989156100002660409044391606535327652779092729960885322784818559918182458283302065323163056002839884945840247607927657021850939085176825119805408357291141838925130746239408040905403327271388764024865137065085235236212840057925089060471664481192506875967007429269490726526143339085430432069527654121592579284516429307829101373666151643720501609302020355936989071701743446795812998879497347520923530605462974994284672;
B[338]<=2560'd288866805134896447062259978217194850437037170880399510225429190514792428114854935947356246721093008799799833095612591381874646592090798252193144500047157790935849499689422859223152270068269136090562870353368970587090771624026693510063785457073460011217352943045801603372826628291657414760765382079400076758860469470652764109859435552151614011045053810321657131542851142232190368253035793461926294171265774882545331945089807825921469401830089926833329371760532223595152214326888080483491193253868312523045677770804151871118755637823122800232671893994352026781734686413743317216105761155462913912120817932499145653985095115339290249652213791074456693196467020524650507809200798015727578871152159593459540303030051152003779091621728413995035505677665749065392127110040743976;
B[339]<=2560'd317640648830935543586196610443773827370044712068348897522578383429216518829957987281322762483651304511733308987153121919749484895319256993278167665771530552181301343280042580046288563755402596797176816768799570270469452193965128572232202209952652828661090371912911607659836118660744433279339756614095290232638637567085859003819893832984191232215692903248042072052653338817204328729604098111556747644054345669174461173021662173597214162158240768931641768971144168274623721211516004896254896867957993778410238490434302077701394630117543114718989420406937581173219896187792278088993100420314557997346689589061501590445920884381188512226837460708566923986684317522339550629038733458999149361207255420539481510363958149893092992781863524568165690012014414950561594765405848152;
B[340]<=2560'd261785104747941177727001333646884974969923880932807337941654690738262645471122767058599901613201724551190872382731961116902463832984852375982106262227414666840055875434983360387251336292944897479049304489045470833300213005277947949453528311336753698562934894996699562699258250639920129634183944070514468762419798544094929999253542008794207299873767287589777813414204289273064806216804422802731921925988895999670808968542248532107505306515395644331537513441781560005887371787779027313230206891067660423569515507384079596458668117570660102039656060157505327811800428786023158258423510317457997100283464679784655344210225097714136223690074377391617273225056529829180751502254629726757328409041394207307954608620734603451126964468795642380802183568411998489660672396795148292;
B[341]<=2560'd344715300444194144340699792701463869963154267545303241411011084673362581617198450098066682680972075793618550630987563915526478280530192325497881754868641494767650551626551087078302041039351657002486549200492006833407022872748225258345802851551215710135117007908927662639135331804571893480910812126999951191867815831769544603064361628669492352649023888222967747146145973905504301197837531104203808864306589231284988242356423665024772314709790226984752621377503021150281206875751200116101057493079912148788783243250159102123073503224672449023738589989588620984708388971970382570773620535380903526272462927185652394704420503788657600318105422148494177162552177905193574287826191262304210873771102040093558471070094652150364434172512605082055002713804393023422338491920045859;
B[342]<=2560'd262010311908211026393804604341950848078332782968288416747299161141317293073905725124888787232878492153259138163461128341225893138176843058426540945104599255505873370259980078377080291197970329318109525361555664732497390166549828126107227722044731058419857290795050876469691095495711057594358888528108469834746828114408450341223123719066686913503386687861252812652670022287008328622293277111745669251196799955891891153202041721808946547400857020497931504481491871018768693131022778464804273203710243012899528561863324911564203340333895844629637686242249476534074555953827293313040729161449482358413315555720962063455266271914616959285213692528002727457967221554055989543296349047015092088423394535848403647164754032814752003153867242337235146208595179177345138686012004912;
B[343]<=2560'd29037009017182740703509297361366423011974600620441062791458802183455453104411743774036747849093284890588194310662106983594389900256866341018657900354111067030663935050575985476005216050372265787185083999252814416578862309231665642044643813379656902865863345710903082328682421360084544128029840873177738272779183934878894816959033485161805186180365711002322858934557078780039125068289514674063176860361521039750503710328895601250846505144705566906345172785743915392707131959395847708680000943012523331264357533508318691329264158322321320573512282072962067407935169683679964295859008498284760631975480434529342293632163672242051141590044644103474237721739701614703099509910031059574867458027128228554393498007690607599577960195554132684591810151980108211451422273360131939;
B[344]<=2560'd27088437478056201010721536992932335213657572890714425110168654032825378907264473943406682712105372744828226782796188145634359152910325854397702900976563563876605755766162027110574900914363577861488486758589580574810127729574545699347261096629629309234162763080627327042842205779163877013163329745475566875449854958354979151462175923437129349535233523050403989720178344469025987149533657418025651228029397209839606352146280952384315059582896785907113965418532120831870140374810025682129851334655679220972108786087459938490515887645160680306364354192578621293370280114717570101433854989442180215058949395357351612781660173654354661803381696084741547932453115219279958990615915305442066419717199005645964733722764662186049431667080014519335765934183735536326798523640463426;
B[345]<=2560'd1798813627411595857540039797543963750891463348939783533457219736036182630540355015840595650331306945483720911439864962863106640480321244616639435086515846700590839536541859954846389050764629859152296556623525398944595476243802367914413500545874307582238038052161386702418800330608937872282414321122834551662590074276730599921610822501271194715693026031500483211195732095660184155245551320957868852598062931061535703897051355614279663082400547890611754656720082471104665319446724428853422743429398082374350279872113807113040690763355234238172348667070454659205061594997884706418831346780319104826183394243942106821267372404044709747291745970115767219530588435340158656374821751739390147268792777572975492715688673000263525876962592457809583842324513840487179923092426757;
B[346]<=2560'd27081322523427676400002663267795189050822784415616359460662730894948581425511486235990469867444091979972767774034683308101990508387897131353524198244900696324054908194347487406569479698551860104715752205181960874031007449018161021759247926613800014089903839682468791107891802640625382391724727367149837708680601259022490647447495421737819858945964038715981603139223396796146392007421679819872414882933934818143463441215721339941530440623986188981733802901573108941330642699445186182247152428375342544412620788320225380779795129900807971585306860996877595852930948106430215238012824129165052983794450280706416023289522935166544799848014629374713727814346520357839562687488338494424744288779127468833960944321670887600819837335915588927982891828016455010531552229019747696;
B[347]<=2560'd112432989393351520276984298050539606857820153986027338401474401490387473680250754027015207966420261568216670099183547550011897066373421700333611268936288209825414799987545386524372232904281930485778654873969504237543806584032398889378165292902427063927662134196460413048847923533187753399668277811787526634118988145192361496726259073425116004071607174492480362663889574767003831863817434786892590903906286270931523809743662672465312894230316804473899991997850009470535020231875348438353333006682910639504103917265290684065039454853522486268301966046959040855483372347134312413435184655081327924260166341264123411694858792899032986040559027164343657876442003474055786631696232256429117629670258201342151880054135160870522259200943020667656618690495228974977455290845760;
B[348]<=2560'd422670592882260642076838129933010681320207337220622153050654309385940456044017979282218045469475024078931608680478753016444271354050306823822254809443448722591010014918721930263380470756803919686096189712779248674913592938658357959970200135407606010454384659557038197847064094915222766036363818680227281850189933261804458847529885874058819739274452069496178285588017982515919729993274435334096766217267149106295497863540565223689088890936501667320962520421961326503336673831378691613237024103221385318522414611111950803375720304011885812018874368781463882293819811622502915582398850358201041172460866519883947489607347917504983689375812453354594446953003512542832958478801435274257713792480375938354664911962722441163971214787371086705279926016373058508117861466421;
B[349]<=2560'd1693032292495350832233695645547157125036511595982662141616850039170127957571877366586842718353752883724914786459458356797773179156721991369789070834053782145800887973365139181634235949228409055656712847538151349065529547248492871734182721043909326463832486757775356020466884637379560169163426747362382124534411039744053907208186221884255776987638185066454460216364176416694804293231953772128661793640298221284269097611961055662945359124593806854948077034182601906253997128850072372248234005553333635449250424674320317751453158796576103091743445218183027188153010455250486312664166780685280071707766804553309062243286380983923818750591101903136184597125445878236299465073129099661988430242565225820664029283827592552681516212559275391259491427463191344858758464959176710;
B[350]<=2560'd3171203279955923418714505557678250280104221256252711347872709313901617127792131723679072039620664942536233874947983486645921330704839116216901702148264369794568099001711484794225974222933705518833390138470176896476643902383617210439666113979922069044807913371460964443122453608576696146074282777200617469295758758533461808718022446005126127115528204590430601394181718463131723255149790268642860590057204707564548866022067943940635593385152506135716378673298687589904801361689437499798850673394830812419946714932513012288894200340985313638506355150446688490795810372952953869245188657478806413948979953082757277874330268011561060251822282829600056617090790747592481093132598019109432401166728666952160903518077502916015061698993899363224982362130597104399969072222724;
B[351]<=2560'd12773995960922336413698189767639283010365339662022546979462191390926870083701462263754303266016630061615045193180019509962751254360081593285415300495100926087602710753113694473853814262018107574514168882005852640590513899083081644360262044080963223924208488245279315477840794682104604758289254854001755346611415528058467719833190283321571444022361367793021221488676340201143872800026292269483411609845949958185309232745010881984726436652859662934436165456446218358834759593363777501272179907709405353456276335327775691382280470599774955761848078104439515225783218518237517151510580951382573249629983349642466140062083453912892294425619884049977399837269273392301467630870622314552450296650318197077016879724235660219096386324134196040492529781874248097520841120645190;
B[352]<=2560'd4020457981730102801956177112418806336012340394412192933511336889402879446521610640533832448412683166151689821654099731161729649686428187730115517884952415503790638285524171210313611114419326239819597849075979471538008889796452313780836641025527019204048127871541090368739562482876907887613861476957290809575375058315886444122488670201622460227721003778288106140301233191434445100336516149733459637478748786738930664144724720720666975201480828317813958643169132511015066069054026475681658852478649178122599156363201885375626696305418288759585627270059408518155310544593019127146764440869858579544236537662896658644045434490354498847668822276669602099548605499173695572105231643258898264256309167464641708025955265549383158036144389153310789510551104505610524023595827;
B[353]<=2560'd4433584377995874312324054983020067281194460802350845586497927891694663756055454985838459886323984529542359178928101557758817759532272678324778375331830256147108693809520075286110466657069569709220164613814037543507662016125037334903322341854772574058772629894394047423001328937158686551691473896784855994321092338813610872346743908275968716812045463248139421686208443804095859304412620093329008160775405103381341875578649076324134665506490748984931294139350338444140752499520403837238417313225161911861717621850062523831689485072114787517528784322379271099590080540379210970029234719852128198877846416611046233712649143683788964173619416035702327706062127902624191648898884798045440978014967383875881410313675634897007337116682974968283374995523308841651319304556800;
B[354]<=2560'd11071054291864590120385783856394281804407857551243123318953159957539993916012669229378491089168258617905922410601591202282999327379986620486810421950743230048073138617562007056859321604911465042979228858245039182069801884950271281212418665491725005079081058612001277610026473846590149951838506200873299438027334345732428544787753747795034581736895073294314327587382407095571085535593432152977079965984383861086133941353984039397720946885804017560960540322231586789378777502447609228175399651496191035177546259043322917504780885767185786771185531926101730693126437257257025977356347296159952025214514992247051468602778706549101133370232159732083582437014691692626048015336817125897790082207053337777254370549670374648904586803292690575005914433277596755892449403101205;
B[355]<=2560'd11071155177431819616665738749868841346168094944602547359664078199167782391661229543186391760905238687324277668471331266952708527176986686977699598477069187119694603426650159779705329743749244425808499721885932977086953081193707160510925179413028990578470070369186877118417822723285894024334517863909712633286499109923772485881646272786215129659929788615080221924659504433986137353183181914784503971176310004107242517969571356700115459871575758822173274889643779814149854436770978902281513267707507370300206360127535300580489412555992240319423692352578612514051589433427831194631155052913572154573656833564117849701359388594033851540464685415568344970673572050571030940988213101063248595196496512983390974596390223301465873658467838004100184727495542540306599887520820;
B[356]<=2560'd11045328472419530722711103601402340070018919999523941448117835433636110000074561052525481086455315268450011203741952650469816874709257075152167692602786114213560037891085543715655574433925880683254214794591226607905007768706736699934909433867021667383091307323376389396141080706711083905397701004356157174628316946495490825537451960051202305036307813524681087212812673057271378480301881330550487588213342209917543798477218218524479396882594469561767392715264184592417096030804112379566791314503457683542350749964339754964940843745993865062265391326965444736383328206015050959418766029591353746429974612639831945661618304786381489016603097947578785981620726777291870006617453794911802313716993936312526141074042252039008824891095404253135196054968242218094804153141008;
B[357]<=2560'd123882203144010400490393439838201321644092535469098744338895630453175621773170970191991788521382359888686382879012334447200744801738777513762612482137680110493835967447039130081818801607191970110926153314140699393491649259743730764865712994129187339494402211547506081866925723363085166809277479866862538967001209225173147315036205645441546492207183955411634889426336131586537722639306291283216154586182907042913575309357448611038130277821721128692031567913493418987267694174429906410553251183973252702239904139990355491134509107644524298132767565187321427041997617123528002246739671353018632865697292903388923101873254187453951813129410517037296373972377837533641138865931739692407138205175242376327602976136790706977372378108441300412192841914987745631797366783750912;
B[358]<=2560'd1816461149530437117425149070977861590030730833980996585509258444762524297583600639042449601316448533430350327324683268349570667152611238374630844197722742817127391020268420417131181593943435767911348417399764004500990118064863652207624756175523539393670366953080405385867943484833438089396890160040235756259108807283446596162077469808441364572307084034453894295778109565244976246097740376654094999654339767358980347894310453523779219185091468908066792457153747843858904838871344413541927964948999755780997932086508172811802767901514438160088478939893159613836359300486167658824295471292424163865741133967356021412081267171524447219629246015096262214401952962216000872361588783293917460902955424547232638202360000593983493394049509542933202856509443545833830437539086339;
B[359]<=2560'd18096018994755728754842244975679952869652557254462855193746350400788123074095218946256357261679239666239662244301092122585881018068648348662919541950674252845427889275435507750234548109145267954417960378313003648104684841790423406105985492307211406951887055036692322258566543046734356911362412427298986617861571578591628567598954085413151906383161769059824152301511594503216066037641798697312925802927992304642284408256667198233935674774157210822639868519261466562714860768664606748675713456423305726950769307265140925640526893326696585004866973806614490473898778216984044605401608945943906898160497788985883003900262316713724289765358939628903380815300224902655726564485523598448150186046229715632986175940035189976033020754832012211481737956763819513326406482329873;
B[360]<=2560'd1809412072784440068320620277432767142439581028751092946201239860120350799358355838450649964466134308494852021332426248697956393677319496576852872212080907179070028848197181890574871566017684291930637565870029420110525768813206360618107716430743394801986291369884518556116514748478024039382499329611575671276514025641250993531028470103436754631272996269267257242532346704760442666563370939721035910152483599916894703378689385474372357018275673308806580444358307446926516989759644900450864562764636200516510945476179768825646728870004046771782291211944862436280516500857694649631916802421241762528741561442196633676337165474511238319005548106208026657084377070287937266950502529635454143196568820976108972884068254035883014558135925315173882458712412348880013329300459793;
B[361]<=2560'd1817287597422576927782569829179471050927950145642858448252387142657262748298202798379083471321887702916372467174235142072529279702574482524016102577264393622842295215878818272154867213005765693821464936756333333721931404422406627329148556900877307668493475057799088060237748923570919369304629885110794805433673621297327098276675412992088460270684867556952393344848420429843445827319013107988045473028973298111436181568606394489530970217214004280197653182387680157461435086693778414341365735949651567649521123680630290229356505276649193794397977650989103321872068042318871450221640507764869108045716576179183252948448014529911256266423743529587204690327239992464127437703523128910959246247608539651015266417626939051407691913646244058621043515407517294001575083626209282;
B[362]<=2560'd27106330757801270861088830763127790607653100441577286721026171886590549507980852630005529280886856821934666456772351884877132182822954409001465425467993280335333102627459438755682241815483264622612463923504326947690527257924013894884493928988487746368157401742669781948808299449758566099590242263600536139968773456212530940932983284732288137737385779693554046968721433677542948953071391383384663754817135085109232246755168221096135400008069272075754713651677500459518691459716348735300502600797734922767988073206711063029985809119095835704262140807383795121282683931420204263534396663123663372242829711175086145993836765775986982296607121135539254999090320093555729687965569415245771634400035331288057190988352002554463838180209588249197455390699044426302393122700660737;
B[363]<=2560'd130881051225700908712188262866135890810792362013229825911195701757236774809292184756008242329989573825503565485293848138387915407913699934215115417632152912055611692935283905076060201906590080348269050040927212881534828724409289337630486688956913720793194646508204423116633229608560144450723413496323416381687551412164137666331745825938545106101190690592361912340389814382902528356496951233812491375772502576734372427469561111170008926380768107398473605020928271611583425425871888951749614270907041752325457851814222512202706554714136401317135411320702945844664876969528717729434928499771008869215809317756825903962945230475075247532120336640803546939873150161204110004409274468327039335896852065882228839001526984630121287015127830824416384775999525524233699240972288;
B[364]<=2560'd28792272545320026746382198515766502915433039936344902507211613091652400455657531789513366693535354506032524205323283159574869206262930096040507018647763164769534235179330848260815472968390303567923953429394190281413214498139698141094894308452049429039975195961062506565117505003592788670431696577314409296709684148045320542864800945894854003561338957206561587307937341669772770005548832713598188564846007388542392970414486812241314256038583108171227061714463534008871197062998557379376653033366125015678146726405942511872540084000026375251994397055402731907272629712039950875194617242244775308072325482932216221472440263619181660878796071279216358540910140290633333460559073005454996021419865824354756790982949060646375555939153464748403296918479085036584969577995182336;
B[365]<=2560'd129647645122353628001074517791869509475019654956688160375070478223654553008002954435445261871782571457969240656712631001314712384218292770473461913538802615100485767042987093381711740519590076167156912247740640885402001889866315298716687190733738478557284091817010643851176786706912841723496658218649578234268345710403441078771406382767172042677289574371056157302973419294463598573135915414043168573181887447309459884634793417731521496941032185455751005281464873679485446989661304155574339768326297914889633595313723429091918138471315110113950557486031288838552920676601791352295337121889673855524910987548854114702940327294529800829077695979753375727406321343934349762242767922077248737016963997748039877709438319429651388445517686917263077433406888943276580798468369;
B[366]<=2560'd1718931977810135088461774374876941676209916755673252929050365147937477156379687190403965149653879144234604808171606747998793380201939131400334354686624524918133083019714049647389508838193077412228076878843544823967016105351387563335276573253486360903696406267549948546379425197314998103710094694652002156370538594730770111385383797269756570299735697872883727832585291437748562608377810054578713456896883444581766767754900896275656876453596326527892578257153199222677106780835391791377538782312432250500816173324748667231404356522930084624405993346580985063566233173968840578478989718733154500753451076208375307233117893657740879934351891628424273546207913025729460436116682783133665483270048076492345053820126528155750593767914157528676151495584827252649666586181894177;
B[367]<=2560'd142177733409606286757219600723675117326535341923480581148682329943790189959872763837317603212496110872620495650337443366806603094768356767284241331515781416877623388174869151653705734443434993331449790567741273110435560290770711608066926335875984246119932532444921618339545546021460517113840462520070266781034182811245664174317712967067213444710542645499242679098245787380114761701690473920528639049472887507133207444815528965396986227110643457272285291916518259013660063837396690872663958865373539014284503827181930890568721964580769626190007613353630283988300101512492012324696848747804930712502195967791490301426086975894171607336433929083385567790766513916380339744936933221762012205655713507587526267692259223098763135371906630152820509989708679311901204201603073;
B[368]<=2560'd22798329097307687844484148277083475097279638052977494428445782389816007969530437702872797396954533102930893867313991092572065930080319388632814580451811861707791741537260331568033461954842944303149745345459808761534052728247742306030664214272774353786571865521296027287647528043944141101232012760368743820530226112005698370620797753389850865961346324327773086819061704798433721824646671559303422877408843059464811392712362858283817591304687828817231813994763719270342241957955496217206145291832763486099598975278022685493187505130163752702750351280605946585967022796084682345964590144288935361271491080094518576247147897274706087855504229505734354828762290278329667838813023499793965699051895655076635441810764903962950684635087934033240065;
B[369]<=2560'd5890709092508123048289110339222766559550543700560683939941330397185633572074130577215319223490990070284501679229699358483378652582826826139183040611788762265947144416390960763241273522834419812211339211993960867547564008108313397411649540529014512029109332532896242810563572767140973300192708927487556324625172067605818685062195575431232612374139335768552863172442441555282981438752642002762630682804102522542387361305253466916864836278051339851575935971817529364023285970628559035253860483641331471095316525998905488745996767240929284721257977081531279039067160819750315387013098889401410883383664904242548726570585256573497737969148585350721419791431326357364984531330187429854930452037431334077953389611400960688384508389024231076352;
B[370]<=2560'd349164516133983252332716805237657968280226581174685237491423208106564036308121799225175458650704874688110095419230177221915826305604644221372583374561721239881477704182445124633958742493235892471474695537525280026510850525753713311169790166670097141490876362053313930949160205347584118201938957762857889424016118636440749072679866800182880087388567715518791714680168418303602245680743724302606994478722262833736293136168710571889499584225032070784912205648526341067986662502716298522945530554126053743256110481549555477458989481604967586078811716166651876421857835870677154245514801417754533736505736620696753731769745440100422246278537556024334589759691409872143236314288089884769562484292450501324417535053053704703162708067954458624;
B[371]<=2560'd21363351290246281412849408225998775653228730359772848071930886796248188470873268932259902118683218844093723896269369050804291032338011177030197820782139993534594100621147679541445957241416991326384742383056041081852460129032070893250071684612235804249164974169579496938770154013360549727521236025754961800948958166602723302308685136438084561475634896367246132930658178128374671695382295297870567668310506762499900944578520108588946672800239589505258516632467767151486707775165771039914189883174228542928329568026629123791204797581470915777235198188185806046890735725020961747351479320843063008331186570384030811894360952376311331837023083777059142929267798132941228298519025177954011503534164550939342009653034684390759672960772863005040896;
B[372]<=2560'd5217104701221436823653762554649857160319371686969910157514097568112800247566979068484759022756197576361087429572312945322949539945801113141205348185989587935386924286176884850346377002948900212381850799103812881394500926076241940345752047037820378103361771419885941470916081207849027373094989976386305192261591815108723664020223575490620224083673185159115528551178347914819985710179792674059663279802922867679326074985861825788083516767271074503273149268041557690694265754098890222320058713275922151942158218702832585085786114974152799004394862196671935858594149084613104563556336469886191799041034509648387489760136452945459145195468759833120250970812702164555014752515273645830255990238295140975605498536624983833826529718691298287888;
B[373]<=2560'd5215666867478140185748632202797783309832312819341049771384778003391157008402020471307210826908266569327152989297666907505128321444063319992147303147262132768520806632800160005046890120993815654560903847966703050139478413688510873492389181069880917374799502035543168033294133019905712869733413026637195228250118804488613213520360285761120822879363984935979672638620050448210062888036857267682082311441998639245453523753649691483895499918644173885653616210021305834380948728985367263337302701778630237984979308796351952036623333235021943088960899685208546040716319908097441948759268519234286540792828646569049501985063695625413712753256952997853944013270224965099303543215512479912736673174926692641043357601289352094346114798873240207392;
B[374]<=2560'd81019570741491303426776730564147229239827060298609623781569942111566716534692170237068491836737989071501856680248912464539529105710923095637532933918524513523942683838763092898951291149824714061689506443177555734678999713860357107190806998556252518989169114194456717756508031518961122087469023554923738099495024399898270133233486639957909760870738718482829633238782592773092694702045350882985422548315906093456311567119658756240775745318596940393428107999374292669596374691719812870040553925718064356038005776664492094913647971116167882038812864994624174121060639272974563296989666462318673888114211135861359926548491413985529711794561805882644061294219518095265402412713033560009003293610036629710901341796702801268505063936;
B[375]<=2560'd5062487855714884506332720991185886570275076312780100261989150323358687338959518523069839940508969801177344478671375307291004508291999242737393205900325880039718736168158091425860454475973663651667314441465002525840957127860465112993079239851177346575438994494576969514509038558897968121492377765234455108769579535752810832125686844452898816238901807571082851950383568086340263688565171768193153246509216415439740865626473670747730340029316476375008440120888464953967340775598111656729349224560478061782806694635195726050562347223577052201873607602366417092889392398674593474781006641773353284753829240048973042475367595008276353792021404233570213646083218473503978417263138904654554823820285414643569198783120291716466234372;
B[376]<=2560'd316323439522980975204659822798492738906757922897432819670573669438458307480953532351468872289040481281295670085224185172708045100771491626666415705397327662138823034664791911723806430289248270895622390702355194114137996982920219126127874235016177874008652136518581382011907990510302839021949159053538836622277307693957185272526364154441186904722311862154454435601846205747852097482687498832689495367896867998764918242022816615512866353660342774599495394575984751164328059662272128201174695656133884359415646242250183159056792098922582311239289997193202882121669478480515793549646975752929064198568632868246369864070349784387213116816165067411461601225111755095507897938427363247073627505794286535117458003750448893440045586;
B[377]<=2560'd19765353071606805099374916873917320986471171578899062206951978624465963991582408994249437997104740028139847010909010185790161777443706181079942071352545442457139003190444616289368512614333565636437900300115936592108412537562122569732722647207336088151776296173998653436004248895347903211589275143087164919214654501454489280389320023895258147131620618513516608899995056528680558340579821501096308566984622639384320674101541714785542698083330693282133744265952960026490587330547636475272992808984722255673299417170199880620280539054928848492040531202445657763997679809941766997980722543165673118401773306407571296675843700740093640731995442146692577307249685550569393900678535200439871150471995655645822396150105912875430145;
B[378]<=2560'd105844015879078622111376856045945063345451107374587511611438975902983563222263827957806097164695604750945663384248480056877132044974957035036089732708637540012113608920109938384109077757173961495711503300296938952067037633319735239635166781710657932451937711437653283088681603176188103625691546421871011459646723462728477298399667038595166842490737079160652034882062930989132140240516218250850422269932158895565688851506164088105813336512862033668581118131460035981383146536550116410054427758365487720140553284123703279170720921462180698231693889231657690992514729671460136891998579534988981364988899096169347279999375162832471137886490887003596072088993003249595234867540143335053396423614080111273572599201796096;
B[379]<=2560'd17754795570684222452498024990272947324141124153796922576859474535435122392255915035528967307060306472071892230065778170370578339052677350288760718683880222150213095150136748653939201146138714876337963361103885992749967534299144299127706827716129375691823350764664123861124836561379060997354333807108509787202967218192940498099847897890792432168294301790994886154529442324522796035911715104717433955687729894457650513383161120397049353292858520413379226979994687564258426368981171430110786988621296173210169557818738301991957249016816123437397029844419160882735416472303857451929007169877911014150024207192789016868914438583102394548767373638804665579766167024175345367512123831848368519131429334187035865463712120848;
B[380]<=2560'd73955390214271253734061289446511865964532218298750074907774039146365771723684205471169834114236433902603978870207386296176398789732847964688657295778066290045333910310919408022195088436384052915033127055076891773068703393858020111612119473669806984034840190110474978332949068531665778860578702666298498993530273366699846323603774655737742285295365182370028020994849189038599351177291399077997561376299361201236144775507863128956428258925604384429409216795173086227551129817336661630282774347755717489918619171636174641235392506363961987747874129089393658947062950201142307061576835529556335477372541058542294130453634684814719278720109762680073365788655094591172072798238662779136011479894937889925198442369384464;
B[381]<=2560'd4601989183336459639191606828456500973356309606278919314330968720502572470283661452377726396844708938076955960271268551595577904430293676959563964988433933847538755513684083481253287759841973675919247546886908291088830501694375357918525428342224861152599290329782869004163787235193518124173694343989756444263251268057764892780478528053435486307640692056428822412093502866881417980560349244988777415304768697544545138625701316748086759969737637102824565924015841588250084526488870903925421196910632512285343955476876605821227458717002601683448497872956796178980669813632216948332867213433044953768133779806436190621010147101930449268140333867074500838080816605427203686373718573945138730833038147380263420246888464;
B[382]<=2560'd4684518926687037760893605525714161606683514176923445398933393274826038122851970510340010013581430937508507883468637915810023115369454851433828237597564250463466379976497800482464043042101734342243408502280323693005027784550068872450505211173567831303932690748538772327049607500640746491250124989378453437467379353756993055402908437960581061007961660583561715802500332615157292424699887373684686521621849947452165868329356438223988657562764083837976643089456828895086701529834889727109772837465542711817379027428703658842975450929083158846477636457847132574132388871482071185487083711768948566737844577498663003311618399052872187745893831413229422510366221277170314503463617189925889446413072307936809717776;
B[383]<=2560'd292586242493234440242830380876841030547809808077622697708637582556583072146590597945611532975283400041108177429977095126998728999565389767404042222847052110325365093255369869424844908579044523908771049274598342170516630019463250154385236794077129319016186636579236403077501053562750728290788662801885182983276635457064177472493466595551806442508717904932644805534807664046120468955645571847483656259670831794021479331091458783620489641075587089608943779943941282292140709632401403901894564855282871652504525057855946643323060563995788066031355667211351990280826648947272296765918199717974790816144982887231288052317190110836042611341085323205567525230134016728675091035973409400642384571130250832620032001;
B[384]<=2560'd1143175509063028536869080292967834050283664652080862936223730434803826870833508300456941962073486356555052187026995835528855068994726773698149484890526544628749329107581280909538812232068295153167302017846357354119991036310133824199533202090512275956968828850950607203691050885643042447443847188034940608478033813389499253955876285906590930146434727003340326780953074286134030103669334709208581041756372667414808216068539604710444406878449446844682719480284391543703652802430465471472999849202650173495870807140645353806162852457796878574622933392376022827193139714718836920978704410092713894191001470332164155665379722349290058817757911308945965566488114425806035586853328273647384306622820950000795648;
B[385]<=2560'd8667230658298935556192638798708448511943263604210819187330477369260760532348937766206224186006640140833876014214901481308900053080695753099917391030966742153367711783099800033981237996389563382104195877250917567467034207210220603071638548233607475369219066015322323483736066267888684264074447948358179881887803668103520834816897964702335289736978577726715373446824546110193951620752914967819071565034828154314028049411504019353753937261516921154432671244853815142299706310384719949720861767856676080377467862577390964766669756256673540422558920912664377002406957460959944728823442651750068781313697271801798986542575631754657395621132224878361223859961098963289887523437483804123547859274499352428544;
B[386]<=2560'd4464571615034770476949257265312503491626110656165841124871128744989709921326976613944669759980438889955375512929167879760733078687151994775266462133915639472887241148185029577537893034259182827585771240816447644050868515353562669390635613467865995462146119295362185950530358838441668678495112685565556559156648941854686107707103236752837299723159559270161876400044860791229626939586025620234590337036160500019733957332673133827413788819481551538266818011289347636037922616388498142196661208877848614727745647461210167190817377725896434254557091796381227905217130143712984902908209498854749112779260736988597902832553247914939192585040651814410047785127734151327491579952151045438647277202046481072128;
B[387]<=2560'd66983139811775772252020953777725520700786021588172022601229788635689862813858951699853563349959919415142057076415408292622955784799109081780928379478146321092764617848102720058793161587632852003088093746520319627825557200206277498506807787998121807983592713443224115154898972645118004556285431157113536434890661677515607129989126037764271073945830732631328776339619506540202902732091801433153693539127277499990034781677629190206968109722938280433272285695567271405017138222753553304078940397845264860399961284455204275216983700437136651542706791498356457207743695300132473473421777341282999214786474124439210647075393166648348480176277178512425303912464605229042146682990134939089545069314964346372096;
B[388]<=2560'd4185480290431868619852565438141202338852557845807287640694888630284142372944430861367900714620895216892601280275388693804303117237402597612036234956499401772787300360761047523810053131627143204101642443841226830411195139790239185205081153954077286860673279708974282312849235655842827205596259717669834237103261026074754654324112439000018138823862573442064867338901315298803757294889455311470981337925005525027069677608468120248129447168512414858873003951144366137070183607314300355501049452950825198791171365095779982194587335005835909737754372538173059444500146993679456444252631197926511366662322401526337652810978780661095765061526356742603320601124583222537065530881622591592488995867235650109440;
B[389]<=2560'd400785353137346596115460704607271546206609682149521948596158173019652256594043233178578984993081364812410356808261979344404873644309089338860218009089417078845798060469010737568774471240242478796077073288516564240049832913009059454510407082864233949107379027995444929807408344244016296052724002596580858389098504250882295234296492856111455818640147273935613434336485551354951710547472331644252805602121543030963669849198835884727818984829629794465582855181119467976764364315387709393352131550221101972850947339531273529202617175236322225951738117212092587224838803994305669124858219873057481951111354463824107815445695361439577559930809237932350794780348404871641023901286469442859949427098991287128562789113491209134709248113367285222228642205108535296;
B[390]<=2560'd12828159211716870479923636824733980678479828995339404417731211781191424518744625796297475967213981712660103585548098936051371552519418034317541039390210278932988063982807511421324657392458809495237932069409154566273430880055935654610401189129115146262906545732866109704089452842660069107372396435804980850078290234087639544956494707655354018432603461661257705437992101452233488268251011824274528979226917287670775198083683171634516540230235022517636298776266748182977213490086554381123213524519194485909094234901710782827722609993447387660525078642831304836460014443614916772159841685155937164476143994403227102554068368447431031767987336596688000596423996506131012504749483885448741613418240029823392497636891981450622720471652904717066125274245291311104;
B[391]<=2560'd12804767449820017847632614557476467791618325434020036711819688484759767437986396786403927946668525922011724960598120010456467940010854220231722321324046634909250798932551937394450685325065668372220725430429611570502556962551173181610488891557163838989532133795882500723534204305720609247282753843930623425359705756211212649523724534301359610913423026437270108374098609467214368393484407352615951268920989067290798249023322334025050094817464505441027451481809386637164943989438640485477623301241926181470652929495566273286145479644741523150740443172562704861243497734694416008041044746774907144858967493029403326996555072138093078564028283252727800626869038724927821090780994555670249788407684590886403416012372963458598381459801101304581174613130474422272;
B[392]<=2560'd109016741454249125990573393814407413037758882684390258038289791454389619750857931050241916266475541557084291851859773360179737269859573391039682769652008640485928735845457460282913905602382112759419822298464255920896662242799450448791815488694588066149924710758290645006272419387578632301412597165638430030285322376022678144829510026640867929129195589031882200608426779247359770913026609881609493308872644045502351841177555540344990262795248360273378972471690094884654798458088849442713662181970020511061626885544835371101867371866298960153178219182170601311975579263444995882894947663009149794365009250680908905974041595830303938292468465524416187158561966675513459984132909629807854367727964714789519968173528200296667421861065165389074096834862664122368;
B[393]<=2560'd103026982330438231806869805262035003116429331390727072872701442756889378589839635819046393120234651255542518143985760046272043000704083457876640687446634768835373616546717461225824654295930382183514279190496072639324225533399125760821184765599001910632307307932791279084597949328049030108626430196851708595394434937175131862352277689637560649357991554866181625459045605166739685531631956562860967817498572497230724903445199681020808458544652359692544133164351256040696410712693109624351791380766301055012589946759763502212612609474160518523276815181766985793532466457983879990657590471222154671529404658449727707843901881884058177670763319208137707076887402816522614357893967088188742754567987167843950979970310397749345775055405581632787819619825932566528;
B[394]<=2560'd6437614734768629700104587567754299210943668019526696299063176055410439651889489047873120005539771651531508369871141645599659224934227839442441154423622968476742734891638264551956397627658047737604210919229572085839356288143291127801185592766583496481589766008751628592875940567242952136767816752502440887880463760509065400968334199021959911397751860235178521288721123901775859926308798321002616226637112983963096459618511926631064660881325364430799581352669768061851335865647459533257514294364285781452846980764582498474083820495432322271594243305230647298332278420629820360694105685283002079697777759968558957622687537251676874429331512891168036709429620109053447377102909251285619741370947156924985082976675320050682191918509386231425845360295334117376;
B[395]<=2560'd23489251465925075230210151185774156554233534484953667316032739986389538193089559149557302552408464722169434480372331282021158185487400436747296586100101689568121091109491216164216046348025254807780332018189755195551081845884846116801386263995284721936099365983312015155384769343691200307020775126092794482177169621527480637485807626099030631073982746959445031837302271108348226641193498410557343758420820839223344249747409683751704502216755923856507628507367907613982379465498618958998325499586378881972340891224682712355961634381718494744644859862290339645747506308275728813211117816575198465692821668189904239464455547260107978430638060352503505315717013220729232741179160383188654656677066546700295667172905194964872885410638778314684851072679280640;
B[396]<=2560'd226950964506300163895327879686879413190268394939194869290553088321072998024929926822283356119754441469267322452740612190720632134237430549970636273531643066667380809714903418634582426262221903966236339768006128768171758922939281836363588542549517792350840357740283219280861541991083171292370311493280956898732405025369993455657848264336907953114661394045363237640186161976053607412361749420903390452588749212685760782457184966907620956799835947674635786579054619985963633572536760350500779964307799625416525450663981610445893442859891567776818212201374657821981749238232348416373677038628011213563064869721112610472799298627250498941059014541602792799554206717116716269377788313600;
B[397]<=2560'd1493041787808189526630419137355951764459199019333429443015935368916255410388342450639531113568373300383417760424307677376374729827081739851909033428853748093224650108279417337941948161432077501504965771326173407160039342449617121192820468052574135487067864363277843503088622357034128883374368177612857557980844234000598752432345514273094489479368350909283754862601454597522727331993775323252315931362475536575839804588519600600044717145558339151144226569816912804471866008611511890807850613335270428343241224131229560470723801762966761574194293710090193003453150169560152801892219652128605765838968530342428826641709929241025506317734903438404818946356036832050983216272339237484529383168179371696575864793467707748749661543209462845040297508864;
B[398]<=2560'd96211974006015123228890870695476079128313546304191348489864588473169337045924697513162309585187823279534156372635601753396951302501769325485138405466641157905672344268797937701775770966987445869504049802192998170055407555536084785417222561564452955480300920592086943248369475817265582333404926398594044410758365914447427400129133912422800904695115137929704727251057607084509002452351362697943301872122893627803292689159997178362819530527080665345249748404428174577696793635198997034959773244751857882703260613181373088995220773678312365247952887676742097299595459036717791794002944036401499015784891148694071313562122408866700818360345940919850740686511888933946055346907858436973475313255039690336385246053771623560871014360311206193768500887201792393216;
B[399]<=2560'd413227281832625178624377940173273591162540363609555784489470831439111381486194876550285338970405736458241855100929749914339507991469281123866255135790414725314116992933493461327318008249176977833691632202369417749102511739199807104687284737448853043909222502590174483278526356759190423843193117454915424270670508742210943504760094337534403671474647328496831420286741485889518529691520555448820079449783785577452925064713791428694456406491778611403899960225825872726972709863869381424874106330782757421325405100439649123114653157779599091092224481382601794963512797563988745246272064415222338923837229267677198597476998978928152463648876511997627373554003411789552860535942826967226625013413075074269829980138370014007444723022904936760433744351670537725392973725696;
B[400]<=2560'd3302627480576900045277944190604976378912910739056775796140643191161137136822816672068975550738343136495291137686282827595474639540795864766607713169999696291636489922363218576064347822565616145566051491435515871058351037410995774910444469806162944074559232763676152985227776630273245227772854649504214651873979915117460815403881342331877048793181732138798885048016705052406437076679439365008816251898557559840287987029374029838950530068998124222079851935265836930656105702942152782964918357375762068822692659282783448733940341625662352147852548888965944775853233337662798168216196585408081340426970722619743594916103074868938535649809155062779862640100326092962992750592;
B[401]<=2560'd860029666044216403279718246047628749594245417734645536424901238578750269875845643737530959674976204741520790673464017687272150225838105516786882402733494310290790381432961839546986537180766809565027488932459829415359056563678469777129075410539602058170849268681149146785530256713049157749344253363564471057948548832682451682725031230755873526152988537918431275580433100936397101397302356183076958291050990862378696908281480947416808744678162377717649924765252621190534655630280640270968324188954923863070954196318832791063304127515956646918467680280215008674126180181364484177087047783769134822520378088972349659344028831538001327319196907653692026535365640087142400;
B[402]<=2560'd53960134473244257663923381946554151675476574431959456740643607384227106989175954832193960162971939150945410540726669142390153105750859694199051305599095912646592092097676592012509785312388552521554318299530906491588030809844953404048593239318209218367788463601464010901864547783898051894545343578870425706955576669698604697631420682104774695764026114434601423466176612317325801850466837444930138611840622729758310249207101035759736350752442970176890729481194649459148131789789764650517804752114319839838962965168334372854629759079433892116772945019168314062976628739080306006800857318432789212814133867374184165598146040082033553001095005440082564273220036287528960;
B[403]<=2560'd50590851170528442469924034036686409671508515735438646481693593018546606398027116718407786623964665902646582612514200169992083457384006918308989623250258589866548495416493092354212367200801155237181460392478548075097822129010185388539021426762398811703376882401932052123980874514307997820839381242222920252349365897538211324649181242969452329581180399793965249944496068246553561384233820653711990483597514375719825826081923396083195191626163166099390653586551092260871091710975168485243430305239794153067038678677162172524895438195413918232076798437791794636846495022780621969804488323643735475689450779351489315726460742447874040617903293296193912439872225527463936;
B[404]<=2560'd197668546878914856118256231353719449244528063708079927970389590305161422454533507139299562021142570032584759073704613052319872352105391271242604804990500728927436872250942926301011496169872362454520294017154772907776480576701034960026898014224320304115225273334957843502137936366316106250721558773044632320522137994770635908293100454508719896253620365964132534002283037030671419646263117525525404810331138440475103393401006700484980253199069521363180279111381436249370939599886305467775043955174616846694958195148009235956674611250963535033391270183485490813974418728554816983513351188433693156275770329263070142571123275668990606157104974148819059448174449000448;
B[405]<=2560'd196800527309160435749293526195914967554374265772324650573058265241665542873582889750711481794933230412591804575787324660603951587772009256225413651943183324312637240889057620129441773488250087530437187649232905081968452630759867560126487448369892761858977526654263024456072561594162958839979662570780546645432824221085394413732056885834157173377919008879891696671855468676519175928728864182910452141827762108609402030216211550216526092192857027717267169654061365913685864829708109646466776804142523708013033118264204481148641435796143039225423227900545852067277746100622059042360458732927433541858800647253562841157053471742650310150159698271070486346630376194048;
B[406]<=2560'd48048515274689558292910177415122923251760005619308829380968291066398851843661479026729405079452228030408532883044228869901226415825360226770973426889342776015004953567658143322581585420305119308606117269216833425183650797968412063231937950422867273824558263102563967396579208549735704630862480331486624049512360037801411534371777743201701288767014915897587730782490150733599980758667586177103249378343201636644327290806243459911054234869942507726740010973036533766006124173071901469340564244760652525762082955399762496545050269699556035979597761446927952030754531354537741328704403227420871395771142523341401172058735482746649294715762023147904959243670781952;
B[407]<=2560'd12512204569718033164482190001764712677756554887152306112512514553358956937386524414177560280328254781529791162326606409904199297026974557072571981275791762822321763705606288719233957055782477650455080803853467832177957652342829647679330121529726111158827218983002351973171042146984360782024877658161325460992343634789264550700284471626528748477217051879386510486406094927399255994771133011912152778708645699286656563985407550799232872227699617960151133620476464496137605510234208524605025795977300190159429785906873223178579081416466243766821583561555159154293203335350385729864768881579653765037920938304206240032951255156854273194218076418358856394997760;
B[408]<=2560'd48875842456855914879678186001164436263438736108671269931148860691762681969721710669953301219014043963504843315050004953866237823828074759259856734546030362361914698818197524612547112150505506938461838465496275426926065408156527119915142101710166547076667215999652779968060363692490133271062071523635558529618303160168703682417276130321837833238730366218822945633575719316715433904741634816053369359534767356755951865113281328260749862374765978251798140688786347228449734372057881406858445693901835689400552651808398500901667181522490793956659410901044663820054484010567446262596387798968425806753661658856345462974166061081619805755641767088833362395136;
B[409]<=2560'd2875751652122056253157370280308016895892202502076527998661658131443732181873918529594339791406834083416059888434147712635875902087383653994687333846877422543652497661902955532809112220435016845821110238420572703780220439929009325705216414750983706710900015207586914646711008138334965891059183308175993566084571477944888626491734947594984528486056252420521248990195843054983051751668873006401149247819367260381361739074342301473547578416783611071479819088447722761442335917907689191123237532075424066344131058715626137309131807964352535516665598457120401099918620689829779968020178768597037225612385552264367066485598601743655575957944374205629379641344;
B[410]<=2560'd11233425558539875176110524770427302100015223594209097958299156258110816118504581897163781683377931261674551931418970510301587541314586336041889335224029644060927216598018764079489635377123473886903438743821451716519739996474923537725959735189686214379475795118697322572878996199725205068441524347197615136847697580421384277796918807240012800578262188913040140002550617834596236424014591039426872912944459276017776231349647499955143990804791703567044459496172395029492242778648452998048621136068422765724280162965883158875893575644993312835262462674984466196804197169555913566227989307374825428519254115884878694819826567655337928590851348275319013376;
B[411]<=2560'd46451651406788871696489030128204993265697670177788861770099039518169007939483465303075847695734625214702597750635218758318066420448602843740834155395149161689812715396734844288847015642421363467089424106414142843624564762728961484161021100749917828122373533376802337308886833796096320582889569888655133622525863725685267528789384152245451971997045732895926066181836794104314532661286497290627851297532054796445503513601118797644630102802637458468608326781800480332268882191919805923864575324636066162561468675344208519314983128786753224538006390287347322687932838853163623147480916435565689400437251666775651828469465464742483758968249206374924288;
B[412]<=2560'd2731867143358834214578654664710124436298605868899388973234972499016861885255040292844793548744451914499448434952247173461417107440271175663936192070686193263347192054571985999776086987399586751491425554719472245276705567602514513808443315877980585099230469859886202265352747831273630421356443763856385597620020675993793492072033246130615561707299635762725145442297629737491896522398108839875731411247004878958791064002735742988969106444628316162203136653183901412407229985682315394469378961619391676605167131076903993072047183110045581383955425064229861204526017067436971790405481132003768333746193070354859716112089827893673767557590740000309248;
B[413]<=2560'd669726491216085512492842139083118432240842883003764896381641615480673947073414366031216543004122187495305346465719420789055915452857600546764196291873048643670698122868470076620425955098667199970402680163179439588416421701699267132454105457003014488186729950936152341435510372419047281536482969001132165220808248713740041467669873031676249016969151080555023680937467822389067943234483873052152747398455784595266988268027649134820907013400905611645010944545149470721959576825682588820216429060428244817654574255494323238099616971737968173946308255722186418445507817653163725689762391228791163314482771416093418444857759282748422301816165761024;
B[414]<=2560'd666796965012748854176328823707991594324221729484568795484506752720125048853068664831304057437273246307537316001948723512177259983237511493728796835384432948223268598886531958056167132301544323776876649679439341593440220330231048060060318582175216792092318455426555120983955013961476238525664118180056799754095774103802247658174989731743590073797111713489424651496813383698007129369204718765831462411008397639563984954625493576319524930339756218380100015184925860234189608896462065463136772694948291307227683048610304310479585022741523565955951827451572918743496163984383930308629686080162437279752675633227580583893123111905064684992044466176;
B[415]<=2560'd2605311529851223425871517378978753962864355180491149373094425968276612862714315293200298648922858863048285647453857871005851057571128272085322372422899244953230369387350786824277530348990462438909475726412316402021238527900483752435684638579525058874884719878205116846339398405825950003883446169852089562597052973682004392773651546120822760120318263865109850915883603566497886982880587789640521842436365717925958971159939631356001706002895770035272158196177322624539197808166919943422279872925854528379910365075898965028001302575372949415586990975794991482656363240779098929616111714216727981141709293823939901777980427028160788962476032000;
B[416]<=2560'd40084359876398503263920403629739058798637770770969660754133210542568859628435807219442772863937765334867915590768758106080573246227559272207544580414660195401720530060030823015297688969968975929218833659972581672122269177685490148414631377849354410764056518147758485580277845913680537457778868139742279674780502323883248137220039236081664216592958811167609175656241092684172430602030111111642002080470946052358520038666325958502390274705963388853872716290644146853122461705412170374015697446534167542869423944984408320659177911988324644376369847441730975057919046187747494678498965634849816791555777384495325373682687311308231184220160;
B[417]<=2560'd20699409315623259706481519202690246122145990772328995031465978655603878777784521239660230481207288135501520802250333331212556943647571162886678321460829358628575448171240004921137020148938553436124610847669609820326911581860372255159483268905386687491405464894728371594831047632212175093447874380601380422915245713141897850011730083692285179717482958745407533151139284839544530133427438800688053936001743086034570445631638999737481797531576820074892603038296143814657434244146765735537413808639528489145474208506825710039824839752663798865202276032231540824859320900863321666065306691009236569723656980386548688868288546518744432640;
B[418]<=2560'd9783704367607217155965650421168079295256024994337022434900955900297462975621699987735723326232031290514423903199134080171537176923859627549590959028128368163682282194606434296468541434880447607378259610025486136855697459809501670415493916711225558490545129113358064903154830578810168108594383007102539159624001209046683013359573641316815605628579831529631836737949019446562260499790088191837853694812603246186028488871234513606259453881352444754517494847328643397225978432205408374542936032603518933844847252104489447577711566828813665033686768342938438096105505818407806126525955632871096987541579052922727112610779702899561725952;
B[419]<=2560'd155248102161804532265799015352372003944753073282127399922613121118285941587328041082010141816604569914898148320257745456510002216022014862691825271081621371542558628617307196958778920057651109299051193602811075102290285106277434211038082090812023131971112559580820782156518766412035008997399771307797913459175829451465868618532013756886987103740346090748090558232918725877502297347386319614033860015982285208293739754657531995406478590083646382071044547190645423450408791631729063336375478191536942736419717458257215154646272710692716098833918453256314814412329954580691474467430161117068031646389871653163720883129309858877916839936;
B[420]<=2560'd149285362750795478616626233088618596115151891446191283922148936167838125378017172010543053037639133657370510290049247410295688405786182594570658753455450633015367922031772071494892081492488605663495058698267672434335678533090669864936587102615420225864863784511666470094926900077116369370497085687869582921257903351593621151642753459487690506647902755154243256732488151499321549480885443757762022363121056281430398741646908837589713189152279239763284781393922709851321660899991947859495994800682114760867401398280576111903582154232265805827436190259964453667109880955330239865971336658984305106909021133870527786397426190909440;
B[421]<=2560'd619441373819961736995062977770230570646509008597609665958377757846483370892313422117359782783531445499446504607341623852809284987131822708692549844871204279301752928217869266433474478485749903316687491003300073216188548664722230161398475954202339036436275779526481419595115200323666274917592498137252425904445542869322084819489019452345156564551241007176353020191374973390167814432034797011357431766399424694293269238720726095712815210825914511697212194344405470274850079907956021305270325932386642022487514841637646591487533954550112469144096636663975288697025127878556191583867047165651513666479456797898627063470102675456;
B[422]<=2560'd38706293626204174917915319523918868819543385905532313764439825136524365713873181338689214009830514492196503106619248213222871764701764222469081812914197872132340410115937559456155849313496343203011407125467782593582241812100212191088791451857699063857025319841848752285137259245785162421894920802188158410581975558296975639948653442027958686229274373514043832367910871283726488171634935898774877987196621407479708526605462842047623184179400868694886414752323452333082162673147291350895090492643268312324462684088891878250414085446792348647946106893756449724529954684477288273978118579256729515181744344733014978448794320896;
B[423]<=2560'd578477138529316728128364394270364147576179648657484124336509229182885963021267760282042011573884135503305267517950476023321678659033464936497185279565103083730285599167920435348006752304653869042478045162098543473662126940082306217180262823295218270126979724171484750926310774509310822212307127316004741868338705071277581774054963705365915582935614226234260147587299764526338324336199062507180527797525068286515420652825069656611897939040979269368676043546124358131156699619291798294144023866238226775782137728218927977084014103240666601467939976567986698912293506434022004057607557388925154300926979124159702825623577690112;
B[424]<=2560'd2259124905050219418599973124010168814431155237605020185632529857477020875723843613741518559465888645980231469587426657031364874100287191067086398053926451168012507731304912618292953569349728138720029440030364294863266522506834489350340245599520260525694538265674089137250866839098830988192400458629777466265388552264603572671407885070783380778070022155060929010481602801392153095443567715613558709843634080327266987457798853633597142040840365082264702728593168157243098328921637676160368722339034400393704572230209676165873405775283465194547541421448453626447577746262465264168895103539188078512803900663524819986703974401;
B[425]<=2560'd2298100263170018917009698555547045711334245033480007977141604099244277528882340229441160715826877080073437184162890913590925572232380849076690031762093579334169572403586269242180832392873207426691766964484129758625917259564997567576982543200307664002657492806571223558998240191997629079879378407315616687496456665244562330260837357542926952045638214025551382896696205190349071325414980900875794656058384807751036509893541280686940115834911680671240600813083223011974527813062348738145814862130479731691105747377258014674570853924201810685304412849339161988961700238801209001688599871200971661166422454551846664011776;
B[426]<=2560'd596116262247883622922233253103634506847506108023856972063112939644088604094397050081285724602178568123637344767639645262161224040361271286972474551165624341470620904812785892568540323691744619907411751618953705060352598024769791559231289866869060469039608086590951094007959795585553383272386891910314453406656654042890746539481664669851549991214093319725955258885556256549197794791125445178516278111284782900215014170510788857100341620079619088235739466112710009270179083673189299751152424806540143722640799620850904962813241993167050038608742820749577696300878597125425204580401337822711093271232160903469203456;
B[427]<=2560'd37121856896787398990369676030576741177812261630039655216356809475175009905790052686797351242246386096245223273086919601558792207886313248310731789625828406944128834458555110123868373803648265443128309347708563191292380329555626536812389537859647910939969030276716733565174628875319940035841892577033987117150422716277619306886244945842228931122122110892838111309752983057943048661038570775376614664682938041692888949752968244521128530152565925974273865819800121773238251337819299363954004818001400321535302964965163120000056705270637774978876587622402607732838876271592880304800238138420724069929831980752437248;
B[428]<=2560'd33004044833135452603370796523296335235966974307234532782697001159823087955912928021969362388076372057136101180267476602002403263332600785616246341001239023202686378009199558579748858411377957562894552560322331432732214353113852653169416710006598266727676742186239048144334337314752906555176984517595659457804152933101116273962775580862742724574708789730981187375396147458415076742681407975248267632753379645203562851521855540520444410955459200408376516299490284661960094260705703291619828574351743061558846135933837924559041127506024499268982002412876378666722864938870093327869516087280561768422518984120729600;
B[429]<=2560'd8061424140310454880900279918290852478258089644720012523176392927296596459535969526984469798231610876626501388243750636663092309017978953358817054163388314512031495479526267346586847016185898541303384668721379290258296901406399087409099314824378023337850964647676398941620583743076749395976036015858435535278770253658470799459865988591786783674967492363067944131571195972822248159478569518661039825940264422927401474105625312467370005008177939045511811446010437663087539245427904262110130901105823026128386749575786130328747199344158769708251703385498162449389827407858181810025835006115675952541402660864000;
B[430]<=2560'd34470947149796480785652005224947285203139703410397759192756712110399638624550160117957566465458884852444725257212270130085004333816232366614237973633625371677516166593972984613955656656660470346771424902269017164954269956475694774728099878205616650151060060425475206591950784809018225935347534470658858269531518265909154840277134026697173309411287044400282734066698021780117068407023330388874160773654466746949593373412709495030151264641622143426551191641628698524636099211582659123658040885448200552791286042125663070166782936307607629825338754503724244936241022682849011256367386100048701748478862744649811802193920;
B[431]<=2560'd551543044290772466999209368707138932527517800189565224279318798526624693754272031503137089454128477479452381310523261903948613766944074276712931988887296310453252522204466459764320006592923099602167319412514199237269277173194692037822697403135621201042440539236598018378690789424022147181068763628849287540693278432312743690270194482674915576885807270821466461440325843580047334889278217775526417550442031768028754858899468705237118847040572760867663783654964520586304500383536992946921229230514235635443814917951068702060661236508673492739234084133471770516247714690877808805329935899173041893796624792482698349248512;
B[432]<=2560'd7656438804794914812417123055421329900673201123420705266701169535676447238388288843555000082405213490121234688485318348365235935767032169425937498517331510705110974510303179889477640182740650318338114739571604364879466049676591703530842446624143420200913165492523331144498976175277927455668872568830307780722580819946824801705593267133870144820755541918661212530394862701856990178340843007756582546416545068833666823972398565005796457989822271820902061024525253729687418927203841733656345175734286917906729775369402334595843655499345300272616160911876692198669168411545145961111473802484706787415031808;
B[433]<=2560'd2000610589549994062289857177190539379137075629005540124183040054452758291095599674164031242406241988930185514111832430317539098219622546527700194149018802847157241882927580211789120109775015627369998748635164193879020382796399075399342689107218627833478110011822949621789394861890948072703190152450839517710154289363380640289553157202754345801107212450301900891765580368545178206252800015191802201642771505331086309012469104322498253058852931417255255665174859668320174147410869828882709026420995289819054589806884821735633731016537984762507291066912297345730188329213264555099713833477785008472064;
B[434]<=2560'd124125716511805493136071219538922243603246833024209656653711539214556179707501950463126304854110668275028613101778598411994161898974202255625634976615579248996578555305558068202398637435573549608566365464516716763695983079260019732484739389076307960493473464310954587955014920922980494030943533185717976845674442539697887684281736660169875917051152392625874327439201164817441701305017872255213365820076095146830687906011951596863454941869247227944935919229003571437845071519255139643090769548948774295202815764409964721043436785602897306952641596492115992422427539745082375673374868254988336889856;
B[435]<=2560'd116795794913119249769295683404946229079500625545310828963074870141971129648805333384512800486013709580249923637156529434431655198725644762616348902854169962538078656085032176836762880817135108147697117484643775789076309115710713502794294533134410631518945731488535053383210129219577284546605425667784736987253195346604910184837386124840758173694446680769995244596933355903554580979870226607527850804675660163360353020394165560653512947430867676675369405614242104158662626641105792164117705791514796915265638177837845067784814398885857290503210565996619591381880277131199540809696103913176092901376;
B[436]<=2560'd456233573971928566894565770248657330766841029366032781227932261803367994460965766773100602726503777947816650918247809546481000727148185052077483190870906352733033270697889462198752925925274236879060108340436951694076494243477145648012995554473434662343200673116297747638271054363616094655681385602970210766438397693996623014417177006786064314369573100232873869847475341607926597851387436457791723479989055904174597169468983819950031402531679543376965257925552223923875871988212876414272841978235399215334726144087267596045502365320535016133061606581144547723492608084974515903969331542770057216;
B[437]<=2560'd7398363015128399884669230311707644889471426425959388266254937342252123075631701528437094807517826366948308128339437000883759789899211841930440438231253765851412776712653197652494893932942423491741146767846077049699145655357286444137853446719753484754791729688294189596342045770523227186207559653695475017135451293270574937514875190133034886944462603932836993144189919951922247108431873944142069841066501538034984786035995392525942720476588560113390696905655176936659943445876355160944643285470635710748219347506628981580244109391445038325836011085281751679490126005694191149879488407404544;
B[438]<=2560'd27306917425803680745399532359653921199618136512962453048781426322097956826706650143635562554371720260976191303055737574515523116112738092892063787213120499983812147569979792676166449863130487661240141831113732327570120775922117716322429264883783157860806691729226497567571789310986101540331166881222980879392533145437189548782891523723235277666681460239804205427634903428525004992015708452733247185446785758582841060762649890668606544329233587501199496435308495382282277740012767963625485783719619443643050379599792460652730850898092801924184359378932353550085681613683249248533601058816;
B[439]<=2560'd106252919470556801233693270090743885491106286213760166912249898509334833706519328435180739996815985436180647373630375695243099296585828671047959304419570206735711721509154483144612947441146617690328182169085481085733723888652537645084600864258159145050930868173662976823266661382756196319021479411263947043329548565611621217337527317471560447414132328685861512731503024915310241701642810618072250913171402345890813947156045715443599843143808416458301330964347794108295665542610768691198871686685115259772289717278864935289710467725163385863494128266386209937291316163403206720237862912;
B[440]<=2560'd415050466676178289241786203694770249443489680948470733538432241950974692702771187923898441695630065314322883802024446257977645580352091709997410288851237297270948410129995018986738617316887617094715594365738842089099212057299003503487870301020815803903959868113645360008785878076346132786148982038559661931238392688733090128675373631276565910207778750372936694906339062760014733291410037619845972731952567875432242552597520222412758964832260373294534116014756713287302407515054675288894231185812467183566641576319124999607760380955944403504280444418332832983817360196300874266443776;
B[441]<=2560'd1621660236201928286499986123289647117862803171289590075386996852052515707607208425049582276581473263455705058004193654448948445777490957636525795524848407505815634063486603689256823900211496589694621202639732778413905899758637521396393287123533319522386560853123547546244455114706854877998326429840478867923840826000710483497586824156636563537204870064687263188229516219230879752931192220645528344570737351546506680204126875943543757950811678272346160039371974933862943437526651603103672217925588483878629925463247613624668491373980794128825925879084932302855072087600336939778048;
B[442]<=2560'd6333161107380288473492103209174136892863661301320424407503063628314557176037370729992778533454328352456802155704634097002232418063569548708112971742529888058696341092063188840900522330230432205825829734681240392399553765647316224291629374429255003048847801372995527879938458532468848548495583362887223285927606778145040219281919891617130342039153308023743407079329522914747303745039701010816751836885950104407296726428949352141326116482792259273978875850873060327594703539174756957186449052323966996684553604212176725356308095569037482084510700797767677774769809897722262585344;
B[443]<=2560'd6331422155892634360270098696092531291624822516333409922957531893942554854193272668733530297885565687904361978176569105217588662933137079232545654121052541368827162643035588880502539965382611233014811592443423135420728627425174721869839048561484412570454604186050075123871843584739993999121933862028093089705188784765644848171540399310167248771169368621714409828985332864919404110150891144950748228329757611548177024800340894845123041814356015958552750084880008540483438167319172099628375216288626464936817438377495342488894161295425311756895275127534660112817481630634458742784;
B[444]<=2560'd24732092643836218448717087237330820698612448024611148978727351061888391795310737713264261674541452721441795223620180090737628818038488129154467242974767881787398462458611609813492453290037348506985266329783479457740754391247143499183942310402496800748286979059026634263474524932005726188427793409229298619478585909330718311842512055476133522779355704264020655995329339655631306853539173044960658806144242209069734853354631283165392074810013558042108643229827617041933517348040560504485958113448884053033990126011510079522730974533731821589980856746361688241680530245196709888;
B[445]<=2560'd1468387807174999947067579053373722106580037753082625660613209150308299146532598150241317050632728977857331014375712641692422247265108141919184077429336956643159925585461025981624458293407677494802717067916004496654163993857384594419987024567674639242476974659020215779808769791463920206522650072037032223993148019705135546751693878562606601142520143576818819416427392293875615456069473329671393508732189000641488273329337307307809197968209726899860785444109800787127468578230095773641635793917242799858081112356826468917067859165146983345418711560751193587704047599616;
B[446]<=2560'd23580580668163234444085240092114506121523886107087525370647800699088975667353240394644562877576083080072362574232783859278518281624477307947869067184948646658974350967398005717979017860952558257061436948078768756626575061815844613099666769907949351305011558053801938647150132698676940533306302106457815266993674642653756090209241233200680856351522362717877697611768732350760236118907846555518272802315893081852123250476735458002864624853697212879099224638019649380189598574187299325014496840470124053964278025095937177893777989248470730128753530665291514989976458625024;
B[447]<=2560'd3404095678729953194445350767193377554772305394818209054158020109413036728030560691502229786231297301535950377300173248329349969560205906740852972831895066909191364981765034092045342735629559938563706579704572727059856586284143796793105409073499553203249706946188296189931228400920953535027642761494899206531188696232621501263587240926961883113713698654099745525294552165978990334427428559611454945374894648443070790799357379404972643861498985295176412028662719109948146151584451227077446466929688576;
B[448]<=2560'd3807419956475406532101045332951036701115542510027811749401465741396419878278743424312594864555870532270478706741486738797532105562499869537920430169867333492273987444511347229364259073288848194772354962190648448961297061838118391471401398145754456971236783406892430868326692318314206608480638958344965696193849656437400299376246544503021164816668012901929452341717901456609229070962659151972712412892656104914010709133793102856475779060656245831294628328610292409191986070635878893370335037751959975100416;
B[449]<=2560'd59100688741659719942749924877821584257333112056241163058458134513405102104647708504128654285546301593760068299084883448909334507017779280843015304270484241080770738343242865448300470126931394107251255798027734587858343388430904599613310586901756627471015808601338149185728800401562984381063362948057101938739346846105795561961637740139653546698862894573795507836801898330166087274512904428559819835463152554352476990038174648152383642149452724393070765640199721884110470775262607929327105085212470822884710422784507905;
B[450]<=2560'd14624524117821039677256367059490237319380646047238685368429784868001898463734153916609127700720873974620968313781895460242019273484123220666544525182638352547645911917807790950852696540890431042227791811266011771308783321459996528727155847700582626139225911078894065080433737255735623958035961742512892666799910941397544174153307877964153500040976408304711230254158054236260598499459600342356098751373102165319391647794245622621261816659529995471925595656247388047584440297082998449253760992574302161542840320;
B[451]<=2560'd4061368421194579437567560047135901422245973094860309456605505289793787599938680848989772930756819129881745804402733733548275651011092921060682120970775010799278814185060937471618982609375822600155012280900289660989469042435887832921251214561447476002831616718480205464066979771585534773627829693594953869332332827272984100695140031900153444560066979434917108920795738828817888851570947046212734579305746803061266890529934181023982305648738335580930421020335642206763752581658849682824222417325308539293397654257610820358649151488;
B[452]<=2560'd1057906232813924660752511189917733576172294503334185907086002986498703309903388070524052322245836536623245074796683122289277605204639909378357101952875300638603507724113775151827066001204387811545698257702941082617838962772838454952614930157451542272055961726872097402512361236226778175421054036684034674513503864115367581159673401926642923108665496603471149218399641087982770952492577723861547209967656781808912951719044431779308896067144016260677295884887400710458173758702278952940963194603373321576475704479928343804772352;
B[453]<=2560'd1104979952541304111038417197626446667439481177524809333230226897933955412163091797319302720083606345723098653183809860562426440960484927352720908489154591371191389959546072146176141926755944013262811476603769634866967391012110919115636972356430096383498059038082002427626857348450747582111620067718746727855597514704902895491029647163740771382691435021510876628931276819715703769900200315672082619199579802705433212058168335807393699611718276159355098390398025226230957287668157811653907952261476296242993300155149143836636695494656;
B[454]<=2560'd1044345983218480729687467758841778890240210388523603063683842197285741710099658298764122361896617494697725043230039835209422400830703812647788374169336294672128499297077143998941615557497807527359197558140373450546931144322185828967856910428084644653255381590771214964434763912722157508253952627616524972764452131805368750334525767570889418089644796759482878001134197114025044575586545760720166000406834482038799895764925777101426166950456521249747723174051452037170828058655500913354745556929815389426169105316207628471432533508096;
B[455]<=2560'd4889444834773350727970927856762950601011131213187756318634190728266983301734138803771683460002539823248871384633975998702720666702478471474105338089394870892685408660212694579398091726744248091971355984703640533654868208760184991223689170397270216258015645848229634855786810979591243181562821525189083457261879748078871167006603285425005873445531916708584391296217863403636656696793555488242356201413074744000081738902709437617592918161230225244698599847142732199478330098633082929258887504534645090450537036540037327138009907200;
B[456]<=2560'd35532923950314040371555233996418615656447617690238539146959371986022792206109678041799221488951283430456014754938233744266582558224172189085871013865500498498907118697460000900058252692829444547957332045328413014521689407863938805410341629192057365368890109778500554930922573071833010205103659946557526948495399908050295616591672457345343194686373971226445887948692820862572106913373574766175859371754302257453488041975891127972226578275030048629901981605157469425742802479364165313833308347102684519865090746045046167182925002621073876938294923133313976514303154556757746635214254300607971499956245637792070314612036186258014208;
B[457]<=2560'd1109565847988063696224845352873564437740752949623496227822692462621524836530211924974680966850216832901387650706957187701203820925171788058092251780530796624470752817589989881936317610481588862676394708303399422503522318497657108201084876503178834828805578537026517985474938764700679041583905587826546584682597745752887150225596825513900477440098656218721715220892267818164293746879907536540899048765619276698530745588548062733509608845613737963337180876586042234868184295600062093015125216275422220120441803315535975666566108807168;
B[458]<=2560'd38255062034877977026177430990952923613463943870659685930130103617759745372704032637476828005426439748524180888007875670453460111263669772904047693340057990799911178895050649262958455479373057822731656893750054002814924384903448855704194997568350050711274871141433994239689221031535170578713176258982274891573520673222003857689470752895932409276548616629710070452621658004581266482973299470515147869125965756226250871673055537281763692155014625099670024432417610399870120614243227040710826780834865676706434971272315409133601221363108458624092249421819204699789868906261771233920753425771776116408478934540379578112755630080;
B[459]<=2560'd614463660781673250365106002283749036033562724732187758088802563991857915060418525501427928489607968127247041478034983017801875056637059141227020814410111718555376336039338625383955145785546643676061364710015250263963015517660536203750500590968760496993925096546935910023338942818120138815266426659363604710196922427545518423796913807718336761512931906249292989460242350588492623574668622276433296197008201090576260983664813654083012670134329079053956198230934015717357071358059129231494258554238557059446286151542652460397520855969501069045367543729151931635389916643997041541591308446807135517679546695197406209605407604736;
B[460]<=2560'd148053840968278043675487748069868570782390191710724277435355876923779975663270771449753700894474177607122735488698616935222721316013452292064184104000889859413355673947174235269136521262670216087466243416738024214100067543868455358191767404861728447576018011618731925805533967487139417475244082497617857419578754590678608912003601167815325173892806523453324120503217984429315693356854396039233162184912500630622436647338574973662195963182960787541565858118838077309008938215564333838893421793410219139290279326789326388147153851208948337638126456898563803892796618413863559635487743778122378669738080554813352574271970319794176;
B[461]<=2560'd2386751587479084783067464634008171421557021195198603656518735358348016781620299735265953848423155179115930140943553938029843353983896682011585063655478525689476423859381859986783100282986498650302541491599250216431075579978194643848945277448271732191865926683992113565907319798475682690855187501758080354557531470186657701798246266882321123730267626851738414780411399363808846173636030456830317770962036011972607822281554934321019574132491628750391091499564170714304553281534768647905457340047945071920238054796970194680691945193289046668323005409793140152529508522619216522976997527427907807475821246135507426446450822918176768;
B[462]<=2560'd841936398104496881132935423046398685275229286403152049668558544893480021002839700525751375760954307627690336016570167637935520443357097454760057775738365821362531695111620736969727580222167890992337650367841149785000257700401558718768638321087751579745211836606976156540240304042183724047315666420426346042272482305208206916051046352846961470636560775488233712129185511565280127884789555138922970705712429087764966292033633692527030562308693310396781891278151004613163733591436242275648175722480511222991108041518415440496295339373653992343383742321268687886510943598888867079028560808341299318507156033944441832125589585438099093136605883298747470262141072517954020573184;
B[463]<=2560'd13523808992651798873823001222073777849446997989673553648465361596418168648438443223972667443404837465696653277170851089602721564966060818140334219443420943866342761897007010230017343731758589194245170669653458336153060977852566989109733791960081203283592390946380085140344545505626855605692995921425108969459352165435380870953884680522073568298418129457742833441912762925655686701129431145235603557781689823695499904846336912640629522599499491004354023907804515667285270618582265438657093948946128932963820817085113147419809796352349701426757322730878378128811411127930255790289351487050427443545430220163663973305755490671584000884544455650344097042959442179211581049602048;
B[464]<=2560'd7024863791154628036614424982945651049763186181362448336321004134464893485265312901412722365035235431798031615811684711166928422262068303475427845913996289055747463839839763374802428806662759225603692159881466484408296272069972636160539748598865460264094868967658891938600935134267741205214574679953056650144811996488874117696231001540311874042979938110987074772540215927135837373848636625350978078665190630145922194517968147960592464941663814181012622029607607370107599820841022308200461047519514544136948322813783635697056827265200677977162729957791734304476898468139427219643945451417397952163451356003752352450848583109574216658618373933870246246191145956825905424337923952191140450542809089512895489579420570671019691183886312340939853709411679973316086918545408;
B[465]<=2560'd7052405550912491353564068444622593558974638321640420593141894269817937695146099565384251062843788570519763978071177184905966148535842517951974185830066757542975873687009736140551750691888288385583111588533466816822931317584104815885209162129237317033070034751130692397316548665206175000804461703802094724860344821364539039246928477631941250605837974623839005781065413476266905477108984799839673781931296060037581322501288905583719753037175567242582537013619633016479520536606991800636864422905687146055964197044863912185206983048366815767656635800773378615840248999703184050338115373718342068121149429645664077468361487232626134379149014285543553951305265387761941790164292354145382614399233848738523198672185141690082929723285971847829918499698587695004801314062336;
B[466]<=2560'd27187490095373768866656252185663885462697105390340268912996236962323234001038299727695846890211354490043333180694043575367443350060536738963733150744583665147575346138489242405936064100247751883775497821036550072476488978227200617378412976145921740567841545903233687191819378417830746024889115842654259628683404488146723535026046661541778508843951584050270970769722529334302864611572300219076535673967088548661933749223216728484001597044670249193913798202681438924434285075728994342264310453319595029459246108350861030156154466013250026291360684501769974995208455532414896304017738223878992358633230309792884328332982752020502965821121529870068170778443020655379695072577828594099938641324610974990732570382405813065757848328412310068091160503710782045791154756384718848;
B[467]<=2560'd7050690496378207249635476162499193882185989810623667608830920116958959703795668509513248516316424635066484533185987051535200839069190870695619994922358613682071546803686754358269511898208498322092726301762234018127227814790622167572236963536291519752787108517213395430180398728798839785780924251377604896610048507888087253277622448104864336095342007120228425969390251828351959926736603256965729503137042421963837992924533443984598596843290722921035068197457230561749161169712173852702766612679022845777729339559966318098721788569010553642688732563745731754843633648484657610195339273370959891725688644889555922220208350537424017443328545612239830573003141247809620115977329005362334196320940946930848634704488185820880145234179012251487252793790043146705070660255744;
B[468]<=2560'd440668157658840634450211847747990773821109300669372193680922265138140020140244865432216943577845542486945899494021708852587240088859272437405628164067283448869288708408975913116312350051188857027343552831224010791632560137814969296412753058123788799251130083105610884822683681508146383431220533319570235276883325073051182168414387460650984788432305854497631747737546624871270224784717923030146598054235538922810741882453841177310366379856064386193892312601676707746536882459923771671605361287219765188714629281609885345934816175696657264519226785870421647162851102966246380876720087582230774720829849367188012580782650315909186964920451817998662221963810822068453587923594934887283379135961066849301343684780241009441685207807532107011140629850072819374080386924544;
B[469]<=2560'd27548065201605893895275016815092551355112543856190167465953844165510375375878170321613918423549900033987297920672303720220921201794285902519344623633300539384264430972961464159189071837886648950623241760550376929974906153466365731872478631595619555247640107945779452176064077480072978801672040924236514097665814488927523671246415426883826648747041756072458507300282048875999321152751198841303018840778344083793124103082102430181942785511315947168269147356951854139705824551574651356442385739277332175743122565756988338508736286912537029638101606964379140904361848599259383873369903186609985138885718528812191942118862424846303701662526702108842257649038179630965040530188512622852650080995390463443886768284023973115139114217520280855668471192154284602168149278720;
B[470]<=2560'd440674461371165429876417531827802870094204256056465902008988901576839948051625062916171308598357151131834561631425752138458998300447891998828306386711709837082390808332393757126442794358774087479746001769500924178699249103353353120853294897536328911656387259522350083931975546234857047499897657292501126177267673486426761462761118766778859965651448407646129236259626531468167173929812958875979920207888100280316599367946812027471599455255873684628394540957662853128528057958037421432423167893804693230831384983584793323197930196665415316493036154199573320854711464607809332851714536916073793597586431079384128328553855198768769555525100973689551487271427348641048352978308000367299430063366895475610692349447719928991403898396083669602268625512876274539792166813696;
B[471]<=2560'd119916828657152135302748932403537743094615025381481930190780897109716353445238682461886686670964511771452348588116668130454187457281287622651502244632898176473099153751968170724180608088886884341520357788056368446898079320770721328504222252077603438257535936157762251684667658452490218082221911227420628428715524209848894844167355920738590300754923803823111431753681817824835736700785413060969301200615569179166807728534655811439475274927087902754980597339007188730095152644878582290014810859646067086502435116150520158030991829363811780294200957115447590438126306385595795149947654003934311776472515608548111546981701851013271208501720235329152879238114429199070803164593615368156444733704793088671791773567512405566323918070149338485399777860960392124788269620658176;
B[472]<=2560'd88578709692552567531994696877192844054783052223455324498549479127214563286009424607940604117219077294303806868877179257242025774254921612342775361998477803604934668523495876239864228164155676319053239799642017254835178982868005502295653941910871130039433974748574143175824383915630838866810152863242525864919192769423851206424498347912575363747125217396478749593138049753389930535618921817668354888967455150844649477852076423553096715743663061601833591804378142618926822988504600105318895208252162615634407099108777587584893917860955301732507642843160740886588738056556931576950838723090587786873599402404789212572061352476379298334711582318176099806303965350486988750431716613533265675130772676106587226677422412888562401276461119536892281723410825078158580544713064448;
B[473]<=2560'd202206737131696770253142860902643793962996942683750308583543319105254822981769702796268132946164238561087553522805316340958825283631763597435511151233359262663685450790138848506647769041587359452525927237058779648360844933594178165703809320448761231703259068714294169004606818550737965761180982510858596647656383340138625035959223261867382604507874807755823789074471540987207680373979829012224512225902640058981537410775544103218081344899009381729670883907217959568407586961627305194911173978175341389038936248771403946953296031334995557653575205291581689267553931804966992606436581531179863671422038051960805935390963919451087546529427121223425468223797094577729502777413704344342888371660252641103935303854732201159988102589579843132690122636785388146795456412904325392;
B[474]<=2560'd232786022690669003021107984954579653930663622802977608384395393438615289176570733506188295287719308549319251778892840119731671444374508670960542346657462880154579154457978640469876003713956369742293505997749852937926872321464855434205473585624782701821443786720067963786963623725361082710698251781816161520823788636310170903613105078541808292253307704238760656168469119930201099778509313670064641045612945005215060517960461596327180215686957622636885036506338147718557854497833261611656256323499173709890918266717383405302772326832851496893981221937806119056421767421904432925912201737688999913463864295387896356704649211732527526052637041642464284398375951306662069751614103011401185277633900286437510746552526793725161447974729420492084813074149827206056071082215997456;
B[475]<=2560'd259973512799914427868665841100064132955334130775296493738914518023112812036433164574316971296901491207608048917976790437254888955224378051613530011747443135025592646598399904913140515501124647107622816329927764490598997601339419138457525635134713323993363947409904089635072616431711563410859117428022952210656178721170609844322238983663937379648165146621512299578964638337208456219270919822931396243756965092485982197320070622012260474364818436675356488635069000513423599651827550420084822821000073333768689736573722525490037267827321993493817423855761996828153618133516622186786394880451514941082818267674850190318922075825774559841232567060427556690436773386507158204384627229466190124278186511150958058092906941919307866616777268449715175453622981018559298392273522961;
B[476]<=2560'd231093884533947889734268991835940435075553562158201233934515684860112863254567669911303305066538767612318902486728687531771043269248765420273525232768286931932256555141189464070353690048276431956135437039422430724429259435047019316965980459275041208251021934067896300133130461931195309862095772950794469124469881628483727728540756152256734804488647494684827817445742134262936475137620869380966679818746391231754785125710406370127824087146114432573115220563348372565174092441489288025965350959192639410044585399751410447713481898966877995397127758115025532700116862477948999992457689009020599501270155252650498394932127156525785810363206527090098692237262091709762772991062942144034432852187572740159087913351560844197253056360959925613500715282156064110877959867545489681;
B[477]<=2560'd117359633464110863205513229926789107402920834876925534334911703923947725433265753532011627462031738292062282952227387643707255948475088731701125800781502889405058420219577532524591169327931991610378478837514425337148132676125251509619950406678706204720306305836312521727696176237638076305550712746421130739934899698614819567650971835505443631771922303883608500274612609037019788818727604382247930814278793614714258211292457296442060918175744094306540580471359706602881382092888064364140962206758094249003625685175962254912162122198950376442843465999898639658817004315799236457465852490000317608367922578789547766291714728237441766842547511403126732629334578760409430019844187637553132031016827052312262662786808943086719385323961226059260889337459106966323680400229086002;
B[478]<=2560'd59586273815900966936186018454575680998241954810537439500449433791868865150274677070150577161144317953513698192472312697946478636708197582740474791298848463707831170586386354806562753527784078763600188858257100775747868904232324626970174569807056419698048801761929937686367231667966839572106398627472788375977314910633239671855791561364656868058760032770353089456553444302823681608353570928808686833372522508777465406276360708615842022440851038725746780203934082230027624674589390777734913279295347956438083142744845515046209292482170181438930905271312335102561275123860641438435970319754031712514917732260690935700291949532862080776916649022927516175064778773093860509456987840759693155067697878577870829524946827188641799009421640654127107420316557293648987760186512981;
B[479]<=2560'd117457926466941821840695740754478637940381819086616500533253102861783707937945987063075407701911892458358792299337024361180259347567819763486701878339667537998096568433418217801374333376001499265036608773365763503872723311172504419501892160311377024027441335248436036103762354449690479052312958637047508217043285479524839896375587619630840327597390946738625575855649315588894540230281944863667297703176429842430230161071736515795047800701276971144671019435601074832706089769670016715834216060193195919051756729653997824106423604272832595842665602904872289009715659758599444404926798643117141059632815942861510042057939511581276281766225174759649183582900716026477436334352452640256054858584053549888708413941194635412601473430260106468279963408643069657303771459850744338;
end

//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)   pixel_data <= 12'd0;
    else begin
        pixel_data <= {R[pixel_y][pixel_x*4:pixel_x*4+3],G[pixel_y][pixel_x*4:pixel_x*4+3],B[pixel_y][pixel_x*4:pixel_x*4+3]};
    end
    
end  
endmodule


// The whole VGA 
module VGA_out_color(
    input sys_clk,
    input sys_rst_n,
    input [1:0] choise,
    //VGA
    output vga_hs,
    output vga_vs,
    output [11:0] vga_rgb);

//Wire define
wire vga_clk_w;
wire [11:0] pixel_data;
wire [9:0] pixel_x;
wire [9:0] pixel_y;

//****************************Main Code**************************
// 这样的话每个VGA输出都有个时钟分频
//优化的时候可以将时钟分频拿出来
clockDiv clkdiv1(
     .sys_clk(sys_clk),         
     .sys_rst_n(sys_rst_n),
     .clk_25M(vga_clk_w));

vga_driver_color VGAdriver1(
    .vga_clk(vga_clk_w),   
    .sys_rst_n(sys_rst_n),
  
    .vga_hs(vga_hs),      // 行同步
    .vga_vs(vga_vs),      // 场同步
    .vga_rgb(vga_rgb),      //4+4+4
    
    .pixel_data(pixel_data),    //像素点RGB data
    .pixel_x(pixel_x),       //像素点横坐标
    .pixel_y(pixel_y)        //像素点纵坐标
);
 
vga_display_color vgadisplay1(
    .vga_clk(vga_clk_w),
    .sys_rst_n(sys_rst_n),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .choise(choise),
    .pixel_data(pixel_data));

>>>>>>> 4766add3234869bdfdd226e07749e9b31ca939a9
endmodule