`timescale 1ns / 1ps

module background(
    input [1:0] choise,
    input clk,
    output reg [0:639] data [479:0]);

always @(posedge clk) begin
    if(choise == 0 || choise == 3) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd0;
        data[47]<=640'd0;
        data[48]<=640'd0;
        data[49]<=640'd0;
        data[50]<=640'd0;
        data[51]<=640'd0;
        data[52]<=640'd2293498615990071511610820895302086940796564989168281123737588839386922876088484808070018553110125686554624;
        data[53]<=640'd1675976290930685468645128323187019804819274807935478584355997288644324119240316295174021690532034581474959799140168891292198173855926923755850975816974336;
        data[54]<=640'd4608938271443963528941588642716363415553844460538933171124528709463054170393956612499412155428494782625729343881662003406464265768870265575791175453900800;
        data[55]<=640'd32262541127990939173762083020509032968594440138823179507501159485634574000849247021006776338229579036834994698149052345903902864697637648985753025844871168;
        data[56]<=640'd58240171439706361472169453622740139551676880264982424390591317149858243932624905087835037248725775054926940671759288438860704227669296539774404515090923520;
        data[57]<=640'd42318407564523126557606423241263499508701606765135631683196970909087290531237324837141462551277584976845020334793376876887606858787731732121488036166893568;
        data[58]<=640'd395530370495227042665516596148738352043683483543209051664862984962215722154818246074688097346266051782000026180473705838717361763032412721084388760520491008;
        data[59]<=640'd875906954421202713545704567525854790768358994252243776699793848151799154343056753832682919968808972452753249328458824810904489328815372625029041313741275136;
        data[60]<=640'd1074300936946527189448081477115531402820708126955742360356077044371693182696136319406376230962391213472250986774014381769145217585253263421021236472190074880;
        data[61]<=640'd2723731004535675457407407214648210750903770826922016861520642014671865412833960365204224421091120348781355315742556081222814866948425965607358914138996736;
        data[62]<=640'd5363542192147591106665945431975488483211153355654328491357949574079026346254569789205797302263463966091837288140978704750469707812894644221288083022638219264;
        data[63]<=640'd2148392389880624983854794822778637342357380469688204162829970252499582343647074513421659901813271610738497426696471688412865232369391466669779185154318663680;
        data[64]<=640'd11157393520650594033816653652288795059042270346749989081083521077635666177081536011080883761299459976071350897937465882988689764126215296351421545708670418944;
        data[65]<=640'd46340318392186936871323099658801396008038326033905033280090403424319477039293533746461577656164197176237198767912607413258782486604516713763506551490862907392;
        data[66]<=640'd6866894267813936637844109936851291657023550013168452068701946928148428461883378977066012880698571175098621288248210288500459301797733256446001671825596088320;
        data[67]<=640'd6866055871643455633919549855401627155405683307443407615500233076853761656628263449134380842739204401454157064456222742542119398180196937364232137528850776064;
        data[68]<=640'd82380932058025304369882760701860083250682292991484941806457284014125123379755651628509720405156100616276445336341233578718530541909729839781497329850521747456;
        data[69]<=640'd123568046953902601885489631601050712319174756009461312869005805972744294597349989309378349784223221026846516048020819811265697562604659577532981444669203283968;
        data[70]<=640'd288324856952856638938360058898595805306574222331048332226622281617419903733234488006034233947574894938995849281914303336068168613552865455582601091901248503808;
        data[71]<=640'd604109837461759778168159595812366405561914221390916897199734931180272979632225765748065127120840811121811655347422247737108184549641653972618942044609571717120;
        data[72]<=640'd604113173047588395015331192328821260737655662434528286280150192127775494254945644991600158879780428058664007014154694790222100112847793335065517706788783259648;
        data[73]<=640'd219675266569980855101283472340255299678830543246909919602823875385570340106129550504925267063655400482168152660230457948423843364412407532088987667975607681024;
        data[74]<=640'd878716280995473004337282926076232960710252933604169513785718377197055657451630564829885256010195180777820288365803555872444941845579307383195420644215244193792;
        data[75]<=640'd1867228394076075483794978113422141474529413092464248978844049179274668247592540852714362839805123260305110545725523235818229294611325658936654682330078214356992;
        data[76]<=640'd2196759186277915900926322250153514691466961015354738301595353246150210141478551945047509799424682666003850921931081454547645667767808867014961711369790485954560;
        data[77]<=640'd5491840118327575789266050286268835412211319625532502477095620565199695451401293084153438916689517108918215411578931448829559414360696935030298648443765439594496;
        data[78]<=640'd3295140691075790202280104419051183345307264370081109106149563130065548234442196278888186533097198155681390201425625669533083696367444166288535752857087247384576;
        data[79]<=640'd12301738147164137008516192307349284430213059126345595918172653360353590957845406813189173483570374230403960158616455187826875596110565138928530713386938705903616;
        data[80]<=640'd10983694272968463208017411114256965826893096936854354198107273535794206413204309036433666244710318396426212727686533691447454945851282655205826496843257263161344;
        data[81]<=640'd16695249082583700151819180632048177262635343246267534392840559284858924655228845405174144134607644664658356352874643028256124293023562727569268576201652675018752;
        data[82]<=640'd15816562523961361330229573309826634226434290288366856178771999537978267005376446045370118187440417277347052876463276094705521338392416505356020586531298431991808;
        data[83]<=640'd36026489125927671166289176420646080071866189211135292775156866507934099707732327272359078617095675212156124947774533078691482697388957364701881514429016937857024;
        data[84]<=640'd5272240021943069727947564190292979055793729966361248715538640052077095891112436303112593429210693090570943905958303872941466164741451264206416949289102920908800;
        data[85]<=640'd29875653048126526639798045377648067050180185090282107520280915163244183757325856740083861989077872004946784096482024153935771661077851379083361887904318372184064;
        data[86]<=640'd63266116017769340614370302764131239925710436011546193109013856643390801955703664349384433193504743177508980454909012615578815823764973452731200254228423507968000;
        data[87]<=640'd31633061360863825370210645136310830404209726733791878434705385420389778471631909814652699262398831417058366293186418192618503535676488482274630290480730283704320;
        data[88]<=640'd63266263503656570665825684773802091766755078915378435853240554166128374162234725728383526188788462984391661037890014737274341293996581484529175727360672803061760;
        data[89]<=640'd70295581671023508211478452617564891644709630344406242109297818921681604012213781017281502757906308516323092188893825690710699206741894451723342734933425752375296;
        data[90]<=640'd140591176749765437835789265421574959863756815093899739696031636517167324564256131031003711274920578246666233112393967661926318979829304773066559488652826841710592;
        data[91]<=640'd56236690588038060701510754154057083807847535199944312387298568698492464460505779782646578450388672046384196427450360965925681982269874295247584323200251139719168;
        data[92]<=640'd337418775931314434710666121368382058581550402986087022736596132649012604514048986252565250960473903116455606423577632442273831910856563706269486414050219291312128;
        data[93]<=640'd84354740910148374275949364164703432233673625957957103591082717251868282624564948702530145342028491063265353316901573768218354216004237376400809978444917485076480;
        data[94]<=640'd112473113019738508644751981776265581042538941086922546215314451586728435496034081217546402872535840442426955979921003800584349379723459316631560600633045759819776;
        data[95]<=640'd309300537899771631082660610980791466418600909513341640781873249643700485657286888528662428914250860760547729443177382375785407577796792937338398326762111705808896;
        data[96]<=640'd56236422431789954785131731391502193504346644638376045558492893439990743552035552631576808305257788610793059377749037847322670386405301057230994913620053708505088;
        data[97]<=640'd0;
        data[98]<=640'd0;
        data[99]<=640'd0;
        data[100]<=640'd0;
        data[101]<=640'd0;
        data[102]<=640'd0;
        data[103]<=640'd0;
        data[104]<=640'd0;
        data[105]<=640'd0;
        data[106]<=640'd0;
        data[107]<=640'd0;
        data[108]<=640'd0;
        data[109]<=640'd0;
        data[110]<=640'd0;
        data[111]<=640'd0;
        data[112]<=640'd0;
        data[113]<=640'd0;
        data[114]<=640'd0;
        data[115]<=640'd0;
        data[116]<=640'd0;
        data[117]<=640'd0;
        data[118]<=640'd0;
        data[119]<=640'd0;
        data[120]<=640'd0;
        data[121]<=640'd0;
        data[122]<=640'd0;
        data[123]<=640'd0;
        data[124]<=640'd0;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd24084754561361768648102764881807084833480156810453237320207177473645930965106688;
        data[156]<=640'd74106937111882365071085430405560261026092790186009960985252853765064402969559040;
        data[157]<=640'd70608395103938906748405107852975316393858956036050582890626880237652602651358048951934797737936631459539297024459407360;
        data[158]<=640'd45391111138246440052546522188883403559323054846082361826329892174494524730641999395236457398525145100652968239135981568;
        data[159]<=640'd1636695300423147339984264753165683763861352068017600084079017597289272743107056999745917197413513491481228221452992242061661815718914536385280605159424;
        data[160]<=640'd1585546547344335296113853409499099363080482373423273381883767816511650089470346914178743826280728800528865695811453009466328567948542369888887919083520;
        data[161]<=640'd1499240499469038150352069204590791393195277157356287282573090901620345529018413437819290550805642078102596582069426496683875338620610981202319829368832;
        data[162]<=640'd1432108391049830273401644278722737849120364334060297247134938174134513807501900800215425895994497321779674193266119508278048795711930628599338634313728;
        data[163]<=640'd1432108391049830273401644278735649098510798877008576842994953233506200279217848201550508752554026776391740998501303430948513796217162926072429574881280;
        data[164]<=640'd1432108391526171299756013210551876448029150614539138435787030598275081770131852063681093028035848772279035276784484252021983740776745069051870915330048;
        data[165]<=640'd1432108391430903094485139424276427473980435159081327369931112343416947798816495883946762667839777955560060319458886669030369564042715836043895660085248;
        data[166]<=640'd1432108391145098478672518065078236569389773955797441806254956279136580565305377704354828703225921280575948257942322540404950830814731467307273244639232;
        data[167]<=640'd1435304159184913523730074650705793697101542978888194795863711066188827681739786745161951189230623421175438922548715131793750926613889998273988660297728;
        data[168]<=640'd1435305037367229710644637299496199212568719915731594059278130643385491741978943949843963127844319033508265347311733950057284828604547490761026662563840;
        data[169]<=640'd1435305037367229710644637299827448417961298273229098846927417863473669561179014619152488000536355792201675587252827406296687614509099521024827229995008;
        data[170]<=640'd1435305037367229710644637299334373618732349678270996364183221587829367760609145726026744782561119957545428387402377148278373136728610751125342621007872;
        data[171]<=640'd1435305037367229710644637299993567271371739555789304069914834457587459522536104288487695019206776728729846866371242131408545259898951552500600571691008;
        data[172]<=640'd1435305037367229710644637299333487199138825454724606894071476206184202028858221877983831414751630822537736703386206619778425774892426268893339512209408;
        data[173]<=640'd1435305037367229710644637300653019438121440510868069007907168480577641826757956539973854350149827416275424392591229598479304825936053175413608078639104;
        data[174]<=640'd1435305037367229710644637300653034558641143412569597725777903431964866886898193444370075328131673110808604221924283288817759997577909217358664431566848;
        data[175]<=640'd1435305037367229710644637299991983623461348028344010791960645046074374778705467357024839583392402874487172079292395303024722442452133379642409980264448;
        data[176]<=640'd1435305037367229710644637299330897443181561344417431113677107966919478585359131666779569300610786589534507938519752671279255654159513994981444495081472;
        data[177]<=640'd1435305037367229710644637300653029495482915038838613054143659807267775516853193537903920654581336503892994637717971373035093841031522860826515937951744;
        data[178]<=640'd1435305037367229710644637299992114802589490987460098161908503990359874513499613344915043052155791646944514578423600700997597789590847215077138546819072;
        data[179]<=640'd1435305037367229710644637299828787438695083915449891531911929626210393274776978887610931890986492201089081971266064718119360062608871443242470722240512;
        data[180]<=640'd1435305037367229710644637299437092528518306659726087176161919758242288498105904759736451027421619171134752812288730275521880220238638370174373946458112;
        data[181]<=640'd1435305037367229710644637299507781500724513233078128733369671170587125172353968989771482801333236989287052402859688069010439927259458017806736643063808;
        data[182]<=640'd1435305037367229710644637299361884422014369541227848242073100429670977541832460348276643557836512441370962158324081713487370893782277483959604217905152;
        data[183]<=640'd1435305037367229710644637299330897384075245286961408227572008944085624655223000009162103830482396664431885916192872312702111210533470150330521170739200;
        data[184]<=640'd1432108391049830273401644278720155599242277425470641325827208866944244833533092231581146358403408170107056582211069222276026431019298813863888485875712;
        data[185]<=640'd1432108391145098478672518065078236569389773955797441806254956279136489502701054623304629250605004095551821760436168061530485590687033354070162791202816;
        data[186]<=640'd1432108391430903094485139424152479479832263546777843247541066662367902466614407770004358331660552339384398933352360265046554038560303752771291930689536;
        data[187]<=640'd1432108391526171299756013210510560449979760077104643727987848138723016573772462518240338453399013185499578619903403200659780537093026911160143901097984;
        data[188]<=640'd1432108391049830273401644278720155599242277425470641325918728819289000624416960959470002900423128542097679766079649740384620074055066005399296163184640;
        data[189]<=640'd1432108391049830273401644278720155599242277425470641325860322923775538239351472084691929209789460840314490041901410321420731253428251615359605793619968;
        data[190]<=640'd1432108395908508742216207382982285076764600472137465827655363918997263672051292261884593880915529765509542663695181323129311614392245719303451800764416;
        data[191]<=640'd1636695299851538108359022035016317859765970218969111736337295113767801112561132908262865464095900002411803365261028630529618247886460062426035715571712;
        data[192]<=640'd1636695300423147339984264753164803680650949400929914618905344030551094012883161424892461219733163082806729873652110221921477370731085546254030396719104;
        data[193]<=640'd0;
        data[194]<=640'd0;
        data[195]<=640'd0;
        data[196]<=640'd0;
        data[197]<=640'd0;
        data[198]<=640'd0;
        data[199]<=640'd0;
        data[200]<=640'd0;
        data[201]<=640'd0;
        data[202]<=640'd0;
        data[203]<=640'd0;
        data[204]<=640'd0;
        data[205]<=640'd0;
        data[206]<=640'd0;
        data[207]<=640'd0;
        data[208]<=640'd0;
        data[209]<=640'd0;
        data[210]<=640'd0;
        data[211]<=640'd0;
        data[212]<=640'd0;
        data[213]<=640'd0;
        data[214]<=640'd0;
        data[215]<=640'd0;
        data[216]<=640'd0;
        data[217]<=640'd0;
        data[218]<=640'd0;
        data[219]<=640'd0;
        data[220]<=640'd0;
        data[221]<=640'd0;
        data[222]<=640'd0;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[232]<=640'd776790931223330254907009681665451926923432634146589683220239250695842456566297925992806072473548014703579287154640580429317990534798152161039138947072;
        data[233]<=640'd660112465837955895739221196300032900889389781067498077708454946475114253791749433487388225928158669858709276934759650228460064616906766016298279239680;
        data[234]<=640'd716054195715451547242569712078821989794218681978577542941493380638397682223863664322544223568358465496659348510484073966487713886108951164052813381632;
        data[235]<=640'd716054195763085649878006605271096505493162353663964368912012892892945166105615811211600999073734541259072868665551139018036680509270078572746034380800;
        data[236]<=640'd613760739218697113804657534100821921254332919828471363860652161097943258383094857179881852931776215206652750007736803826650701570673207073343417614336;
        data[237]<=640'd716054195572549239336259032596121955099334801158207852061356801448792842080559168270882818182321596549367850604942333938021886517261835439313086578688;
        data[238]<=640'd716054195715451547242569712158871736014912852844908269353886756848687318187997569458551373113494279167753218908851100250178044746260928142723719888896;
        data[239]<=640'd613760739028160703262909961365203591672173316149811168137838111293297354117583164902912030002727744934092442451961619166581540213446845762221897678848;
        data[240]<=640'd716054195810719752513443498454979356758800439428213205417422927204079958898775110336209128697962308883265212617858920508814207947400500444495681159168;
        data[241]<=640'd716054195810719752513443498434320710063628303715722104264378486736449078009609937506835143563140728989218382396221405478484941207118017931440805642240;
        data[242]<=640'd716054195810719752513443498506624652298210471454580631817978684638221256651682055343100676463891433662762449512291550250352994498084041687198964121600;
        data[243]<=640'd716054195810719752513443498454979339520422719331634086085317577553004449140326088157082167534735801866357466995654626418694858991575285603261409656832;
        data[244]<=640'd716054195810719752513443498475637968977217134947546067972745522638726218803218737963866474074639029707315953979441524666868439552122893476093667311616;
        data[245]<=640'd716054195810719752513443498516953967026682825744689537321206210830870755031356310792626601131510055948434664690725965774794625032834905303444631846912;
        data[246]<=640'd716054195810719752513443498475651838503407857783457612004023740012272049318143742879487223216607915566096410483134765841002218758775178906054867025920;
        data[247]<=640'd716054195810719752513443498516972889851300130421028016039157347335497661769359591841987425384638752091307413007997007491500789825376896002756962156544;
        data[248]<=640'd716054195810719752513443498477129571367123143256409622961880200894187855801381105167642950423942030140195393554408533171113187586288060610244853628928;
        data[249]<=640'd716054195810719752513443498688349581229667683819234323872614482215359658453377902801690390410282977332645815467658880462739171969499039438989399425024;
        data[250]<=640'd716054195810719752513443498467889978237535413865193261722516837795240857176937423000817673609967888972696308019079950730225735760304001403993255313408;
        data[251]<=640'd716054195810719752513443499012744682755095901190603710942458311937664230556259154779137599693269315475229028829709518779086258855941445733184438272000;
        data[252]<=640'd716054195810719752513443498434320749542647963546615847128590290717972407571799454286011043581789429640321044974277537475434800497574688132935473692672;
        data[253]<=640'd716054195810719752513443498764848812664846345737906278997849975982598580447173321169773869957056320881961665510260061692698207071969379802162304909312;
        data[254]<=640'd716054195810719752513443498599584702492099270351629887921327346536436747285995343650763722514606921429714685427165654562488330188806306396538197245952;
        data[255]<=640'd716054195810719752513443498434320828500781206688941497732121774492216533516931710521477415365599104042734973635925821243467354688783545621977073975296;
        data[256]<=640'd613760739123428908533783748022824438419078804462979289892749333281482296153378453386459831809598151032801689536472321311761208179628544868692954972160;
        data[257]<=640'd716054195715451547242569713067823772213345384943196004009009088356959474312158081546613895513026045545123624799960285426309255936814095547164780396544;
        data[258]<=640'd716054195572549239336259033530702395488284809835556403921171256902278259661830482876894470727609808971837699942243493575529123185142255009438730551296;
        data[259]<=640'd613760739218697113804657534711433314465665878071032689821669780823587264776888397084705101346608823682554815902795910942811073993053114987340172886016;
        data[260]<=640'd716054195763085649878006606577392162570678021919213997529348213847026587804420199614273285468072257559282186656092761864256846949472257882743004725248;
        data[261]<=640'd716054195715451547242569713398351835412481939453995422825402414182293085580568833513668095081506865077682764765641214345568902369610989501851463843840;
        data[262]<=640'd660112465837955895739221196294868401133216110672097662729025665818992141539655197441886213985069293820361315308564429184927505435222358720396723748864;
        data[263]<=640'd776790931223330254907009681665451926923432634146589683220239250695842456566297925992806072473548014703579287154640580429317990534798152161039138947072;
        data[264]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[265]<=640'd0;
        data[266]<=640'd0;
        data[267]<=640'd0;
        data[268]<=640'd0;
        data[269]<=640'd0;
        data[270]<=640'd0;
        data[271]<=640'd0;
        data[272]<=640'd0;
        data[273]<=640'd0;
        data[274]<=640'd0;
        data[275]<=640'd0;
        data[276]<=640'd0;
        data[277]<=640'd0;
        data[278]<=640'd0;
        data[279]<=640'd0;
        data[280]<=640'd0;
        data[281]<=640'd0;
        data[282]<=640'd0;
        data[283]<=640'd0;
        data[284]<=640'd0;
        data[285]<=640'd0;
        data[286]<=640'd0;
        data[287]<=640'd0;
        data[288]<=640'd0;
        data[289]<=640'd0;
        data[290]<=640'd0;
        data[291]<=640'd0;
        data[292]<=640'd0;
        data[293]<=640'd0;
        data[294]<=640'd0;
        data[295]<=640'd0;
        data[296]<=640'd0;
        data[297]<=640'd0;
        data[298]<=640'd0;
        data[299]<=640'd0;
        data[300]<=640'd0;
        data[301]<=640'd0;
        data[302]<=640'd0;
        data[303]<=640'd0;
        data[304]<=640'd0;
        data[305]<=640'd0;
        data[306]<=640'd0;
        data[307]<=640'd0;
        data[308]<=640'd0;
        data[309]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[310]<=640'd204586912945874764240387462872684461939791862714291309128701634107400620581789783294404734467263753122353208725382371822087818297065713413500142878720;
        data[311]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[312]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[313]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[314]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[315]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[316]<=640'd716054195810719752513443498444785882909390677394503417248096665387912638568274816216319923546195994976306584519426322962481530122975535690971336409088;
        data[317]<=640'd716054195810719752513443498455968487483977001750781907060838224134704709211147073704256992800668164780831664868630583039747908261161583167644333244416;
        data[318]<=640'd716054195810719752513443498474537234532114649602277376614592304150941807458703701962780977343526620605754526330208115812089993145710677900868284579840;
        data[319]<=640'd716054195810719752513443498469181083417895511379387966348654761088606061502328738306483090926155365809885569869539490452204505213097378866499214639104;
        data[320]<=640'd716054195810719752513443498460143208844760463077529821080196447904555248326788557900137008901452003884198374928910000939410338251252270873223882604544;
        data[321]<=640'd716054195810719752513443498527281705674757012943335194389606949037152868359891240043216593653491645666403208387701926563269058460469809487764755841024;
        data[322]<=640'd716054195810719752513443498496294707137714219955397731849003363864599373346113716124368161452497813606465404624444234571178191844129520710124740542464;
        data[323]<=640'd716054195810719752513443498434320710063628340411699960038642707334417784651430246326352683510526311075218355571800711260941025649074145058756830953472;
        data[324]<=640'd716054195810719752513443498558268704211799916019206224453643091529109337873841922197184505931979417130605302723257670802630712437700647551437725761536;
        data[325]<=640'd716054195810719752513443498516952706162409451976667229383883273086102694855356451481973609612325014781178703990715379981662365375319896323895735615488;
        data[326]<=640'd716054195810719752513443498682277239580970957473452572422737403252585741964642850032475924422476581956582228806857619203036121907734186946087295647744;
        data[327]<=640'd716054195810719752513443498434421638533521882075411746585902044686871280811745016078464176196770890654219677253771343330134798667677997582164607107072;
        data[328]<=640'd716054195810719752513443498520180528360673233561419094502815395445687106779796414844980695166071443563498360276778173398667954563354747162810074005504;
        data[329]<=640'd716054195810719752513443498996605656726023935176777716230020742777013287689054251465974486966298616100244663611899227079591643839540565529680693690368;
        data[330]<=640'd716054195810719752513443498573762205327292022636158609571585341487229762413136362358988649101210667449267486323672056625660151417107876774568232222720;
        data[331]<=640'd716054195810719752513443498682216713136626426241962318096820975062643994920880194237175984206851725341056316457898984997855816749784111530799062319104;
        data[332]<=640'd716054195810719752513443498599584702262693814274499031200694035285404404923758357194094993893866283716026817139533485184985118062016148369030003032064;
        data[333]<=640'd716054195810719752513443499425904673101307019081430866693741199808277343705677208242846533457381245478574006576665460295014574276902122092042165157888;
        data[334]<=640'd716054195810719752513443498764848716623583836033777364462676998056899305882677914285810678489932238168967027307797086834675354174885748935025999478784;
        data[335]<=640'd716054195810719752513443498434320870134880584172952545574899093982716409234873420460666315864822867744868192177266560455333762829457981149911869030400;
        data[336]<=640'd306880369728433813490920999973032091888177539338973819344566951264887624718129768309910498613285543059810870937169556231544353114825081807705236045824;
        data[337]<=640'd716054195524915136700822141345505175867727173326085351914563933581537959374124886357715011359114410977876207797533991045274121520973040230082134671360;
        data[338]<=640'd102293456734924946615096645243179359725951523280409852558940553728898963952424449823390596571164643963785372080723646075007308202677695252159801589760;
        data[339]<=640'd716054195763085649878006605965398942080639623315187204597609793783644828853910759009133843173107130558328372115095816278527908203806702671000424677376;
        data[340]<=640'd477103080205620143594376346681221689084677641687696716643995623368367979783064278499825532192613900514358981828142414339007477591187015844279068131328;
        data[341]<=640'd40757545357465589008840466789133681118391266897917571308776845053923947707004850323457321705794696241597790325850590410003784231118969220988854599680;
        data[342]<=640'd380403801969710437049663090959704244799164306710836292282002467361635696256651293438701146087377121643369484786329698804929741386998927764517787009024;
        data[343]<=640'd0;
        data[344]<=640'd0;
        data[345]<=640'd0;
        data[346]<=640'd0;
        data[347]<=640'd0;
        data[348]<=640'd0;
        data[349]<=640'd0;
        data[350]<=640'd0;
        data[351]<=640'd0;
        data[352]<=640'd0;
        data[353]<=640'd0;
        data[354]<=640'd0;
        data[355]<=640'd0;
        data[356]<=640'd0;
        data[357]<=640'd0;
        data[358]<=640'd0;
        data[359]<=640'd0;
        data[360]<=640'd0;
        data[361]<=640'd0;
        data[362]<=640'd0;
        data[363]<=640'd0;
        data[364]<=640'd0;
        data[365]<=640'd0;
        data[366]<=640'd0;
        data[367]<=640'd0;
        data[368]<=640'd0;
        data[369]<=640'd0;
        data[370]<=640'd0;
        data[371]<=640'd0;
        data[372]<=640'd0;
        data[373]<=640'd0;
        data[374]<=640'd0;
        data[375]<=640'd0;
        data[376]<=640'd0;
        data[377]<=640'd0;
        data[378]<=640'd0;
        data[379]<=640'd0;
        data[380]<=640'd0;
        data[381]<=640'd0;
        data[382]<=640'd0;
        data[383]<=640'd0;
        data[384]<=640'd0;
        data[385]<=640'd0;
        data[386]<=640'd0;
        data[387]<=640'd0;
        data[388]<=640'd0;
        data[389]<=640'd0;
        data[390]<=640'd0;
        data[391]<=640'd0;
        data[392]<=640'd0;
        data[393]<=640'd0;
        data[394]<=640'd0;
        data[395]<=640'd0;
        data[396]<=640'd0;
        data[397]<=640'd0;
        data[398]<=640'd0;
        data[399]<=640'd0;
        data[400]<=640'd0;
        data[401]<=640'd0;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd22835963083295687686091080188131599678433132544;
        data[406]<=640'd22836137307867241909738992724944393428252229632;
        data[407]<=640'd45671926166590717540745122690701737417425027072;
        data[408]<=640'd11425168305238367630390631743024032890990100480;
        data[409]<=640'd92102251995524685136327182220460836482002714624;
        data[410]<=640'd174235205715414699939639567012653407666176;
        data[411]<=640'd79973270849186984475343595013176781527727472640;
        data[412]<=640'd758237586915271256831821758006986185344286720;
        data[413]<=640'd188399493930006087410775984133357220008931885056;
        data[414]<=640'd10634488215193846815244531305132589056;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
    else if(choise == 1) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd0;
        data[47]<=640'd0;
        data[48]<=640'd0;
        data[49]<=640'd0;
        data[50]<=640'd0;
        data[51]<=640'd0;
        data[52]<=640'd2293498615990071511610820895302086940796564989168281123737588839386922876088484808070018553110125686554624;
        data[53]<=640'd1675976290930685468645128323187019804819274807935478584355997288644324119240316295174021690532034581474959799140168891292198173855926923755850975816974336;
        data[54]<=640'd18016743004716045104939568706166646234830913194566828459917631673408091544086843037861291450401948673299982734405370585939836303642089739931020670818844672;
        data[55]<=640'd42318397475031701438889607385923245877036691254239602651234569147285240898305566161081713485969712312403657740930550414975923248456038202051341749537734656;
        data[56]<=640'd57402183344188992557480846249111134803883445987125003633414363911957637828907724366345008656219299889741061112297913938112867822288523357300753250694201344;
        data[57]<=640'd42318407564523126557606423241263499347310989384703844829702022658899048385630712785314992999361375193054543958740802212534772278779117267377539787870175232;
        data[58]<=640'd395530360905215115021967377632711409942006648779440471063266579816800946473045629048871445053568278627989595852987097636404105016876635012054155033330057216;
        data[59]<=640'd875906954421202713545704567352562934563026676853642611817926797221644961654863567688143481820911674474299584801504605189711145700733634866251699676946366464;
        data[60]<=640'd1074300936946526427302439310125071297515937130994533697009700542908227236054607196059323136753822689742996809766773833370569381539617161493151705275232681984;
        data[61]<=640'd2723730804743768237183904232934132161590198535360849222019756894908502785821633132584250944977698014866267721515232107944067370552804837045185415225540608;
        data[62]<=640'd5363542191748007292225498426358644037797628068518507929096833266769054255422522206636867302888064784899710315832520857566929660082277303334339182503433076736;
        data[63]<=640'd3142916103311877827994774634041287214440824010129971401946070220615944633674407965106679014548230495399058990158957803742790727468293186791713320095186944;
        data[64]<=640'd11157391883955290085745718645693946645242694238428966059551126335989982129014637808743606319664413813119272322494123819208654259517587023408725019044406624256;
        data[65]<=640'd46340318392186936109177457491811105143390564853932790665686560000254254661569666650423555483369856326553091574677262891816660630792352920929528114164621377536;
        data[66]<=640'd2096606884159293981315126535532627615023078102265478175759719763157201612263761929777286175608312879866159756539412255745900722075555602617940478057775104;
        data[67]<=640'd6866055053295803659884082352104202948505894945454718108404934879957895628581040891606397478280400890069828080887171596984391567232311544567374210143564595200;
        data[68]<=640'd82380930421130208514591602192456812614175954239596008503794331118824453286272729634887977963833354862728303274743662591346725013435792896395326352926655381504;
        data[69]<=640'd123566370976313023803090396825458558807077497481013248406508153003950354552629039991956389071662517411689116159875761730931895855458626834206801549764222517248;
        data[70]<=640'd233406472398421153322362982492754957452371837391271051293079320198475871542681979470129447661822803978026991749405005742697438182615596978466919612056934023168;
        data[71]<=640'd604109837461759778168159595812365051719290138961786243677184080065183411059435054900128032160108089138751203381785997749605204012738286105816714796771764600832;
        data[72]<=640'd604113173047588382820268264222886635157617763925308602241732751467439116477112097925475867510607460983621322460590903413775070191378235877211246055920150511616;
        data[73]<=640'd219675266569980855101260213501077829681437464241079911053085166377405662230442034181704214865795090685004559815270726763607027574337217172861509719847012925440;
        data[74]<=640'd878716019124224372645561183594217863774359502483167172018946154157074302914062729473940378033073734968744706476903378722072150697136375429262006661899186339840;
        data[75]<=640'd1867228367888950619673161100430435175904078019780503412171713751340883795768287523978524475459543415189443776886969609436705478006197723396692008709323596234752;
        data[76]<=640'd2196759186277915900926322250153512660702702110476281457737819979581075412135074665551500504044479750609692663029874974417062491293293797985828882601537181843456;
        data[77]<=640'd3734451812585640249554143841281928450105880192824227291225780984914582739891778147297281175169046805351828243620487176111287055629663337589635468384718758608896;
        data[78]<=640'd1537749138130371623117224962205775229342215845254144378050768554988013656470221484966380435991139240104230028220114544953081115824182065800004499654551648862208;
        data[79]<=640'd8786961745176465666816578199949556679295545572633687054749229839962912457951089140447432383293854575979817958002147119417324729918099622086327887568555216994304;
        data[80]<=640'd10983694272968463208017411114256965826898261436610528015286585374138212436952968448019324691735979715139294022930567373836714236557842930868698303187202758148096;
        data[81]<=640'd16695249082580503456914996506659553199402015551421791061288099602174596231441956973274026555710445567353584232040205477320890597725521914834538813215415933599744;
        data[82]<=640'd1757456916010675963431116897263003454217930426518018828788947740877615651905808648266690413449289711337892111023783134693021225513345144367168930891265539571712;
        data[83]<=640'd36026485773975688680639901527139830520404657341293837627058522077043738777291319753972334416627100670430268025266568532069969983950486661715239027820604686336000;
        data[84]<=640'd3514850144973642398087560138975016262599364512174704303161934339965326802369341883727908966006340731650767137022466249985703598557385084030274527494533533401088;
        data[85]<=640'd29875653048126526639798045376228416843826357165641766152489070646843781580116908296303110864128845455995782506093753715415935597082546797563620705583817795043328;
        data[86]<=640'd63266109313865375643071752977118740822787372271863282812817167781610080094821649312610944792567594094057266609893083522335790396888032046757915281011599004925952;
        data[87]<=640'd3514830033244166381687035798056207455250404591228774179863247277137251617984081560625554648336540389400059265172303182244137258777918140076375065009842498306048;
        data[88]<=640'd175739108367236480040979677000488704101778534884202464425131953194331274773152521036697160974466964807039099562106772512003321904383933565984467335724821647458304;
        data[89]<=640'd56236476063076019515195519781046155012777856211980571718136330521586745378286078675400513575088202484271654880263712893850577998137566993457519853062412287606784;
        data[90]<=640'd140591176749765437445189623810992435795624837489163965356149666762333898095672649144284224911363478561203128175860853594687231528725570829239145539523128057659392;
        data[91]<=640'd224945904252176205082262517795428012740351067217645091963793851838006239238882506518049539620670322340683642412762174233918148560550936107459003180443837531160576;
        data[92]<=640'd337418775931314434710666121368382058581550402986087022736596132649012604514048986252565250960473903116455606423577632442273831910856563706269486414050219291312128;
        data[93]<=640'd84354740910148374269756930822096636120398362898369227892939495922741412985713164212095828237142016513974768879467824348471207636164236838640447402853665597292544;
        data[94]<=640'd112473113019738508644751981776265581042538941086614718041905119717882505495251709234694217409485329140333609937700334099244527421821785361515272197189243978645504;
        data[95]<=640'd309300537899771631082660610980791466418600909514572953475510577119084205660416376460071170766452905968921113612060061181144695409403488757803551940537318830505984;
        data[96]<=640'd56236422431789954785131731391502193504346644638376045558492893439990743552035552631576808305257788610793059377749037847322670386405301057230994913620053708505088;
        data[97]<=640'd0;
        data[98]<=640'd0;
        data[99]<=640'd0;
        data[100]<=640'd0;
        data[101]<=640'd0;
        data[102]<=640'd0;
        data[103]<=640'd0;
        data[104]<=640'd0;
        data[105]<=640'd0;
        data[106]<=640'd0;
        data[107]<=640'd0;
        data[108]<=640'd0;
        data[109]<=640'd0;
        data[110]<=640'd0;
        data[111]<=640'd0;
        data[112]<=640'd0;
        data[113]<=640'd0;
        data[114]<=640'd0;
        data[115]<=640'd0;
        data[116]<=640'd0;
        data[117]<=640'd0;
        data[118]<=640'd0;
        data[119]<=640'd0;
        data[120]<=640'd0;
        data[121]<=640'd0;
        data[122]<=640'd0;
        data[123]<=640'd0;
        data[124]<=640'd0;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd24084754561361768648102764881807084833480156810453237320207177473645930965106688;
        data[156]<=640'd59285549689505892056868344324448208820874232148807968788202283012051522375647232;
        data[157]<=640'd70608395103938906748405107852975316393858956036050582890626880237652602651358048951934797737936631459539297024459407360;
        data[158]<=640'd1067993517960455871195206506167264853458172803453249877212770887222672897722282443732794302529536;
        data[159]<=640'd1432108387429638473108440397114039512156502156033335282210436980904339081275380817489034594535054759240168097957780675895876963965085456942287741255680;
        data[160]<=640'd1634297613668868485164156015396216578334004517111613362205129064985160865023598932487272848798129216410472244711290238003745525127225051113767361839104;
        data[161]<=640'd1432108394384217457882226801255574326011139464744983649041783449188805675173431695226038861926105717710692194195001296951384522668838884790609488379904;
        data[162]<=640'd1432108391049830273401644278722737849120364334060297247134938174134513807501900800215425895994497321779674193266119508278048795711930628599338634313728;
        data[163]<=640'd1432108391049830273401644278735649098510798877008576842994953233506200279217848201550508752554026776391740998501303430948513796217162926072429574881280;
        data[164]<=640'd1432108391526171299756013210551876448029150614539138435787030598275081770131852063681093028035848772279035276784484252021983740776745069051870915330048;
        data[165]<=640'd1432108391430903094485139424276427473980435159081327369931112343416947798816495883946762667839777955560060319458886669030369564042715836043895660085248;
        data[166]<=640'd1432108391145098478672518065078236569389773955797441806254956279136580565305377704354828703225921280575948257942322540404950830814731467307273244639232;
        data[167]<=640'd1432108391049830273401644278885434731737677583139590510899697009561482395899614769493789849643746645578004719839213789355280175744699826568721206345728;
        data[168]<=640'd1432108391240366683943391851601619368030742766333927284091709935377258825841755387755023006139996733793087972122933635263791174054830127011530100703232;
        data[169]<=640'd1432108391240366683943391851932787872881544914369532746030153642378346110315479267891213889398277586815048074848824201678868331002210464713621700083712;
        data[170]<=640'd1432108391240366683943391851439793765575186021972537001975082814418431365900148917796436548155402928625066224028133069778591550624334934584063128764416;
        data[171]<=640'd1432108391240366683943391852097696301894721300657310169440440291010802036052354946265695403268860819323901807682606887736049493626825319704900285759488;
        data[172]<=640'd1432108391240366683943391851436325104722463131847189983357910680153990639517166386655697802812652825225351447018382036542098500500671860454687275745280;
        data[173]<=640'd1432108391240366683943391852758439573882462609540164844889184258255521395328665233478876428054350936568592542451206802170221647341217223133501964943360;
        data[174]<=640'd1432108391240366683943391852758454694402165513535183429747091589205869860762080608186200982928488693054363076974248251870455480179949672581674121035776;
        data[175]<=640'd1432108391240366683943391851436347810133124628554912045016995682792950372117323359224234050582462315933974616390479971711216107968677422227345995988992;
        data[176]<=640'd1432108391240366683943391851436398293952276754886694679738749233495776634893562143924461255720267917347978930242223379402132907988712518980241656381440;
        data[177]<=640'd1432108391240366683943391852758449650944940247175441577215031711861624836036121848420102488350309449414175145035366400014318496270684891491090137350144;
        data[178]<=640'd1432108391240366683943391852097534958051516186622932203928043192673568193247427188323179442600676475226127943314644601783706513087399220109464341315584;
        data[179]<=640'd1432108391240366683943391851932916469218065658024399015447463948022914892991142494164425735624336524730464001216137266799473331018338780953464333664256;
        data[180]<=640'd1432108391240366683943391851542512683980294282207596853941880865913209292374330624151226263653084747640685832721066597117359182906917748229587519668224;
        data[181]<=640'd1432108391240366683943391851602872656675393251684714943904496310492013522598519222722702951934295630385870967567779878798513803820407135863865962659840;
        data[182]<=640'd1432108391240366683943391851467304577476394740390682301184707769031484908245125617811059271175132344711277951347270769406224545795318454304192096894976;
        data[183]<=640'd1432108391240366683943391851436317539537270486124242286683616283446132021635665278696519544222751078836949278101551891706255513177061869120807258554368;
        data[184]<=640'd1432108391049830273401644278720155599242277425470641325827208866944244833533092231581146358403408170107056582211069222276026431019298813863888485875712;
        data[185]<=640'd1432108391145098478672518065078236569389773955797441806254956279136489502701054623304629250605004095551821760436168061530485590687033354070162791202816;
        data[186]<=640'd1432108391430903094485139424152479479832263546777843247541066662367902466614407770004358331660552339384398933352360265046554038560303752771291930689536;
        data[187]<=640'd1432108391526171299756013210510560449979760077104643727987848138723016573772462518240338453399013185499578619903403200659780537093026911160143901097984;
        data[188]<=640'd1432108391049830273401644278720155599242277425470641325910385119929934569407605405930278087475461727557224091197044109104064528251235378250768967532544;
        data[189]<=640'd1432108391049830273401644278720155599242277425470641325860322923775538239351472084691929209789460840314490041901410321420731253428251615359605793619968;
        data[190]<=640'd1432108395908508742216207382982285076764600472137465827655363918997263672051292261884593880915529765509542663695181323129311614392245719303451800764416;
        data[191]<=640'd1636695293373300149939604562666811889736206156746679067232740723557148242244809719794113566873585091269302936828770594755214855647371245708762662567936;
        data[192]<=640'd1636695300423147339984264753164803680650949400929914618905344030551094012883161424892461219733163082806729873652110221921477370731085546254030396719104;
        data[193]<=640'd0;
        data[194]<=640'd0;
        data[195]<=640'd0;
        data[196]<=640'd0;
        data[197]<=640'd0;
        data[198]<=640'd0;
        data[199]<=640'd0;
        data[200]<=640'd0;
        data[201]<=640'd0;
        data[202]<=640'd0;
        data[203]<=640'd0;
        data[204]<=640'd0;
        data[205]<=640'd0;
        data[206]<=640'd0;
        data[207]<=640'd0;
        data[208]<=640'd0;
        data[209]<=640'd0;
        data[210]<=640'd0;
        data[211]<=640'd0;
        data[212]<=640'd0;
        data[213]<=640'd0;
        data[214]<=640'd0;
        data[215]<=640'd0;
        data[216]<=640'd0;
        data[217]<=640'd0;
        data[218]<=640'd0;
        data[219]<=640'd0;
        data[220]<=640'd0;
        data[221]<=640'd0;
        data[222]<=640'd0;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[232]<=640'd770397590192283102817140170538835522329259505150411822303279697242529695245195046002799685574473983146643961599703939665628113080606969752731856666624;
        data[233]<=640'd660112465075810253572230905435385139709417538453094234284389724097390386695711411314593885078474562665473932413317528372647900824072787578972037709824;
        data[234]<=640'd716054195715451547242569712078821989794218681978577542941493380638397682223863664322544223568358465496659348510484073966487713886108951164052813381632;
        data[235]<=640'd716054195763085649878006605265932005736988536484652530568006869144285754519957364185939680360653246015039186276291848311476404846398272228800539394048;
        data[236]<=640'd613760739218697113804657534100821921254332924415468595840795184319585048987268738773011831268338462681830428781582556003620317710710313293594790723584;
        data[237]<=640'd716054195572549239336259032596121955099334801158207852061356801448792723509459789259098704445632947652950208856478036322084310112695811336268335284224;
        data[238]<=640'd716054195715451547242569712158871736014912848257911037340368936190781307546401473706522142986264773530752840604582822950986245390901313328363564171264;
        data[239]<=640'd613760739123428908533783747723284561819669846476611648565781078939270133949827327412482222507784611344649550557121527904178720485958666292289809154048;
        data[240]<=640'd717652518874151265864066222402269279027787839846796175861619257523818687142082218814817992679711572310004459761804083586737166733379098454488554405888;
        data[241]<=640'd717652518874151265864066222381610632332615704134305074641825222183666954728432874421828783111629005463041302381036565731968423454677141348080196517888;
        data[242]<=640'd717652518874151265864066222433256575542502603155916248852776122527065707065293418314348292950721787322273339470492072799817557309478448322165157658624;
        data[243]<=640'd717652518874151265864066222381611262764714851032969703153489812878113119591359665287229035812233413687691056484277674090381605018292200832336385802240;
        data[244]<=640'd717652518874151265864066222422927891246204535366129038416941852957986868373829670928928751727755942778123671315338700284483335127892308009649321279488;
        data[245]<=640'd717652518874151265864066222464243889305289847408319664706551807231782615080806708559487265778625417614943554355564108103210552528348846075417647382528;
        data[246]<=640'd717652518874151265864066222422941760753155997363957340645349445284091451629662381206239642585659882684510732393112810272150190683876353548242328223744;
        data[247]<=640'd717652518874151265864066222464262812119968119874359281204074661850797047518956100846188507001715740008955873382393081498081187779401915774669946880000;
        data[248]<=640'd717652518874151265864066222424419493636110543674992046593395335460949492590608146411639578177457561994558275334553558205843422834747255462656196214784;
        data[249]<=640'd717652518874151265864066222635639503498655084237817294316810812535102180971864697945624697763048565361384137290870518038527754274647884562071155638272;
        data[250]<=640'd717652518874151265864066222404850940396143799638307386426094989071733526486589153511271329430645730213427859000577672767480467749415025584543981633536;
        data[251]<=640'd717652518874151265864066222960034605024083301609186681386654642257410547349926520011929742823092108272697347875369729277014107534145586338041394364416;
        data[252]<=640'd717652518874151265864066222381610671811616575624536626906963505192944409669247814058411920152646564110017106347736831105814939583791750588168174305280;
        data[253]<=640'd717652518874151265864066222381610750538709446680531595425660786388142555758700960183774004641841009710024683102583580712716851135856975197608228159488;
        data[254]<=640'd717652518874151265864066222546874624761086670770212858365523676856183064079662707158119253235780059224649630232176024489037295469165907686078732566528;
        data[255]<=640'd717652518874151265864066222381610750615854520402718549706966991657617018741970816461631098917102044983181923321716996129796342907773975464120745459712;
        data[256]<=640'd615359062091592216613532686273089398809781513253488720619549955218643520191551141955034632786888413165207026731655975418862765051326585983191669014528;
        data[257]<=640'd716054195715451547242569713067823772213345384942636067823464637304320113742015970473715136309880874393107405608024440974814555383516938193572275945472;
        data[258]<=640'd716054195572549239336259032869646426698036064099729672523823473981338174497956614008596886782128718219689104807718113148033925018302225314633891184640;
        data[259]<=640'd613760739218697113804657534050377345521502898846628600636780254417950656343317943091826616036579940120191214515466948119651692478179729438173118332928;
        data[260]<=640'd716054195763085649878006606577392162570678021919213997529348213845994544955425281045347321330072263140128408022846312743591821606798464981227737710592;
        data[261]<=640'd613760739218697113804657535372489361905711875515149648154049558929288904442922753673565904696322360166717555886654962126530863102552070968934947356672;
        data[262]<=640'd723246708519546522626682618670205396500675612725442615919424513077918360251981926363039977843433436239411934400499687063337328814172885954387196772352;
        data[263]<=640'd699271665029450193210545745979964961631808973825901891781574733255418805392616575960024611918592011130701290564316571091104395585953990657037628866560;
        data[264]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[265]<=640'd0;
        data[266]<=640'd0;
        data[267]<=640'd0;
        data[268]<=640'd0;
        data[269]<=640'd0;
        data[270]<=640'd0;
        data[271]<=640'd0;
        data[272]<=640'd0;
        data[273]<=640'd0;
        data[274]<=640'd0;
        data[275]<=640'd0;
        data[276]<=640'd0;
        data[277]<=640'd0;
        data[278]<=640'd0;
        data[279]<=640'd0;
        data[280]<=640'd0;
        data[281]<=640'd0;
        data[282]<=640'd0;
        data[283]<=640'd0;
        data[284]<=640'd0;
        data[285]<=640'd0;
        data[286]<=640'd0;
        data[287]<=640'd0;
        data[288]<=640'd0;
        data[289]<=640'd0;
        data[290]<=640'd0;
        data[291]<=640'd0;
        data[292]<=640'd0;
        data[293]<=640'd0;
        data[294]<=640'd0;
        data[295]<=640'd0;
        data[296]<=640'd0;
        data[297]<=640'd0;
        data[298]<=640'd0;
        data[299]<=640'd0;
        data[300]<=640'd0;
        data[301]<=640'd0;
        data[302]<=640'd0;
        data[303]<=640'd0;
        data[304]<=640'd0;
        data[305]<=640'd0;
        data[306]<=640'd0;
        data[307]<=640'd0;
        data[308]<=640'd0;
        data[309]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[310]<=640'd204586912945874764240387462872684461939791862714291309128701634107400620581789783294404734467263753122353208725382371822087818297065713413500142878720;
        data[311]<=640'd613760738932892497992036174976134355966872118469674407814113055119417345132374102654813496008001772766214044241327380698239975365301387545166208827392;
        data[312]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[313]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[314]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[315]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[316]<=640'd716054195810719752513443498444785882909390677394503417248096665387912638568274816216319923546195994976306584519426322962481530122975535690971336409088;
        data[317]<=640'd716054195810719752513443498455645706249216138177074917164337847650413495987043420765153160381100583828079559719301877370587891032232095271147739807744;
        data[318]<=640'd716054195810719752513443498453879235507419380885030023238568209156304161116069913860135702491201439629619796773170952985848890494223452525086304632832;
        data[319]<=640'd716054195810719752513443498510497081467286048813882673100702951077881354187596314511773640630805727762155028983613816104686710516071829618063174533120;
        data[320]<=640'd716054195810719752513443498460143208844760463077529821080196447904555248326788557900137008901452003884198374928910000939410338251252270873223882604544;
        data[321]<=640'd716054195810719752513443498527281705674757012943335194389606949037152868359891240043216593653491645666403208387701926563269058460469809487764755841024;
        data[322]<=640'd716054195810719752513443498496294707137714183259419876007859178091465048512722663379328334759999833805043974433678217155421262723832670948113755668480;
        data[323]<=640'd716054195810719752513443498434320710063628340411699960038642707334417784651430246326352683510526311075218355571800711260941025649074145058756830953472;
        data[324]<=640'd716054195810719752513443498558268704211799916019206224453643091529109337873841922197184505931979417130605302723257670802630712437700647551437725761536;
        data[325]<=640'd716054195810719752513443498516952706162409451976667229383883273086102694855356451481973609612325014781178703990715379981662365375319896323895735615488;
        data[326]<=640'd716054195810719752513443498682277239580970957473452572422737403252585741964642850032475924422476581956582228806857619203036121907734186946087295647744;
        data[327]<=640'd716054195810719752513443498434744419768282745649118736482402421171162494035848669017568008616338471606971782403100048999294815896607485478661200543744;
        data[328]<=640'd716054195810719752513443498520180528360672884949629464011945630600911020862581413767102341587340635449994773464501007948977127920534674423705717702656;
        data[329]<=640'd716054195810719752513443498831341654677359009438988984845728250751230595399040954295930091273722750741024138770869931854569551962827351533791681183744;
        data[330]<=640'd716054195810719752513443498568597705571117911889023924498425831553495752160349493373008716848145533793862362408284626593044442791861272334534858244096;
        data[331]<=640'd716054195810719752513443498682216713136025199340772216790481268029865924641872019504655454319950658852344070947469645236329109806197610742822886965248;
        data[332]<=640'd716054195810719752513443498599584702262693814274499031200694035285404404923758357194094993893866283716026817139533485184985118062016148369030003032064;
        data[333]<=640'd716054195810719752513443499425904673101307019081430866693741199808277343705677208242846533457381245478574006576665460295014574276902122092042165157888;
        data[334]<=640'd716054195810719752513443498764848716623583836033777364462676998056899305882677914285810678489932238168967027307797086834675354174885748935025999478784;
        data[335]<=640'd716054195810719752513443498434320870134880584746327199572416971885421633060395155659807563156893148679265402023997279477454964846962619427443290669056;
        data[336]<=640'd306880369680799710855484106793991606815030501076763680436902581899057953303635566656631382197081352848945907415008763377082799821359458943348521304064;
        data[337]<=640'd613760739028160703262909963319642702360957109387239577243211078328533778236478806517612820973929906066910998918547738826236082253914121697165618184192;
        data[338]<=640'd102293456734924946615096645243179359725950936144764159100633581358749766618167605902753369491196967141042489028467367422896442277928099059984043606016;
        data[339]<=640'd511467282579040372460434677197512054772106434783894694398887777683205499804609093785730877190317093938089118226762781376498788721480370995835831320576;
        data[340]<=640'd463517230514644945403403635537161829322059742570818762195456572280078361975720658521061960032081583455871415023902052716166488001030753226626093285376;
        data[341]<=640'd40757545357465589008840466789133681118391266897917571308776845053923947707004850323457321705794696241597790325850590410003784231118969220988854599680;
        data[342]<=640'd305282044807272297358259442042921005743881775842346186293723637886603009040190077170326453720151994149802200483234037215585421063200410814574330118144;
        data[343]<=640'd0;
        data[344]<=640'd0;
        data[345]<=640'd0;
        data[346]<=640'd0;
        data[347]<=640'd0;
        data[348]<=640'd0;
        data[349]<=640'd0;
        data[350]<=640'd0;
        data[351]<=640'd0;
        data[352]<=640'd0;
        data[353]<=640'd0;
        data[354]<=640'd0;
        data[355]<=640'd0;
        data[356]<=640'd0;
        data[357]<=640'd0;
        data[358]<=640'd0;
        data[359]<=640'd0;
        data[360]<=640'd0;
        data[361]<=640'd0;
        data[362]<=640'd0;
        data[363]<=640'd0;
        data[364]<=640'd0;
        data[365]<=640'd0;
        data[366]<=640'd0;
        data[367]<=640'd0;
        data[368]<=640'd0;
        data[369]<=640'd0;
        data[370]<=640'd0;
        data[371]<=640'd0;
        data[372]<=640'd0;
        data[373]<=640'd0;
        data[374]<=640'd0;
        data[375]<=640'd0;
        data[376]<=640'd0;
        data[377]<=640'd0;
        data[378]<=640'd0;
        data[379]<=640'd0;
        data[380]<=640'd0;
        data[381]<=640'd0;
        data[382]<=640'd0;
        data[383]<=640'd0;
        data[384]<=640'd0;
        data[385]<=640'd0;
        data[386]<=640'd0;
        data[387]<=640'd0;
        data[388]<=640'd0;
        data[389]<=640'd0;
        data[390]<=640'd0;
        data[391]<=640'd0;
        data[392]<=640'd0;
        data[393]<=640'd0;
        data[394]<=640'd0;
        data[395]<=640'd0;
        data[396]<=640'd0;
        data[397]<=640'd0;
        data[398]<=640'd0;
        data[399]<=640'd0;
        data[400]<=640'd0;
        data[401]<=640'd0;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd22835963083295687686091155745995325592756551680;
        data[406]<=640'd22836137307867241909738992724944393428252229632;
        data[407]<=640'd45671926166592015614959756397608870041507332096;
        data[408]<=640'd11419593118938734974605247813455870800613605376;
        data[409]<=640'd92102251995524685136327182220460836482002714624;
        data[410]<=640'd713798081558695355229084985473875756514803712;
        data[411]<=640'd79973270849186984475343595013176781527727472640;
        data[412]<=640'd758237586915271256831821758006986185344286720;
        data[413]<=640'd188396706326222447116603965185342682481500880896;
        data[414]<=640'd10634488215193846815532761681284300800;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
    else if (choise == 2) begin
        data[0]<=640'd0;
        data[1]<=640'd0;
        data[2]<=640'd0;
        data[3]<=640'd0;
        data[4]<=640'd0;
        data[5]<=640'd0;
        data[6]<=640'd0;
        data[7]<=640'd0;
        data[8]<=640'd0;
        data[9]<=640'd0;
        data[10]<=640'd0;
        data[11]<=640'd0;
        data[12]<=640'd0;
        data[13]<=640'd0;
        data[14]<=640'd0;
        data[15]<=640'd0;
        data[16]<=640'd0;
        data[17]<=640'd0;
        data[18]<=640'd0;
        data[19]<=640'd0;
        data[20]<=640'd0;
        data[21]<=640'd0;
        data[22]<=640'd0;
        data[23]<=640'd0;
        data[24]<=640'd0;
        data[25]<=640'd0;
        data[26]<=640'd0;
        data[27]<=640'd0;
        data[28]<=640'd0;
        data[29]<=640'd0;
        data[30]<=640'd0;
        data[31]<=640'd0;
        data[32]<=640'd0;
        data[33]<=640'd0;
        data[34]<=640'd0;
        data[35]<=640'd0;
        data[36]<=640'd0;
        data[37]<=640'd0;
        data[38]<=640'd0;
        data[39]<=640'd0;
        data[40]<=640'd0;
        data[41]<=640'd0;
        data[42]<=640'd0;
        data[43]<=640'd0;
        data[44]<=640'd0;
        data[45]<=640'd0;
        data[46]<=640'd0;
        data[47]<=640'd0;
        data[48]<=640'd0;
        data[49]<=640'd0;
        data[50]<=640'd0;
        data[51]<=640'd0;
        data[52]<=640'd2293498615990071511610820895302086940796564989168281123737588839386922876088484808070018553110125686554624;
        data[53]<=640'd1675976290930685468645128323187019804819274807935478584355997288644324119240316295174021690532034581474959799140168891292198173855926923755850975816974336;
        data[54]<=640'd18016743004716045104939568706166646234830913194566828459917631673408091544086843037861291450401948673299982734405370585939836303642089739931020670818844672;
        data[55]<=640'd42318397475031701438889607385923245877036691254239602651234569147285240898305566161081713485969712312403657740930550414975923248456038202051341749537734656;
        data[56]<=640'd57402183344188992557480846249111134803883445987125003633414363911957637828907724366345008656219299889741061112297913938112867822288523357300753250694201344;
        data[57]<=640'd42318407564523126557606423241263499347310989384703844829702022658899048385630712785314992999361375193054543958740802212534772278779117267377539787870175232;
        data[58]<=640'd395530360905215115021967377632711409942006648779440471063266579816800946473045629048871445053568278627989595852987097636404105016876635012054155033330057216;
        data[59]<=640'd875906954421202713545704567352562934563026676853642611817926797221644961654863567688143481820911674474299584801504605189711145700733634866251699676946366464;
        data[60]<=640'd1074300936946526427302439310125071297515937130994533697009700542908227236054607196059323136753822689742996809766773833370569381539617161493151705275232681984;
        data[61]<=640'd2723730804743768237183904232934132161590198535360849222019756894908502785821633132584250944977698014866267721515232107944067370552804837045185415225540608;
        data[62]<=640'd5363542191748007292225498426358644037797628068518507929096833266769054255422522206636867302888064784899710315832520857566929660082277303334339182503433076736;
        data[63]<=640'd3142916103311877827994774634041287214440824010129971401946070220615944633674407965106679014548230495399058990158957803742790727468293186791713320095186944;
        data[64]<=640'd11157391883955290085745718645693946645242694238428966059551126335989982129014637808743606319664413813119272322494123819208654259517587023408725019044406624256;
        data[65]<=640'd46340318392186936109177457491811105143390564853932790665686560000254254661569666650423555483369856326553091574677262891816660630792352920929528114164621377536;
        data[66]<=640'd2096606884159293981315126535532627615023078102265478175759719763157201612263761929777286175608312879866159756539412255745900722075555602617940478057775104;
        data[67]<=640'd6866055053295803659884082352104202948505894945454718108404934879957895628581040891606397478280400890069828080887171596984391567232311544567374210143564595200;
        data[68]<=640'd82380930421130208514591602192456812614175954239596008503794331118824453286272729634887977963833354862728303274743662591346725013435792896395326352926655381504;
        data[69]<=640'd123566370976313023803090396825458558807077497481013248406508153003950354552629039991956389071662517411689116159875761730931895855458626834206801549764222517248;
        data[70]<=640'd233406472398421153322362982492754957452371837391271051293079320198475871542681979470129447661822803978026991749405005742697438182615596978466919612056934023168;
        data[71]<=640'd604109837461759778168159595812365051719290138961786243677184080065183411059435054900128032160108089138751203381785997749605204012738286105816714796771764600832;
        data[72]<=640'd604113173047588382820268264222886635157617763925308602241732751467439116477112097925475867510607460983621322460590903413775070191378235877211246055920150511616;
        data[73]<=640'd219675266569980855101260213501077829681437464241079911053085166377405662230442034181704214865795090685004559815270726763607027574337217172861509719847012925440;
        data[74]<=640'd878716019124224372645561183594217863774359502483167172018946154157074302914062729473940378033073734968744706476903378722072150697136375429262006661899186339840;
        data[75]<=640'd1867228367888950619673161100430435175904078019780503412171713751340883795768287523978524475459543415189443776886969609436705478006197723396692008709323596234752;
        data[76]<=640'd2196759186277915900926322250153512660702702110476281457737819979581075412135074665551500504044479750609692663029874974417062491293293797985828882601537181843456;
        data[77]<=640'd3734451812585640249554143841281928450105880192824227291225780984914582739891778147297281175169046805351828243620487176111287055629663337589635468384718758608896;
        data[78]<=640'd1537749138130371623117224962205775229342215845254144378050768554988013656470221484966380435991139240104230028220114544953081115824182065800004499654551648862208;
        data[79]<=640'd8786961745176465666816578199949556679295545572633687054749229839962912457951089140447432383293854575979817958002147119417324729918099622086327887568555216994304;
        data[80]<=640'd10983694272968463208017411114256965826898261436610528015286585374138212436952968448019324691735979715139294022930567373836714236557842930868698303187202758148096;
        data[81]<=640'd16695249082580503456914996506659553199402015551421791061288099602174596231441956973274026555710445567353584232040205477320890597725521914834538813215415933599744;
        data[82]<=640'd1757456916010675963431116897263003454217930426518018828788947740877615651905808648266690413449289711337892111023783134693021225513345144367168930891265539571712;
        data[83]<=640'd36026485773975688680639901527139830520404657341293837627058522077043738777291319753972334416627100670430268025266568532069969983950486661715239027820604686336000;
        data[84]<=640'd3514850144973642398087560138975016262599364512174704303161934339965326802369341883727908966006340731650767137022466249985703598557385084030274527494533533401088;
        data[85]<=640'd29875653048126526639798045376228416843826357165641766152489070646843781580116908296303110864128845455995782506093753715415935597082546797563620705583817795043328;
        data[86]<=640'd63266109313865375643071752977118740822787372271863282812817167781610080094821649312610944792567594094057266609893083522335790396888032046757915281011599004925952;
        data[87]<=640'd3514830033244166381687035798056207455250404591228774179863247277137251617984081560625554648336540389400059265172303182244137258777918140076375065009842498306048;
        data[88]<=640'd175739108367236480040979677000488704101778534884202464425131953194331274773152521036697160974466964807039099562106772512003321904383933565984467335724821647458304;
        data[89]<=640'd56236476063076019515195519781046155012777856211980571718136330521586745378286078675400513575088202484271654880263712893850577998137566993457519853062412287606784;
        data[90]<=640'd140591176749765437445189623810992435795624837489163965356149666762333898095672649144284224911363478561203128175860853594687231528725570829239145539523128057659392;
        data[91]<=640'd224945904252176205082262517795428012740351067217645091963793851838006239238882506518049539620670322340683642412762174233918148560550936107459003180443837531160576;
        data[92]<=640'd337418775931314434710666121368382058581550402986087022736596132649012604514048986252565250960473903116455606423577632442273831910856563706269486414050219291312128;
        data[93]<=640'd84354740910148374269756930822096636120398362898369227892939495922741412985713164212095828237142016513974768879467824348471207636164236838640447402853665597292544;
        data[94]<=640'd112473113019738508644751981776265581042538941086614718041905119717882505495251709234694217409485329140333609937700334099244527421821785361515272197189243978645504;
        data[95]<=640'd309300537899771631082660610980791466418600909514572953475510577119084205660416376460071170766452905968921113612060061181144695409403488757803551940537318830505984;
        data[96]<=640'd56236422431789954785131731391502193504346644638376045558492893439990743552035552631576808305257788610793059377749037847322670386405301057230994913620053708505088;
        data[97]<=640'd0;
        data[98]<=640'd0;
        data[99]<=640'd0;
        data[100]<=640'd0;
        data[101]<=640'd0;
        data[102]<=640'd0;
        data[103]<=640'd0;
        data[104]<=640'd0;
        data[105]<=640'd0;
        data[106]<=640'd0;
        data[107]<=640'd0;
        data[108]<=640'd0;
        data[109]<=640'd0;
        data[110]<=640'd0;
        data[111]<=640'd0;
        data[112]<=640'd0;
        data[113]<=640'd0;
        data[114]<=640'd0;
        data[115]<=640'd0;
        data[116]<=640'd0;
        data[117]<=640'd0;
        data[118]<=640'd0;
        data[119]<=640'd0;
        data[120]<=640'd0;
        data[121]<=640'd0;
        data[122]<=640'd0;
        data[123]<=640'd0;
        data[124]<=640'd0;
        data[125]<=640'd0;
        data[126]<=640'd0;
        data[127]<=640'd0;
        data[128]<=640'd0;
        data[129]<=640'd0;
        data[130]<=640'd0;
        data[131]<=640'd0;
        data[132]<=640'd0;
        data[133]<=640'd0;
        data[134]<=640'd0;
        data[135]<=640'd0;
        data[136]<=640'd0;
        data[137]<=640'd0;
        data[138]<=640'd0;
        data[139]<=640'd0;
        data[140]<=640'd0;
        data[141]<=640'd0;
        data[142]<=640'd0;
        data[143]<=640'd0;
        data[144]<=640'd0;
        data[145]<=640'd0;
        data[146]<=640'd0;
        data[147]<=640'd0;
        data[148]<=640'd0;
        data[149]<=640'd0;
        data[150]<=640'd0;
        data[151]<=640'd0;
        data[152]<=640'd0;
        data[153]<=640'd0;
        data[154]<=640'd0;
        data[155]<=640'd24084754561361768648102764881807084833480156810453237320207177473645930965106688;
        data[156]<=640'd59285549689505892056868344324448208820874232148807968788202283012051522375647232;
        data[157]<=640'd70608395103938906748405107852975316393858956036050582890626880237652602651358048951934797737936631459539297024459407360;
        data[158]<=640'd1067993517960455871195206506167264853458172803453249877212770887222672897722282443732794302529536;
        data[159]<=640'd1432108387429638473108440397114039512156502156033335282210436980904339081275380817489034594535054759240168097957780675895876963965085456942287741255680;
        data[160]<=640'd1482454398797580680866649042122612815302120059747903671214493780776674881095288810163559527736042930252138552617983715178619500728112098446507706941440;
        data[161]<=640'd1432108395908508742216207382984869848371083949973791335889913893944253409365507739571627543625473932097162883237885540663008850254506841665261971439616;
        data[162]<=640'd1432108391049830273401644278722737849120364334060297247134938174134513807501900800215425895994497321779674193266119508278048795711930628599338634313728;
        data[163]<=640'd1432108391049830273401644278735649098510798877008576842994953233506200279217848201550508752554026776391740998501303430948513796217162926072429574881280;
        data[164]<=640'd1432108391526171299756013210551876448029150614539138435787030598275081770131852063681093028035848772279035276784484252021983740776745069051870915330048;
        data[165]<=640'd1432108391430903094485139424276427473980435159081327369931112343416947798816495883946762667839777955560060319458886669030369564042715836043895660085248;
        data[166]<=640'd1432108391145098478672518065078236569389773955797441806254956279136580565305377704354828703225921280575948257942322540404950830814731467307273244639232;
        data[167]<=640'd1432108391049830273401644278885434731737677583139590510899697009561482395899614769493789849643746645578004719839213789355280175744699826568721206345728;
        data[168]<=640'd1432108391240366683943391851601619368030742766333927284091709935377258825841755387755023006139996733793087972122933635263791174054830127011530100703232;
        data[169]<=640'd1432108391240366683943391851932787872881544914369532746030153642378346110315479267891213889398277586815048074848824201678868331002210464713621700083712;
        data[170]<=640'd1432108391240366683943391851439793765575186021972537001975082814418431365900148917796436548155402928625066224028133069778591550624334934584063128764416;
        data[171]<=640'd1432108391240366683943391852097696301894721300657310169440440291010802036052354946265695403268860819323901807682606887736049493626825319704900285759488;
        data[172]<=640'd1432108391240366683943391851436325104722463131847189983357910680153990639517166386655697802812652825225351447018382036542098500500671860454687275745280;
        data[173]<=640'd1432108391240366683943391852758439573882462609540164844889184258255521395328665233478876428054350936568592542451206802170221647341217223133501964943360;
        data[174]<=640'd1432108391240366683943391852758454694402165513535183429747091589205869860762080608186200982928488693054363076974248251870455480179949672581674121035776;
        data[175]<=640'd1432108391240366683943391851436347810133124628554912045016995682792950372117323359224234050582462315933974616390479971711216107968677422227345995988992;
        data[176]<=640'd1432108391240366683943391851436398293952276754886694679738749233495776634893562143924461255720267917347978930242223379402132907988712518980241656381440;
        data[177]<=640'd1432108391240366683943391852758449650944940247175441577215031711861624836036121848420102488350309449414175145035366400014318496270684891491090137350144;
        data[178]<=640'd1432108391240366683943391852097534958051516186622932203928043192673568193247427188323179442600676475226127943314644601783706513087399220109464341315584;
        data[179]<=640'd1432108391240366683943391851932916469218065658024399015447463948022914892991142494164425735624336524730464001216137266799473331018338780953464333664256;
        data[180]<=640'd1432108391240366683943391851542512683980294282207596853941880865913209292374330624151226263653084747640685832721066597117359182906917748229587519668224;
        data[181]<=640'd1432108391240366683943391851602872656675393251684714943904496310492013522598519222722702951934295630385870967567779878798513803820407135863865962659840;
        data[182]<=640'd1432108391240366683943391851467304577476394740390682301184707769031484908245125617811059271175132344711277951347270769406224545795318454304192096894976;
        data[183]<=640'd1432108391240366683943391851436317539537270486124242286683616283446132021635665278696519544222751078836949278101551891706255513177061869120807258554368;
        data[184]<=640'd1432108391049830273401644278720155599242277425470641325827208866944244833533092231581146358403408170107056582211069222276026431019298813863888485875712;
        data[185]<=640'd1432108391145098478672518065078236569389773955797441806254956279136489502701054623304629250605004095551821760436168061530485590687033354070162791202816;
        data[186]<=640'd1432108391430903094485139424152479479832263546777843247541066662367902466614407770004358331660552339384398933352360265046554038560303752771291930689536;
        data[187]<=640'd1432108391526171299756013210510560449979760077104643727987848138723016573772462518240338453399013185499578619903403200659780537093026911160143901097984;
        data[188]<=640'd1432108391049830273401644278720155599242277425470641325910385119929934569407605405930278087475461727557224091197044109104064528251235378250768967532544;
        data[189]<=640'd1432108391049830273401644278720155599242277425470641325860322923775538239351472084691929209789460840314490041901410321420731253428251615359605793619968;
        data[190]<=640'd1432108395908508742216207382982285076764600472137465827655363918997263672051292261884593880915529765509542663695181323129311614392245719303451800764416;
        data[191]<=640'd1636695299470465287275526889583993979175984097661909814625262502578939179013113897176468293671057948815185693000307569601712165990043073207372594806784;
        data[192]<=640'd1636695300423147339984264753164803680650949400929914618905344030551094012883161424892461219733163082806729873652110221921477370731085546254030396719104;
        data[193]<=640'd0;
        data[194]<=640'd0;
        data[195]<=640'd0;
        data[196]<=640'd0;
        data[197]<=640'd0;
        data[198]<=640'd0;
        data[199]<=640'd0;
        data[200]<=640'd0;
        data[201]<=640'd0;
        data[202]<=640'd0;
        data[203]<=640'd0;
        data[204]<=640'd0;
        data[205]<=640'd0;
        data[206]<=640'd0;
        data[207]<=640'd0;
        data[208]<=640'd0;
        data[209]<=640'd0;
        data[210]<=640'd0;
        data[211]<=640'd0;
        data[212]<=640'd0;
        data[213]<=640'd0;
        data[214]<=640'd0;
        data[215]<=640'd0;
        data[216]<=640'd0;
        data[217]<=640'd0;
        data[218]<=640'd0;
        data[219]<=640'd0;
        data[220]<=640'd0;
        data[221]<=640'd0;
        data[222]<=640'd0;
        data[223]<=640'd0;
        data[224]<=640'd0;
        data[225]<=640'd0;
        data[226]<=640'd0;
        data[227]<=640'd0;
        data[228]<=640'd0;
        data[229]<=640'd0;
        data[230]<=640'd0;
        data[231]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[232]<=640'd770397583999849760210344057263572462741985033908380594482749765423523275089886115848845666170790612201606787362986699587154282263830894949456144236544;
        data[233]<=640'd660112465837955895739221196300032900889389781067498077708454946475114253791749433487388225928158669858709276934759650228460064616906766016298279239680;
        data[234]<=640'd716054195715451547242569712078821989794218681978577542941493380638397682223863664322544223568358465496659348510484073966487713886108951164052813381632;
        data[235]<=640'd716054195763085649878006605265932005736988536484652530568006869144285754519957364185939680360653246015039186276291848311476404846398272228800539394048;
        data[236]<=640'd613760739218697113804657534100821921254332924415468595840795184319585048987268738773011831268338462681830428781582556003620317710710313293594790723584;
        data[237]<=640'd716054195572549239336259032596121955099334801158207852061356801448792723509459789259098704445632947652950208856478036322084310112695811336268335284224;
        data[238]<=640'd613760739028160703262909961416847322213149723665464301812999775343346159634745888323221367388659241821478795595236040267995165175633900186115487301632;
        data[239]<=640'd613760739028160703262909961365203591672173316149811168137772926142054650562822574640882929901574097945495132491941262672202200011854418987624028962816;
        data[240]<=640'd716054195810719752513443498454979356758800439428213205417422927204072370348414853582025849549888779512536140716143873088809318055174957849631598313472;
        data[241]<=640'd716054195810719752513443498434320710063628303715722104197628891863920637934765509189036639981806212665572983335376355234040574776473000743223240425472;
        data[242]<=640'd716054195810719752513443498485966653273515202737333278408579792207319390271626053081556149820898994524805020424831862301889708631274307717308201566208;
        data[243]<=640'd716054195810719752513443498434321340495727450614386732709293482558366802797692300054436892682410620890222737438617463592453756340088060227479429709824;
        data[244]<=640'd716054195810719752513443498475637968977217134947546067972745522638240551580162305696136608597933149980655352269678489786555486449688167404792365187072;
        data[245]<=640'd716054195810719752513443498516953967036302446989736694262355476912036298287139343326695122648802624817475235309903897605282703850144705470560691290112;
        data[246]<=640'd716054195810719752513443498475651838484168596945374370201153114964345134835995015973447499455837089887042413347452599774222342005672212943385372131328;
        data[247]<=640'd716054195810719752513443498516972889850980719455776310759878331531050730725288735613396363871892947211487554336732871000153339101197775169812990787584;
        data[248]<=640'd716054195810719752513443498477129571367123143256409076149199005141203175796940781178847435047634769197089956288893347707915574156543114857799240122368;
        data[249]<=640'd716054195810719752513443498688349581229667683819234323872614482215355864178197332712832554633225772563915818245210307540599905596443743957214199545856;
        data[250]<=640'd716054195810719752513443498457561018127156399219724415981898658751987209692921788278479186300822937415959539954917462269552619071210884979687025541120;
        data[251]<=640'd716054195810719752513443499012744682755095901190603710942458311937664230556259154779137599693269315475229028829709518779086258855941445733184438272000;
        data[252]<=640'd716054195810719752513443498434320749542629175205953656462767174873198092875580448825619777022823771312548787302076620607887090905587609983311218212864;
        data[253]<=640'd716054195810719752513443498434320828269722046261948624981464456068396238965033594950981861512018216912556364056923370214789002457652834592751272067072;
        data[254]<=640'd716054195810719752513443498599584702492099270351629887921327346536436747285995341925327110105957266427181311186515813991109446790961767081221776474112;
        data[255]<=640'd716054195810719752513443498434320828346867119984135579262770661337870701948303451228838955787279252185713604276056785631868494229569834859263789367296;
        data[256]<=640'd613760739123428908533783748683880446688290643161706230603361777696112686784888529493841782263276133766893125751176030152911436847226692683000493113344;
        data[257]<=640'd613760739218697113804657535041961298706575321003790293152111782051315932604369890633612945924696369482142196729038188755776516116458019660655759458304;
        data[258]<=640'd716054195572549239336259032869646426698036064099729672523823473981338174497956614008596886782128718219689104807718113148033925018302225314633891184640;
        data[259]<=640'd613760739171063011169220640871336860447754633683228360422776178019342914649815566706026969733474683420614005482876815503663432241127605785840228237312;
        data[260]<=640'd716054195763085649878006606577392162570678021919213997529348213845994544955425281045347321330072263140128408022846312743591821606798464981227737710592;
        data[261]<=640'd716054195715451547242569713398351835412481939453995422825402414182293085580568833513668095081506865077682764765641214345568902369610989501851463843840;
        data[262]<=640'd660112465647419485197473623578706460838222903234585278508432617132023875432081480918528322002656347816366758415139829057946748005826465063021223870464;
        data[263]<=640'd770397583618776939126848911831248582151998912601178672770717154234661341541867104762448495745948558604989115102265638659248200367413905730793023471616;
        data[264]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[265]<=640'd0;
        data[266]<=640'd0;
        data[267]<=640'd0;
        data[268]<=640'd0;
        data[269]<=640'd0;
        data[270]<=640'd0;
        data[271]<=640'd0;
        data[272]<=640'd0;
        data[273]<=640'd0;
        data[274]<=640'd0;
        data[275]<=640'd0;
        data[276]<=640'd0;
        data[277]<=640'd0;
        data[278]<=640'd0;
        data[279]<=640'd0;
        data[280]<=640'd0;
        data[281]<=640'd0;
        data[282]<=640'd0;
        data[283]<=640'd0;
        data[284]<=640'd0;
        data[285]<=640'd0;
        data[286]<=640'd0;
        data[287]<=640'd0;
        data[288]<=640'd0;
        data[289]<=640'd0;
        data[290]<=640'd0;
        data[291]<=640'd0;
        data[292]<=640'd0;
        data[293]<=640'd0;
        data[294]<=640'd0;
        data[295]<=640'd0;
        data[296]<=640'd0;
        data[297]<=640'd0;
        data[298]<=640'd0;
        data[299]<=640'd0;
        data[300]<=640'd0;
        data[301]<=640'd0;
        data[302]<=640'd0;
        data[303]<=640'd0;
        data[304]<=640'd0;
        data[305]<=640'd0;
        data[306]<=640'd0;
        data[307]<=640'd0;
        data[308]<=640'd0;
        data[309]<=640'd818347651926401364867860531027859302980412246347365957156818765625425707407666262335017876778370782588144461999299885136316053899419224610999241801728;
        data[310]<=640'd204586912945874764240387462872684461939791862714291309128701634107400620581789783294404734467263753122353208725382371822087818297065713413500142878720;
        data[311]<=640'd613760738932892497992036174976134355966872118469674407814113055119417345132374102654813496008001772766214044241327380698239975365301387545166208827392;
        data[312]<=640'd613760739313965319075531320408458236556858239776876329526145666308279278680393113741210666432843826362831716502048441626146057261718376763829329592320;
        data[313]<=640'd716054195810719752513443498434320710063628303715722104197498521561283459818039193581312856818028331273796925381034693845184096528777295296745846079488;
        data[314]<=640'd613760739313965319075531320408458236556858239776876329526145666308279278680393113741210666432843826362831716502048441626146057261718376763829329592320;
        data[315]<=640'd613760739313965319075531320408458236556858239776876329526145666308279278680393113741210666432843826362831716502048441626146057261718376763829329592320;
        data[316]<=640'd716054195810719752513443498444785882909390677394503417248096665387912638568274816216319923546195994976306584519426322962481530122975535690971336409088;
        data[317]<=640'd615358330717580352115474814315222422238080564829122425834567840102243219446563420275275897428995966208651929301538854069800459322758017509896310751232;
        data[318]<=640'd717652518874151265864066222401169157776406781303612993682764539476050477909737279092927845621024232427088115818831163483776739172427593129943260725248;
        data[319]<=640'd614484972783308354601367197207582443663893777813673676951305862195928385756748065530829907666586237896733387609573780529165794494026850970117852889088;
        data[320]<=640'd717652518874151265864066222407433131113747863496112791524392778224301565120455923132929152031274796681666693974570211437338186929456411478080838696960;
        data[321]<=640'd717652518874151265864066222474571627943744413361918164833803279356899185153558605276008736783314438463871527433362137061196907138673950092621711933440;
        data[322]<=640'd717652518874151265864066222443584629406701583678002846452055508411211365306390028612120477889822626602512293479338427653349111402036811552970711760896;
        data[323]<=640'd717652518874151265864066222381610632332615740830282930482839037654164101445097611559144826640349103872686674617460921758868874327278285663613787045888;
        data[324]<=640'd717652518874151265864066222505558626480787316437789194897839421848855654667509287429976649061802209928073621768917881300558561115904788156294681853952;
        data[325]<=640'd717652518874151265864066222464242628431396852395250199828079603405849011649023816714765752742147807578647023036375590479590214053524036928752691707904;
        data[326]<=640'd717652518874151265864066222629567161849958357892035542866933733572332058758310215265268067552299374754050547852517829700963970585938327550944251740160;
        data[327]<=640'd717652518874151265864066222382034342037270146067701706926598751490908810829516034250360151746161264404440101448760259497222664574811626083518156636160;
        data[328]<=640'd716853351245270371852832533576643400055388644243690201841522016738993242491110919001143686354779174302846176815794138351443741916964917227524263510016;
        data[329]<=640'd717652518874151265864066222778631576946346409857571955289924581070976912192708319528722234403545543538492457816530142352497400641031492138648637276160;
        data[330]<=640'd717652518874151265864066222515887627840105312307606894942622161873242068954016858605800859977968326591330681453944837090972291470065412939391814336512;
        data[331]<=640'd615359062377396832426154044603644161898242535820509412563324743096608060297893304897345407064588946738847181114143603515218919217342832814763326570496;
        data[332]<=640'd717652518874151265864066222546874624531681214693082001644890365605150721717425722426887137023689076513495136185193695682912966740220288973886959124480;
        data[333]<=640'd716853363439600646524677188316731723675578660205953099308361143989941438870815068241597331819765499423190922271032540390475808958676019893080575442944;
        data[334]<=640'd613760739313965319075531320738986243116813772094931589791324142803895124745031834445708488104747733258001818428810834615637314907826830402109482991616;
        data[335]<=640'd716054195810719752513443498434320870134880584746327199572416971885421633060395155659807563156893148679265402023997279477454964846962619427443290669056;
        data[336]<=640'd306880369680799710855484106793991606815030501076763680436902581899057953303635566656631382197081352848945907415008763377082799821359458943348521304064;
        data[337]<=640'd613760739028160703262909963319642702360957109387239577243211078328533778236478806517612820973929906066910998918547738826236082253914121697165618184192;
        data[338]<=640'd102293456734924946615096645243179359725950936144764159100633581358749766618167605902753369491196967141042489028467367422896442277928099059984043606016;
        data[339]<=640'd511467282579040372460434677197512054772106434783894694398887777683205499804609093785730877190317093938089118226762781376498788721480370995835831320576;
        data[340]<=640'd463517230514644945403403635537161829322059742570818762195456572280078361975720658521061960032081583455871415023902052716166488001030753226626093285376;
        data[341]<=640'd40757545357465589008840466789133681118391266897917571308776845053923947707004850323457321705794696241597790325850590410003784231118969220988854599680;
        data[342]<=640'd305282044807272297358259442042921005743881775842346186293723637886603009040190077170326453720151994149802200483234037215585421063200410814574330118144;
        data[343]<=640'd0;
        data[344]<=640'd0;
        data[345]<=640'd0;
        data[346]<=640'd0;
        data[347]<=640'd0;
        data[348]<=640'd0;
        data[349]<=640'd0;
        data[350]<=640'd0;
        data[351]<=640'd0;
        data[352]<=640'd0;
        data[353]<=640'd0;
        data[354]<=640'd0;
        data[355]<=640'd0;
        data[356]<=640'd0;
        data[357]<=640'd0;
        data[358]<=640'd0;
        data[359]<=640'd0;
        data[360]<=640'd0;
        data[361]<=640'd0;
        data[362]<=640'd0;
        data[363]<=640'd0;
        data[364]<=640'd0;
        data[365]<=640'd0;
        data[366]<=640'd0;
        data[367]<=640'd0;
        data[368]<=640'd0;
        data[369]<=640'd0;
        data[370]<=640'd0;
        data[371]<=640'd0;
        data[372]<=640'd0;
        data[373]<=640'd0;
        data[374]<=640'd0;
        data[375]<=640'd0;
        data[376]<=640'd0;
        data[377]<=640'd0;
        data[378]<=640'd0;
        data[379]<=640'd0;
        data[380]<=640'd0;
        data[381]<=640'd0;
        data[382]<=640'd0;
        data[383]<=640'd0;
        data[384]<=640'd0;
        data[385]<=640'd0;
        data[386]<=640'd0;
        data[387]<=640'd0;
        data[388]<=640'd0;
        data[389]<=640'd0;
        data[390]<=640'd0;
        data[391]<=640'd0;
        data[392]<=640'd0;
        data[393]<=640'd0;
        data[394]<=640'd0;
        data[395]<=640'd0;
        data[396]<=640'd0;
        data[397]<=640'd0;
        data[398]<=640'd0;
        data[399]<=640'd0;
        data[400]<=640'd0;
        data[401]<=640'd0;
        data[402]<=640'd0;
        data[403]<=640'd0;
        data[404]<=640'd0;
        data[405]<=640'd22835963083295687686091155745995325592756551680;
        data[406]<=640'd22836137307867241909738992724944393428252229632;
        data[407]<=640'd45671926166592015614959756397608870041507332096;
        data[408]<=640'd11419593118938734974605247813455870800613605376;
        data[409]<=640'd92102251995524685136327182220460836482002714624;
        data[410]<=640'd713798081558695355229084985473875756514803712;
        data[411]<=640'd79973270849186984475343595013176781527727472640;
        data[412]<=640'd758237586915271256831821758006986185344286720;
        data[413]<=640'd188396706326222447116603965185342682481500880896;
        data[414]<=640'd10634488215193846815532761681284300800;
        data[415]<=640'd0;
        data[416]<=640'd0;
        data[417]<=640'd0;
        data[418]<=640'd0;
        data[419]<=640'd0;
        data[420]<=640'd0;
        data[421]<=640'd0;
        data[422]<=640'd0;
        data[423]<=640'd0;
        data[424]<=640'd0;
        data[425]<=640'd0;
        data[426]<=640'd0;
        data[427]<=640'd0;
        data[428]<=640'd0;
        data[429]<=640'd0;
        data[430]<=640'd0;
        data[431]<=640'd0;
        data[432]<=640'd0;
        data[433]<=640'd0;
        data[434]<=640'd0;
        data[435]<=640'd0;
        data[436]<=640'd0;
        data[437]<=640'd0;
        data[438]<=640'd0;
        data[439]<=640'd0;
        data[440]<=640'd0;
        data[441]<=640'd0;
        data[442]<=640'd0;
        data[443]<=640'd0;
        data[444]<=640'd0;
        data[445]<=640'd0;
        data[446]<=640'd0;
        data[447]<=640'd0;
        data[448]<=640'd0;
        data[449]<=640'd0;
        data[450]<=640'd0;
        data[451]<=640'd0;
        data[452]<=640'd0;
        data[453]<=640'd0;
        data[454]<=640'd0;
        data[455]<=640'd0;
        data[456]<=640'd0;
        data[457]<=640'd0;
        data[458]<=640'd0;
        data[459]<=640'd0;
        data[460]<=640'd0;
        data[461]<=640'd0;
        data[462]<=640'd0;
        data[463]<=640'd0;
        data[464]<=640'd0;
        data[465]<=640'd0;
        data[466]<=640'd0;
        data[467]<=640'd0;
        data[468]<=640'd0;
        data[469]<=640'd0;
        data[470]<=640'd0;
        data[471]<=640'd0;
        data[472]<=640'd0;
        data[473]<=640'd0;
        data[474]<=640'd0;
        data[475]<=640'd0;
        data[476]<=640'd0;
        data[477]<=640'd0;
        data[478]<=640'd0;
        data[479]<=640'd0;
    end
end
