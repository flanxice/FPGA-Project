`timescale 1ns / 1ps


// VGA Driver
module vga_driver_color(
    input vga_clk,      // VGA驱动时钟
    input sys_rst_n,    // 复位信号
    //VGA
    output vga_hs,      // 行同步
    output vga_vs,      // 场同步
    output [11:0] vga_rgb, //4+4+4
    
    input [11:0] pixel_data,    //像素点RGB data
    output [9:0] pixel_x,       //像素点横坐标
    output [9:0] pixel_y        //像素点纵坐标
);

// some parameters for sure in the reference Table 
parameter H_SYNC = 10'd96;
parameter H_BACK = 10'd48;
parameter H_DISP = 10'd640;
parameter H_FRONT = 10'd16;
parameter H_TOTAL = 10'd800;

parameter V_SYNC = 10'd2;
parameter V_BACK = 10'd33;
parameter V_DISP = 10'd480;
parameter V_FRONT = 10'd10;
parameter V_TOTAL = 10'd525;

// counters for H and V
reg [9:0] cnt_h;
reg [9:0] cnt_v;

wire vga_en; // 使能控制rgb数据输出
wire data_req;

//*******************************Main Code************************************
//VGA 行场同步信号
assign vga_hs = (cnt_h <= H_SYNC - 1'b1) ? 1'b0 : 1'b1;
assign vga_vs = (cnt_v <= V_SYNC - 1'b1) ? 1'b0 : 1'b1;

// 使能使RGB输出 // 范围内输出
assign vga_en = (((cnt_h >= H_SYNC + H_BACK) && (cnt_h < H_SYNC + H_BACK +H_DISP))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;

//在范围内RGB赋值
assign vga_rgb = vga_en ? pixel_data : 12'b0;

// 请求像素点颜色数据输入
assign data_req = (((cnt_h >= H_SYNC + H_BACK -1'b1) && (cnt_h < H_SYNC + H_BACK +H_DISP -1'b1))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;
// 像素点坐标
assign pixel_x = data_req ? (cnt_h - (H_SYNC + H_BACK -1'b1)) : 10'd0;
assign pixel_y = data_req ? (cnt_v - (V_SYNC + V_BACK -1'b1)) : 10'd0;

// H counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_h <= 10'd0;
    else begin
        if(cnt_h < H_TOTAL - 1'b1)  cnt_h <= cnt_h + 1'b1;
        else cnt_h <= 10'd0;
    end
end
// V counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_v <= 10'd0;
    else if(cnt_h == H_TOTAL - 1'b1) begin
        if(cnt_v < V_TOTAL - 1'b1)  cnt_v <= cnt_v + 1'b1;
        else cnt_v <= 10'd0;
    end
end
endmodule 


module vga_display_color(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input [1:0] choise,
    output reg [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;

// some frequently-used colors define
localparam WHITE = 12'b1111_1111_1111;
localparam BLACK = 12'b0000_0000_0000;
localparam RED = 12'b1111_0000_0000;
localparam GREEN = 12'b0000_1111_0000;
localparam BLUE = 12'b0000_00000_1111;

reg [0:639] R1 [479:0];
reg [0:639] G1 [479:0];
reg [0:639] B1 [479:0];
reg [0:639] R2 [479:0];
reg [0:639] G2 [479:0];
reg [0:639] B2 [479:0];
reg [0:639] R3 [479:0];
reg [0:639] G3 [479:0];
reg [0:639] B3 [479:0];
reg [0:639] R4 [479:0];
reg [0:639] G4 [479:0];
reg [0:639] B4 [479:0];

always @(posedge vga_clk) begin
R1[0]<=640'd0;
R1[1]<=640'd0;
R1[2]<=640'd0;
R1[3]<=640'd0;
R1[4]<=640'd0;
R1[5]<=640'd0;
R1[6]<=640'd0;
R1[7]<=640'd0;
R1[8]<=640'd0;
R1[9]<=640'd0;
R1[10]<=640'd0;
R1[11]<=640'd0;
R1[12]<=640'd0;
R1[13]<=640'd0;
R1[14]<=640'd0;
R1[15]<=640'd0;
R1[16]<=640'd0;
R1[17]<=640'd0;
R1[18]<=640'd0;
R1[19]<=640'd0;
R1[20]<=640'd0;
R1[21]<=640'd0;
R1[22]<=640'd0;
R1[23]<=640'd0;
R1[24]<=640'd0;
R1[25]<=640'd0;
R1[26]<=640'd0;
R1[27]<=640'd0;
R1[28]<=640'd0;
R1[29]<=640'd0;
R1[30]<=640'd0;
R1[31]<=640'd0;
R1[32]<=640'd0;
R1[33]<=640'd0;
R1[34]<=640'd0;
R1[35]<=640'd0;
R1[36]<=640'd0;
R1[37]<=640'd0;
R1[38]<=640'd0;
R1[39]<=640'd0;
R1[40]<=640'd0;
R1[41]<=640'd0;
R1[42]<=640'd0;
R1[43]<=640'd0;
R1[44]<=640'd0;
R1[45]<=640'd0;
R1[46]<=640'd0;
R1[47]<=640'd0;
R1[48]<=640'd0;
R1[49]<=640'd0;
R1[50]<=640'd0;
R1[51]<=640'd0;
R1[52]<=640'd0;
R1[53]<=640'd0;
R1[54]<=640'd0;
R1[55]<=640'd0;
R1[56]<=640'd0;
R1[57]<=640'd0;
R1[58]<=640'd0;
R1[59]<=640'd0;
R1[60]<=640'd0;
R1[61]<=640'd0;
R1[62]<=640'd0;
R1[63]<=640'd0;
R1[64]<=640'd0;
R1[65]<=640'd0;
R1[66]<=640'd0;
R1[67]<=640'd0;
R1[68]<=640'd0;
R1[69]<=640'd0;
R1[70]<=640'd0;
R1[71]<=640'd0;
R1[72]<=640'd0;
R1[73]<=640'd0;
R1[74]<=640'd0;
R1[75]<=640'd0;
R1[76]<=640'd0;
R1[77]<=640'd0;
R1[78]<=640'd16882841531918873291250251565564139913819776544706983493661416868226824712570182907381492335146696704;
R1[79]<=640'd17376254537216603520283501579689306452293001289371370283519183479633757469225510874436796577229045760;
R1[80]<=640'd34993875609492269879877640612175772293536108189769042330042382660951425767464234131026187870281924608;
R1[81]<=640'd69989887206020460669837676246057714139186819084060441312854712363510673754654248902602398702650785792;
R1[82]<=640'd139983912886923018102959992846671131785595680908132948640451197120136503060027197796270466894345011200;
R1[83]<=640'd279967959273035781262800135382198899168198524485298544571700515930373495008787256882575310223820455936;
R1[84]<=640'd7198262071269318799409855121164446798547567114230080153089086747711795224138669533192284170027130570394836727058462130671723248028265349409561668293787684154900480;
R1[85]<=640'd139983912886923018102959992846671131785595680908132948640451197120136503060027197796270466894345011200;
R1[86]<=640'd3273390607896141870013189696827599152216642046043204773512990082141161526528498975571203069274147693665906583681159045440054924997310443599603611729920;
R1[87]<=640'd35091527597436931785922200359950658499183637522754949738185893746340359151868259179728727578237565652471488922756331199060601250656594990727953946003246719455723520;
R1[88]<=640'd9037418030478372893789809754239600358097447571244890132572797794402643311689402724528288997936595403426860387523266046409351022817463696719673933736609596264104853504;
R1[89]<=640'd5398696553453472354676594280158184825492050341538408280743928359512784536118620019745959807291384925905219951641259201286324079904135971687221849992726929205100544;
R1[90]<=640'd14756345861915242297113864154572193165155188740105027698815006548543594891502520906387589327368269828587018385472039908291176945245459626611537018832141271659389648896;
R1[91]<=640'd29483315222662668496425021432556870481072198772010436701438674877709814728419694543342168182917247371346995310053927534211597360926877029007300217280644241215792873472;
R1[92]<=640'd29483765114042112995891478797982029039688995258924810243178048582744057993532548984782713533436076288935278549490655657698229653982194195427350617773539930879324848128;
R1[93]<=640'd3832930474357839129121037349543383225414463114709015887515683941710662814452711128748945488227986352714398800321279009379875584851121239912806545702038695819527617249280;
R1[94]<=640'd58968035477192378122112608134997878509252648213530285790768917964786690601662514153883585459107763632213022152353768780949702552520292181341313393213890821644340953088;
R1[95]<=640'd943490471765193775298565992542541157647241103174317376495723992210612421097231234247870921370414502492010358571479763780873227829843930355302221936465334742872884248576;
R1[96]<=640'd1886981200988602496902126804164108806175360350805817776068277919003675982549533594227691452110583317088167321001600941047891977593894490450636277379572960070383379152896;
R1[97]<=640'd3773962424279222337084047026593320997680619337831941394987382895690630693048800207814379128577691854430062321891365263629323619010182594573166086324568545303612429959168;
R1[98]<=640'd3773962424821541352241178410287955813853039737950250366766022665326597488213559162460214287021879987505316742812390294978836873897295363840917419691737571129055672008704;
R1[99]<=640'd3773962424821541352036781923956016222503329659329542823059881495925074378810958895730909880464227005408306971171464264419515994128038312327434531719851642681177759809536;
R1[100]<=640'd7547924849643082704483096674982336517864916914444123130113638903022824762328455975950032522258651937287716530269831980658181068577162032725125929714589745128512501579776;
R1[101]<=640'd7547924849643082704483096674982336517864916914443961812143709597601302624113659307813771068945706182681677176705818245231324436046428212110097932628028337816228927111168;
R1[102]<=640'd7547924849643082704483107405992978229088212288684449322916973140929373371023900034358308446617284891656004160276471304627897791480827554457603672534200309316988392439808;
R1[103]<=640'd7547924849643082704483108808340959816350347479636481134972745833039719508402655645849914123990725125495364512298939400958445788312811302979689918647236625968400282157056;
R1[104]<=640'd37739624248215413522415495849711553578621665444774363561979138092520464804527533225750884655616867691620510221601371360687264190554535020498541573853429516328605484843008;
R1[105]<=640'd37739624248215413522415545797688358634497367550330047354851647184642225541918966967181495622494353936044774180497487518991071458294058750436894175742926775455456260259840;
R1[106]<=640'd60383398797144661635864873277520806842662972545912793916535700945414442255229046505710611091203906314542445584901940907051525308695458223181777648088362650659232208125952;
R1[107]<=640'd267951332162329436009150375201389770156414028034229815748096745938089904098616873341985331100753434283129233989503499485142835636640758871168235051573984922345331704725504;
R1[108]<=640'd384944167331797217928638567254325188915106547010127757842460765775757830629737259740330917657811595292532761476854576295101355691674130680927457015982762275146906912948224;
R1[109]<=640'd262290388525097123980788043377327115993616073363340456037807156948644134685732180065371900833633259095032835290590200758583585182548368709592561783017185739087706455015424;
R1[110]<=640'd35852643035804642846294768518964313237113891764081496619525460877729467999901542451321174900574046705825840377373443708750911134247760717749449227935477981729369880526848;
R1[111]<=640'd37739624248215413522415545809703874953572904179379589226729915759433353009108079348981849307180444087965678275153006703525580235530050550097252907186061313066356627734528;
R1[112]<=640'd13208868486875394732845441033363370548029043512633319992764722898291555983868260500632464438561622074669489734522337856564504778392356978473219597666254945222055459553280;
R1[113]<=640'd13208868486875394732845441033458731788656627136673069598381041728670464684307059057678291281702717869363370412195381860320762527132042222918032022934277294216509621534720;
R1[114]<=640'd3773962424821541352241554580988222373238566301575694922763761823375714529343139373667337695032914740920599010876043603372735376318391774062325040118016906109412505026560;
R1[115]<=640'd494664576908633889662357283593875368153082901703968732300536235555611768390623230985577421234775293200133392978893820323735158889619997185778094401543388388402620170648944640;
R1[116]<=640'd30191699398572330817932436647905778985908530412603599683929910711187614324406694246562492114351068068733201713747370258134860743292461427659515877911997787405467611299840;
R1[117]<=640'd15095849699286165408966218323952703422240845530939777179562047260894029200075667506315016018088373526531732291985486985900216673079491447106720912438561959815672078794752;
R1[118]<=640'd3773962424821541352241554580988082820203501545052500149135732079031543003940875445723231065339679719693062599272252018355791551354597381259474378791570874651348219985920;
R1[119]<=640'd114162363350851625905307026074894947879523447242233665112720182116843043370070667198666192588357291126548046853882981910832507518409699379321195286690463809447452538306560;
R1[120]<=640'd13208868486875394732845441033458755047495804596094135826496320509939555611937326324490655200186246302730782463193546872718226351104011505924633277407421449879849468428288;
R1[121]<=640'd109444910319824699215005082848659774577751537932656597625782891154551708382745275092804037235689830590588591176018949690902718872273678240458887746701636124097496651661312;
R1[122]<=640'd49061511522680037579140209552846751299066297163958125842546165450123642972241091639910210394569706649445418241555447757579082949175635522182960942947409809636490028777472;
R1[123]<=640'd3773962424821541352241554580986780325209563817506047928774075553040949359419712918877980692758203240983190088359865058135759333670548219471129103857773016911634961006592;
R1[124]<=640'd7547924849643082704483108908795328011657325582586775144702588609955228011860132830201590841186965684020232332459794831810923648175255374117424031698289281313267045629952;
R1[125]<=640'd3656026099045868184984006000165666128851738306151946357848711357077901061516630121305453775700650438662766134099486665792405697283331123442081417263972497845462895689728;
R1[126]<=640'd33611852846066852668401345486902952758411111172744483017997403444874316823672198769813835078572798123457657600904405531780189519020570112763770567608926562841692886532096;
R1[127]<=640'd18869812124107706761207772904916783120413208954036961130036605591736809431785711143840283517342646457970037890916004643048509736377474105778956550054312761561560268144640;
R1[128]<=640'd185865806667370666704658163917099262111097202483365704411326239783310869003697868734999350885519135649028187584017960373330985673861855838803744600728462167943462531366912;
R1[129]<=640'd126634191718200095571205598692259648139423039230781767198281524042761496237229739046457075954993466026319569441916455593200998732314443958086731599424586975942298031932303212544;
R1[130]<=640'd127625445585483001975640383498686916602289519091634274857645010779410933470404914702012244043103421668150061023989420316448578494007399830950118720276358661520782446983913668608;
R1[131]<=640'd989563117374545631949834682781413136324888368291699895616493412374865687086163235608066548887645845241413962373664106438634377708494696894254170123139281959019286714652819456;
R1[132]<=640'd864207181471673314393779205819306796797674234679428569352392620201074744709512572253185407726129358871195634400538544438769022226283005669222217764349269119333578965067497472;
R1[133]<=640'd988838538701141196190014525815660117923232430699839514590704073558041621317230849949900602531405998915854924247138034894420571499022204488961910993217279744314246835671662592;
R1[134]<=640'd494660626041720404611254155716423349518150528955765706083801460981631569952131186357411272857382886497619624264873111261866751362579830868032365221276015122416531868624093184;
R1[135]<=640'd2473301921361262822406306388709165115476448508212554215205264321986648920033353425879015850099166858682996370323065476772999271765366014491306192427792428143446522393278808064;
R1[136]<=640'd35600119647292943149374435712071894833486963654283303774604333011257152947018463105781274701024510001793250134448700645892863779031012518370566958482204171310079191667793985536;
R1[137]<=640'd13546093578445622735896875748957584653284662170697063816960161211424734094747645477424486915098336682586597144648676278018721199806331000904638490049040531279975616747662746830352941056;
R1[138]<=640'd8716903953620346982776979291886296691243025938970103656204372261725344438473708850141751194805737238862334093013975647246008977989806115748412784706068345637962566976767530546794709647360;
R1[139]<=640'd69687163640560300729471852577682079556763804105867268700792490680318805831935500552991634367067482837172230162264056931771397949060624880739656115885346953835963477290395554408243031703552;
R1[140]<=640'd84951994920127167245795661449134002579916004397648589072048425882427965634831205147388586648011726525661880623768590464785096926686464051805339031704028452829382058653947322618706132992;
R1[141]<=640'd36032387946968732516894647597529525894800379101298188416156028443377339473746287758065488913459683202581200125085680187320714418666466536117790268161984134672388412251805961948629737406464;
R1[142]<=640'd41743188832620411102388454950311863558536079019024779916254116728754394100410260772804307604599959771042461739870569803206761955406745600209277455207884972687047233184058924068347741995008;
R1[143]<=640'd146288146384117230735501184067038315021052045462417334428498404827276717868990177944307195886622874795196812754873253524058493796890972757132623826839161004334718308629165356254932437565440;
R1[144]<=640'd2515463309754715206738884845932258045548295545438197227929162012364016785570042669972198037634730373457314044262887271327437810769669555842800594749100989440399646687632102387521152876544;
R1[145]<=640'd38235970585843011530128796468778572394367750137984243378227212408582334809800121773365006716769956657767053397922068534200150875686127929762342336659666332561466873978608872017996283904;
R1[146]<=640'd3709666918579618923603082041049933443313861822533423924008426855665721830809856071287766382639745409752443254683650647472086925164184724567467226185316854294443418073555241475910926336;
R1[147]<=640'd423250588025872425829673858088357656544543210296203717633211286113688454057318389670575485568756261106961502622592359077831306659265956937670938725299436358293087571208648765099474944;
R1[148]<=640'd132784498204192497493081200197489918917253939904642087032931168842936093653377995003598981460716309330066519949203589235503540676800039982096086538557580641000775384021416167421771776;
R1[149]<=640'd1429985148292108422111989037314198555608244475264840743002965374416195796023358220515609420650339060165908065778536164220854014062323207107554330624753905345517789904896;
R1[150]<=640'd943497804467456607174601142108679510363963569230895382130273365782047960199768982261120718927434111632298466464580606600680543918385966733592863930328930694327340892160;
R1[151]<=640'd3599131035634557106248430806147366919947059365515344066424713359585296521144927977702057962751543192483164747323287320412532853187429483518639211973271327357272064;
R1[152]<=640'd1799510599435997508246495547867293355409525891022021141497243865394784510061283201048142321797668692751995756793681138754279138560806437422291007643029538902900736;
R1[153]<=640'd787309914045059366991844238844696376324808990631507883752718666216640904722306321614797827557374601919578451795130429988365817233975106276097053708535839661752320;
R1[154]<=640'd899288493477109872662629004359896354019557643402173546068400355376537416299846725719804762456833620804324072880839764153557428325982637244898146844468796238856192;
R1[155]<=640'd1572907061073916146859800492370705373181927884911773418699542426679212612037056197419614153014148066783158971250018740208025102569977449847856222492034140355952640;
R1[156]<=640'd55399775216961536726118311839822379877535372871657305895882198179039631508593481336660391464034892061612687410072167077610102937664985592954341170959650375335936;
R1[157]<=640'd460744172336440271136525261499083098427759019623958011027976897692335045361315453567379173830181283117692035682419259381229294444160733497970353696219179247334326272;
R1[158]<=640'd110760506897231080609482664529076911826089059839001283812670715043656414945415668021808283273774975579885158677986639544762761034419269829003895430671881113436160;
R1[159]<=640'd26392143654225887212355103350636745250111612811334505221778640119345920631164788515185394484426432938216849784292609011395248041232187373832124570909637374640128;
R1[160]<=640'd13292071731891332601410501446835312474195285861784657941030278436398958099790390569232951864478940267189158208927444007399362451094996368168237959080372189790208;
R1[161]<=640'd90617152575602520430966632614396596572640198059986375013958942282056603073347689108894059585045249395152709148440541644725523715840873062007062178106676911013888;
R1[162]<=640'd62428577183691204288822202457831746279954826101164132013793665488078934725737677901507300392326959164944773934897712067575012043788187796097967370841152697663488;
R1[163]<=640'd13221707555874993851831937508777669841963587020265443113011597842767143959947520559954741149661051882998538328313154453384810836690167917053619982541241236586496;
R1[164]<=640'd66780858900214010848120727547816797379380681642532168951192963835089749158678068942064088888560114893767356292054401877937382619871823210860176498878642223316992;
R1[165]<=640'd57118642785772247731686602616205282442626470820874164885662508164690576553576245078539276988798665096101081729529045393542278769653745533190081394278677209939968;
R1[166]<=640'd93854655509598179697017454094839398562166482226388367928941592756743292583545150522067222699505008715380947746670491404302678797092911778423786331852242944;
R1[167]<=640'd93854655509598179697018156969339303541592551539476417936251094989371144614980468785447854038601754679982410360722546519780904835616249217519692638171693056;
R1[168]<=640'd3351951982485649274893484072376574863183992413037164767199874001731466986990387670790757409025015606220214444967615215833805606854523904213679508769734656;
R1[169]<=640'd16759759909306497824151536243907306590373731475387730612108157411299567610278214473491857715478224693068173874972569020027199275449898389191253250308833280;
R1[170]<=640'd3299373145846317496106341755496024228864913695653428733830660581137926145825172753697229353324679236429392226709888286868590766578427225785236726074048512;
R1[171]<=640'd3351951982485649274893418048070264770476217844893608778950749629947027218837950491671992425468156003403001080714912914343379759826055674120769113337888768;
R1[172]<=640'd2506496564539973882529117739515470638021442404316997588852914266683763909510883605665805099510711935365907531947479898956727516279565683147631470185545728;
R1[173]<=640'd378383495398579695166720692423753594422214543544973124024425387552428874418724470095523288371854995921742308180925078440490837549049001671483576989777920;
R1[174]<=640'd189140600751543525422390149556078449160180380276702404548001785819699434924191753642646955696286683539546947999919195043014262248476536526075875383312384;
R1[175]<=640'd831434730722893147924732835454312620850242799430748269949262911667500122105929708289358936461956286373998529595200160919254835982443836674097828583178240;
R1[176]<=640'd366619708282073872912398845365393397312449744247983231320974983359283611140113554129790830043661323445756502819043711616198371704107815341084370729435136;
R1[177]<=640'd418993975578155631708325781123345295347096231320943637234399580612605734743354556961215920745785730262768553711648609104829740292571411526927131500085248;
R1[178]<=640'd209496995040512528251947650201872315540027470212021156494603229380330831843245823268562611263294851185396152580519049974340437479667815088528492010143744;
R1[179]<=640'd52374246641601417351598368055337720440514948087390698725170688742030775550663247183096105659333938125195753377444766765107572364849470645282832885219328;
R1[180]<=640'd13460182177912996466912001323033343811539640460493783148481621943051488829986592373866153176681668301441879597505769311598583586771662137376525914503905280;
R1[181]<=640'd13460182176157039701542653565675586590846777943079752147345654297054416346956772771670445419888188916482920978030423828737023701415512858137901911014113280;
R1[182]<=640'd78561373809141718455227303749712322861482758284526980481796747563300032916890797776199273466422354845839766356792447364357498416506314982227918440103936;
R1[183]<=640'd183309872484381883111826312374030427832628829701504869256676737221378423579535693729635977682049486970420258084959353541079689436309564716166620192440320;
R1[184]<=640'd47464159326983493167350844443487956001198179655684600374491865884229920117326851333856197922160877297689174158175209714073391477873123540349349345099776;
R1[185]<=640'd523742495702508470561775954749228493509753459360632281090514814793088483471742774911216587999644916973894790027374360869920711211766022514361655994875904;
R1[186]<=640'd52374246604589812639564466387013475842412952490511386541041868709297053315396180816076045855739256475637998657849641174190363218284181620710082816770048;
R1[187]<=640'd51146715761383061972610112734453395345878801060271735220702246953635220473265355158939323161846321142392690283810914622815580739502670410518790469058560;
R1[188]<=640'd208269464940397831029485788423408317342433007140478912848469328123085163578284610277856595308403276937537613187321589997166933778667971313329738667261952;
R1[189]<=640'd169807125297618169508792228107173599640441281155414337277537644094043318032775777442603426791992933158620900440951515828282117663510292444687097189629952;
R1[190]<=640'd5929798832307834260607951367670136005075353593694411536995369477549263729448957321474810365239343542325114565164164326201875910104629505312917169373184;
R1[191]<=640'd40037973545083567590412396543760594927635048350096437618854519449053852504727469155331094291630645651712582284481140760266020900434776135793493680324608;
R1[192]<=640'd24574404588087865341614863051656526265652227735338373444530137867720006391166268742517852926366115283089481574050392236607956946865571792863329517568;
R1[193]<=640'd72401034126981983556616073994384812564197133372177472464929639759741967984540230732971615591484300282140833994231814166976769967521792;
R1[194]<=640'd68142213476812411932303629807540896285279230034736105046331601631854073669794675731473162246052968177133659713666284415019671521067008;
R1[195]<=640'd277345481707382766203441739491551567963118378348623124239828468202470578796352241211974025222452907580271255860022799727874505965568;
R1[196]<=640'd186070713484659809936583493090698243192857409754921127304416411667826176652771167216988888223850945461230700810617858697788130411589664768;
R1[197]<=640'd713475062891440151854406384282803704697664946923934833583686113989643134085987758449142562883944375663502084293920158784516259840;
R1[198]<=640'd26114976232752529184397838890140322703896830362617776630122712727372094106359318332088176977935341430962662699435440377920503685738545757303538363477231778058807714668575422089325046661120;
R1[199]<=640'd35774604030988437628712220594762150749175765729140835127517439225016172364438616480247540171929154933700880260806079696465543199561697341625729076835048961899059954689347973100932171237949440;
R1[200]<=640'd67110585617167563430353237339878494508411339295364608274438735500676496793282331403363486092316889027425598735850240296217796465235260903786967092081303199764542160905512468514755034809892864;
R1[201]<=640'd142576167321161604828319839607242888831054489596240823244511488292152275690812112912184359781896717265590364528192081639227828653440388728938475562807994993630467097556578371457487784980250624;
R1[202]<=640'd1140610154405313836574276627074938274799795604647604377265919043523131936527600367361334728255066740822872915125952937068570624220161789489915948901276729027205321166236624966552445548341755904;
R1[203]<=640'd4562440617622191102815960691767740024070776219299670556051447481343223299931694999295517774555548691483781104341791192895234073448408702055306676059035129263358559057261984273140420383309037568;
R1[204]<=640'd4562440617622191166318041269987329144104798491094086597478386006369356244233062850705346615446776351860154304225780707219601307817481793447624864210297522632074376327075921385561720797433692160;
R1[205]<=640'd4562440617622195218517506404963739057862977246738736335561626843348805995458420005874548410036091090173262915465741202135823609512577315503871783178740035132108613319102489706259943376342220800;
R1[206]<=640'd4562440617622195218517506404963739057862977246738736335607054263617149297556010493931931376600606764624684663654229393745544278565043589736597925382207499025817185521071204567551782543641542656;
R1[207]<=640'd4562440617622195218583203542855032449722798228884580144376764251169104094861401816270721125809163814038076182642357424378731758549711137843125540036573518511537799821116306648108035484749398016;
R1[208]<=640'd4562440617622195218583203542855032449722798228884580120565300506144203498323541033669560061396142527611675848160515558991841966732567357562362245400250555140180094875320499583748495474631376896;
R1[209]<=640'd4562440617622195218614119843039170516480387231136911406648677407898000242280901477777425207990318073349872230995781726632611464110005832157481482702587330248644523294155980781032320584204156928;
R1[210]<=640'd4562440617622195218637307068177274066548533155357627968540465188225160004512134762798517914635336858409846085461193612627313818162225700265299193776644149974018471938764738153319242990134231040;
R1[211]<=640'd4562440617622195218637307068177274533361530322453786347680404598821024011230824874402150646912594455846765052932351338596835557162102830009255634085352585190874536913985250622771313737696542720;
R1[212]<=640'd4562440617622195218639692212429762034081651829005388917899573340043348606101430552222004496996871026653507928499728409152962560727172630105802954463684301866724169055576491804379820759713841152;
R1[213]<=640'd4562440617622195218640658346810519055107599269506024591092485472543013427849166500457616522984776556170376851752093786779138736977103540874702367325797199095066103554693479413499034899065077760;
R1[214]<=640'd4562440617622195218641169726097297537173342080030827012925479252858231056638208541423098912964112961745236635052937375846028902490129509943332542960617230390667215702002453166870522205065707520;
R1[215]<=640'd4562440617622195218641170719752592117233186188169233758989725481899821192110192307791458210583774040636797552671125054345882110945544179574307023271175261785029006834965018091386904806531530752;
R1[216]<=640'd4562440617622195218641171605678696538679417072872833864225511632178887255270245674976235291660837295364325134792564579390905953938347600138445505945800341208996246503523712407486121477230559232;
R1[217]<=640'd4562440617622195218641171605700291324893225233858586139611605440631577726546826906769721952250310738752292479697221906270581586342870049271280282239679926473565021177379356934749675274469638144;
R1[218]<=640'd4562440617622195218641171605700291324893226870562621228159205487998571545098480777102135584212971571585535732385572320189870559946690193355364561789859631201580709934418335934424211294053728256;
R1[219]<=640'd4562440617622195218641171605700291324893227689325465759386699958069748183560759949927210647953610105472645632049195862621538108240213986538848281675787644930745543083827053171117817250527051776;
R1[220]<=640'd4562440617622195218641171605700291324893227740622037938179084304132153863522068685988175328224416056390312792613304274907926778057083872078148351774063777117699170501828189533182921402413481984;
R1[221]<=640'd4562440617622195218641171605700291324893227689896745744094526536412580476612909383879204108061299826079871355660638890825555216722230003399467312398035973325962955073694032646640597303105159168;
R1[222]<=640'd4562440617622195218641171605700291324893227752834318267015245913296962226472935274076691262329783198551334818667758517170849883967721347262528942951306731664641879268820670316771717500660744192;
R1[223]<=640'd4562440617622195218641171605700291324893228466491010857653597944981141735029098098652215460683508054161489044704740985279828768430658956401301485857021801467167126151391494481295021168897556480;
R1[224]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360263644831615583063638016;
R1[225]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264679866896343894364672;
R1[226]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264236280346278147395712;
R1[227]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360259432056436581411595392;
R1[228]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360259505122836935870524544;
R1[229]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360261643720170389717142144;
R1[230]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264462433106403130403392;
R1[231]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264666067866606710597184;
R1[232]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264830359180392559347208;
R1[233]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360261046610411662312736328;
R1[234]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360263257621125137390652420;
R1[235]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360263060480554911555159040;
R1[236]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264148964556015625511938;
R1[237]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264032816722725115529216;
R1[238]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264484617837276351808256;
R1[239]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360189139323445326404569352;
R1[240]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360186780734841324264802592;
R1[241]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674359961395510364074305935364;
R1[242]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674359961985666560551053316612;
R1[243]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360112727855892572893906182;
R1[244]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674359999946490930211456163872;
R1[245]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674359034534123350236493918738;
R1[246]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674358318025707773129925206282;
R1[247]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674359263070532816223651436584;
R1[248]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674359801790413176107946086449;
R1[249]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251974391945560573087993511143196688;
R1[250]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251964250743325628979957325526501442;
R1[251]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251928756518104792582534768476823681;
R1[252]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214186922746396160252355242820486381154536;
R1[253]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214186922746396082793591549495810308313128;
R1[254]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214166973954542095287152616408000905648484;
R1[255]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214186922743702368842360408081888034834624;
R1[256]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214186922743702349336966193388561856515200;
R1[257]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214182921990078895963865608719380513661954;
R1[258]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214184928914226730314291044530883444052032;
R1[259]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188199904375894707981233222158984909712;
R1[260]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214187919588798666729042175762830592033568;
R1[261]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214176953538963067619597428424458082633304;
R1[262]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214181937963703124987391607803729929257996;
R1[263]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214187540633287539901194772522192571425724;
R1[264]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214177617423903420916740303827776776333204;
R1[265]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214058475640158074573627246666618272377873;
R1[266]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214144927017610850276499250787129663365552;
R1[267]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722127053563771194448713465089674254885459896;
R1[268]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722127075290916160888371216010952917762385553;
R1[269]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722127064667545083002208213982329961937729720;
R1[270]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214187905360529871447832775551307199609180;
R1[271]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213501995141057522850622242600037583046372;
R1[272]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722208403409424064296239542530468759006238320;
R1[273]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722170631724719733478303756356679409598840700;
R1[274]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722146131393975754368838539625657684167860062;
R1[275]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722188324412994355579511890936616397529796534;
R1[276]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722212826530130561962365771130522288734314464;
R1[277]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214016604651774110665181763064033060535770;
R1[278]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213932785610056767177061955833218761997805;
R1[279]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722192239919632542975121992509999434871045164;
R1[280]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720820306517664480352495210210569631002224531;
R1[281]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721516896426993833084081282173159888023682801;
R1[282]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214166888533424838835473961047985538432796;
R1[283]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722116037929822899594895946500745367906254750;
R1[284]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722205978544728737778230823271512291779182461;
R1[285]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721945864908218823708339970142668970868793228;
R1[286]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319699777287424039013506604145600398817685993926;
R1[287]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722148720885921115933146682931444476982393852;
R1[288]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722202913698084946006202505227834331476556286;
R1[289]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722204616366861028753105935840208753894944634;
R1[290]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319633009716613638835335283000442531033763645324;
R1[291]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319655311141473849315152462405290986244500748142;
R1[292]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721418203493840744050193733446696857839957950;
R1[293]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721768553838945138836460828332229022345917434;
R1[294]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319621501315706560098692719812152254274169010034;
R1[295]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722197843825679412019530812065712449881955296;
R1[296]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319716201308366967888909062665138664326926237420;
R1[297]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719382222299136979682111683225287639929782140;
R1[298]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720819149808685789807483248799395148612566966;
R1[299]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721516970847244882193016562364282786991964024;
R1[300]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719402013038837037807077104080203781051572156;
R1[301]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213491793022634306072813209966102441420688;
R1[302]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722207706180636742905085542864760282082311990;
R1[303]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722178152333194337406024974410634706481443695;
R1[304]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722077880734816313962149089093689768809102428;
R1[305]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722011111286788916558983926882475259235728474;
R1[306]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722179214506835164403272100958540674659318862;
R1[307]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275164626427508419004221661452227775630435243888614481465191890716081457605039302880649817928961296753324492081668757637889215;
R1[308]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275156879677874158278452693694711766594812254771235993794653398738011835662173252357431819538942812986062035277576085804996727;
R1[309]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375425444049190546360682135110894540349921527696560300006078569;
R1[310]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375425444049190546360673543184118676958767455238794017706356785;
R1[311]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722176033833416465654789708068526836552611889;
R1[312]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375036263741596571974917100127374638656482379984752502474852980;
R1[313]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213387990232932747902553198353896525586654;
R1[314]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375425444049190546271480755111867404815378748373416514844131534;
R1[315]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375425443666066661144211542588352052718770140726171614463185478;
R1[316]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375425443666066660430590277605204885406327431501420666139107936;
R1[317]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437997869537434483440965232039483611225898960627593591578688;
R1[318]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437997486413549289258477871748742782321379216127869811869265;
R1[319]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375325009655176589035520701840157942505459696629126364824225282;
R1[320]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375375226421169196456034794050374182876730165181743089671773106;
R1[321]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375381504337042839235740020620634939724234630448465433966948761;
R1[322]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437973636951693759215471621485624314698132933390746707063369;
R1[323]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375412888313224231668034729863607957137403278675879429087706848;
R1[324]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437971433989351089425974800965554546043078024151493664065584;
R1[325]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310687842003082082482294241307813945815742178344415999815958063269707282551;
R1[326]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310687842002670703622796327384590164303053704278574776397732934818008544999;
R1[327]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310687842002259333711527903952843839830107448310441215473085787324211425007;
R1[328]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721272590821756336669765310869126698118508810457488391409460074638;
R1[329]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310687841975931260831072719270627010287693820547311182977578807267161553110;
R1[330]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688273361817283876507011250554105820014178005720062364731897594901194459;
R1[331]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721169746786971651779740786048625888654312494118151275913379870395;
R1[332]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310685253848202014469389162077448973096956456295076339560176361780528310127;
R1[333]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704714793405547407721334854999689768738266915921592420694258393445455;
R1[334]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704695047360370221323731807546245822497750541302744294202535475834431;
R1[335]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688271663965211671482487732660789633351281808525072714355039807181978879;
R1[336]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688487341970177253453589821515372270826489071765258977994226075428616318;
R1[337]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688489028599496239960307060533294732121068793003760237261627806423858942;
R1[338]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310686979073328145921129542667643212358647100988747985578537150356755192575;
R1[339]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721259736754930212410621153795162869443809370069451731627510739583;
R1[340]<=640'd2281220308811097609320585802850145662446614253624279965289596258949637583604338693252956405658685699889321154786797203655344244310012926755940702597089085220109337508039367517704923879589163837;
R1[341]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310686978863382066255256565514878165365073654245435733259754882915235146367;
R1[342]<=640'd2281220308811097609320585802850145662446614253624279965289596258949637583604338693252956405658685699889321154786797203655344297176889402355363828311140311407934225661583942084602223601762049055;
R1[343]<=640'd267330504938800501092256148771501444817962607846595308432374561595660654328633440615580828788127230455779822826577797303360558452142358729609429197224890125412377457502217307726813685387246447;
R1[344]<=640'd71288134650346800291268306339067051951456695425758748915299883092176174487635584164154887676833928121541286087087412614229052264035217964588634303948912679805404111764958463050066774470441851;
R1[345]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817792082077443838416964060770643043543706307114754240037051709172390381765415073475791305348948198882838319233253177;
R1[346]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817792082077443838416964060770643043543706307114754240955416825979597385681886181518490359560765752977530483295129463;
R1[347]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817792082077443838416964060770643043543706307114573051981156820645385025502625903802219701289021919620710067402456423;
R1[348]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817792082077443838416964060770643043543706307113871303425993366327586219676046593472104485166777235041684018689359655;
R1[349]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817792082077443540950865490281021328883403419118201360578095801834820372607591351234514981211154205142070449669283627;
R1[350]<=640'd142576269300693600582536612678134103902913390851517497830599766184352348975271168328309775336169850444818476779194807411517139937434963518050907542997326976938800328990114663008531063248263981;
R1[351]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950541721000272732043598020626163579604383946085991908057463519719591098510836329040308628018739805946397538334286420795;
R1[352]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542336506312825409810385901238386153832080704874333529232094844993859700580848883930122661945623126114912810900528575;
R1[353]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542335454165748327133099806751078792209092440568577739250023843363293813470631038307160459096316405637547528983157054;
R1[354]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542336656619550707335712486165144348349650456918030091207192341788866903703910975283029513466277052047847771275267355;
R1[355]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542336506312825409810385901238386153832080704874346143207509262179270800176421740584364015713364456425601846159081903;
R1[356]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542325796958647961130866725206864794455235871761881445163499038825807594820431231263364931224874939066848994145601572;
R1[357]<=640'd249508471276213801019439072186734681830098433990155621203549590822616610706724525335281268785676945554769452406557015888208369032426248222374689818742018736641553013829574608793747345644716812;
R1[358]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542278638223576824839655901031209757388523718044873322051398304505731583052083113343714785941863677472646327129082240;
R1[359]<=640'd249508471276213801019439072186734681830098433990155621203549590822616610706724525335281259817948973944420562479297884705964032559876123936187114085526068307452627404541446372507373320596887552;
R1[360]<=640'd285150295074505543140848360535683730178344941501705716678355937916664939445905474797115792484326274011133112280928314147124919661344123929133812726270161045630513877448117369836800668235470848;
R1[361]<=640'd271628677533663022093418193340795337098266569918999657935162972148527388889994419472617121180221264828010517509429957134852219308457430164570773043293391954299529386113732738560683553947921408;
R1[362]<=640'd247285000165164537920220770452936475563626198097002011085375149793516553308292650181284251201916848743877190304448616682639553378700188797596343356425232291602671589023689426983737804867108864;
R1[363]<=640'd262876075264417236928029318178957261923605695889511585908713443251702251934986278714534512862948397936153609668688978966360299681792231453452432991000787071146550720511737981899144734479482880;
R1[364]<=640'd169309859430774352527134496176902105267137116727107181426795899286127211470681445746737889316765170653119305962236865191092420055600768203177594732267278808376656909907188146296997443128000512;
R1[365]<=640'd249508478711367666285013267661248496664519222112966977801975765003049745215580112403262032089390366616863903496319431609314291023725798398634889108851505200842532360080757704950588545093861376;
R1[366]<=640'd213864408195929991658296950060417643825546806477806856220519539611393597699888271136703135698354629611764645181929804734014501513287239261951405692273193255540243438429469748815383819681005568;
R1[367]<=640'd564236863096669394085222334476994753172538375464927942591530134071789338162186813788856067625610654573685018354406387828311354566941478337733802625922199830649084780677063454197286912;
R1[368]<=640'd6482858277383226120547003211261904050071842677360098449341056685160929146211565258006081058515518663212310618028731722486088823378313758385088670464847873921677159431940394910226432;
R1[369]<=640'd58645000115691914402798803064230074297814728166033561727302886132199526665786686404759822314157434173517336352985392047241518887583439711573851598095543892682427425966257398218752;
R1[370]<=640'd505881970696738014159950764291511603336548954821276561557342620243938144915692932647555708473985361828748086659365555844192909635354997091855754207528520947927795486092966232064;
R1[371]<=640'd142352111545703422611150154651919284852536661326147506332575600677216354846600554493993840446054623625630769280627303337210067371698724077458208743089748730519814753423378874368;
R1[372]<=640'd3214563011471780675498937237636450732696463906011988779482109045527164746523830774758907806106511622124536667463981393559676235827605759953759765188350529126815002406292684800;
R1[373]<=640'd48302945075290904335045575516216672583735697099743003668889076205086943610740303224674102260234216891053381487042577224859138528984513195558552365544123831882653157413617664;
R1[374]<=640'd14859977047679900745544283087217156626910449843038948804901410214726098695020906222474398837811228014510160528641214888375755014731687595805900289995810559967890868535296;
R1[375]<=640'd5660943637177393699455536720100818050193677157436056431377806406101097625784187568667840008499813684632261906574118493099120402227241778763206687551032728108498753159168;
R1[376]<=640'd7198262016350785305701710230712284792465857640005420166898579213319179256347469739074110125139573717992177492965828147095079404346178715739095529920062510157438910464;
R1[377]<=640'd230231858517471542344904264815464145414485715513885035404703297290320666147418400704815832557065314656611719571651804165721672058830370978199780716420506721183596544;
R1[378]<=640'd22494170814556442838141900128023984537172369799127000702248609894034600530124055419476516568134399766485147578911228639154744329200426694165263528647829755011268608;
R1[379]<=640'd56208963345897931798948343583298334529644141822409953282690189278597664522322832378022201219745068678579001162317432239785872355773369969612176874230502674923520;
R1[380]<=640'd27665134675074856604053600060717870161138720570223011266081404200161892775609726152315177897090003714749275197497720674520837556950737012593699997029792380616704;
R1[381]<=640'd82377676670066769256322650007099507614808652818759580055985330568799349450707792513845004260500246733868537132510204674492918724427230206095704579064624840704;
R1[382]<=640'd104748499452676539840414291451978951361386593053120061915311973266776845989151232475046279419543141799901558589371927385379397085234938993610233422544896;
R1[383]<=640'd104748499452676539840419595638108801551851071999286688162670244794595569109209744626989164428687794729363479208297949371461582190924824752687819543019520;
R1[384]<=640'd50839847878886953418642038546266320413706841100295486075617400277251444853731244775270849623214390706405997878746955751252505088879823481535066441515008;
R1[385]<=640'd12786682062094304179578066324113675056571805301265638241699418836599353402436695778794203655553408073684945971846516813779816934545463494050043658240;
R1[386]<=640'd3196670515523576044762980717278705342867423488865123255451604550004681459344011292690555809174489174066598042999651825531142301281074729663835668480;
R1[387]<=640'd1598335257761788022078983644586552326866501000887474919456756524594912664642929243487846657849677926315457489534855124173726166896731505203672514560;
R1[388]<=640'd399583814440446296138488973865367967158397847614501585450095535528839624998095764734895419071795610464505376786058351561459881137947933841477861376;
R1[389]<=640'd99895953610110331797338381303570107426637226930771033299436291571638322006813859116808836637940487034630176080156207159828078109737584617832054784;
R1[390]<=640'd24973988402437083010515827438501707679946830322992548691912099002764764224591311375779434656651707616927305287373153010316107125767121416520466432;
R1[391]<=640'd6243496914561271043087830622693023028094508369726644168321977183907391479478789817124881540430995595848965081141128926164725876560677414933364736;
R1[392]<=640'd1560874089087282696015434635146594671243938594643141942746044026905636802946086318498315073532374999977261975877097815959990307941931624303689728;
R1[393]<=640'd292663740521410852016660759688974860964871608660641859011100476471441147142124802838247812570405241784154525071482851478811994448348730263339008;
R1[394]<=640'd1523919142907141231001334272261530423736650875215801552879397600334925881666225470319661295108886201982022819974525580347471176581963499700224;
R1[395]<=640'd136516083251477377870759728130170582727293675202942817444473409593224246211861959601657895378109835169840316284928;
R1[396]<=640'd0;
R1[397]<=640'd0;
R1[398]<=640'd0;
R1[399]<=640'd0;
R1[400]<=640'd0;
R1[401]<=640'd0;
R1[402]<=640'd0;
R1[403]<=640'd0;
R1[404]<=640'd0;
R1[405]<=640'd0;
R1[406]<=640'd0;
R1[407]<=640'd0;
R1[408]<=640'd0;
R1[409]<=640'd0;
R1[410]<=640'd0;
R1[411]<=640'd0;
R1[412]<=640'd0;
R1[413]<=640'd80695308690215893426747474125094121072803306025913234775958104891895238188026287332176417290004307232371974124148359168;
R1[414]<=640'd10086913586276986678343434265636765134100413253239154346994763111486904773503285916522052161250538404046496765518544896;
R1[415]<=640'd3782592594853870004378787849613786925287654969964682880123036166807589290063732218695769560468951901517436287069454336;
R1[416]<=640'd945648148713467501094696962403446731321913742491170720030759041701897322515933054673942390117237975379359071767363584;
R1[417]<=640'd275814043374761354485953280701005296635558174893258126675638053829720052400480474279899863784194409485646395932147712;
R1[418]<=640'd19701003098197239606139520050071806902539869635232723333974146702122860885748605305707133127442457820403313995153408;
R1[419]<=640'd7387876161823964852302320018776927588452451113212271250240305013296072832155726989640174922790921682651242748182528;
R1[420]<=640'd1846969040455991213075580004694231897113112778303067812560076253324018208038931747410043730697730420662810687045632;
R1[421]<=640'd192392608380832418028706250488982489282615914406569563808341276387918563337388723688546221947680252152376113233920;
R1[422]<=640'd28858891257124862704305937573347373392392387160985434571251191458187784500608308553281933292152037822856416985088;
R1[423]<=640'd7214722814281215676076484393336843348098096790246358642812797864546946125152077138320483323038009455714104246272;
R1[424]<=640'd4509201758925759797547802745835527092561310493903974151757998665341841328220048211450302076898755909821315153920;
R1[425]<=640'd225460087946287989877390137291776354628065524695198707587899933267092066411002410572515103844937795491065757696;
R1[426]<=640'd65759192317667330380905456710101436766519111369432956379804147202901852703209036416983571954773523684894179328;
R1[427]<=640'd0;
R1[428]<=640'd312694321174586587028646462234739719157112810850413784756837656456094047978601863412183616998766690525441399731074891776;
R1[429]<=640'd10047511580080592199131155225536621520295333513968688900326814818082659051731788705910637894995653488405690137528238080;
R1[430]<=640'd0;
R1[431]<=640'd0;
R1[432]<=640'd0;
R1[433]<=640'd0;
R1[434]<=640'd0;
R1[435]<=640'd0;
R1[436]<=640'd0;
R1[437]<=640'd0;
R1[438]<=640'd0;
R1[439]<=640'd0;
R1[440]<=640'd0;
R1[441]<=640'd0;
R1[442]<=640'd0;
R1[443]<=640'd0;
R1[444]<=640'd0;
R1[445]<=640'd0;
R1[446]<=640'd0;
R1[447]<=640'd0;
R1[448]<=640'd0;
R1[449]<=640'd0;
R1[450]<=640'd0;
R1[451]<=640'd0;
R1[452]<=640'd0;
R1[453]<=640'd0;
R1[454]<=640'd0;
R1[455]<=640'd0;
R1[456]<=640'd0;
R1[457]<=640'd0;
R1[458]<=640'd0;
R1[459]<=640'd631873750011343120187508166102022593913370572403294667525865865216;
R1[460]<=640'd0;
R1[461]<=640'd0;
R1[462]<=640'd0;
R1[463]<=640'd0;
R1[464]<=640'd0;
R1[465]<=640'd100433627766186892221372630771322662657637687111424552206336;
R1[466]<=640'd27605871823058775274685614514467385938507091648240943104;
R1[467]<=640'd0;
R1[468]<=640'd0;
R1[469]<=640'd1779227322945296964554040898521508962181356120855162126336;
R1[470]<=640'd0;
R1[471]<=640'd0;
R1[472]<=640'd0;
R1[473]<=640'd0;
R1[474]<=640'd0;
R1[475]<=640'd0;
R1[476]<=640'd0;
R1[477]<=640'd0;
R1[478]<=640'd0;
R1[479]<=640'd0;
R2[0]<=640'd0;
R2[1]<=640'd0;
R2[2]<=640'd0;
R2[3]<=640'd0;
R2[4]<=640'd0;
R2[5]<=640'd0;
R2[6]<=640'd0;
R2[7]<=640'd14821387422376473014217086081112052205218558037201992197050570753012880593911808;
R2[8]<=640'd3794275180128377934137907385222178947880172326887168553606313780073994781116596224;
R2[9]<=640'd28948022309329048855892746252171976963317496166410141009864396001978282409984;
R2[10]<=640'd28948022309329048855892746252171976963317496166410141009864396001978282409984;
R2[11]<=640'd347828580560531852659086279186253910699861789874521850571651955268864337510400;
R2[12]<=640'd15914343595566951398623233717023127597849709749739248070971503263887560116094557193502720;
R2[13]<=640'd30019120336939001004172732863072349025982433454374078734656876113325894370590720;
R2[14]<=640'd101332212859169899677199322521598138261699948794773101008393352639327164694528;
R2[15]<=640'd12531845824705989301507139832157345171965852207559732271451986519880428375380915001172756004864;
R2[16]<=640'd50074418494611761683416531670151311694241871660940519671752224573198917638899217073402196000768;
R2[17]<=640'd12222215869445409104896766487942495384689010216236642810894515026923018923067336961260781568;
R2[18]<=640'd4074083623837049771383660292823318476734199900934968021979160711667853922178893185453916160;
R2[19]<=640'd123860296646158730849283846191605178579924570363680991023859915468852100878977441202176;
R2[20]<=640'd75093294349619196605188622330840954020811571517867144687785046090051840739007905053460576337920;
R2[21]<=640'd17917957945766133338818838600953564257534526749625761840576654342243291175942685439373039251770977550336;
R2[22]<=640'd50079574916004353658137413147470832004207791098880647605326140298236059198177788658587703181312;
R2[23]<=640'd1318041150745077065276524953423627497715731577628719446433852999487804331748996450906283745654530172989337841177050888117413066359136219796454407814485662236672;
R2[24]<=640'd9394743721477722862853975531906411869022490635090759450824975568212742734438706692683119879104719177906126848;
R2[25]<=640'd9404204879452915907458145123068448449362212115272992385798825107819213487223675695362995731476674868655685632;
R2[26]<=640'd21088658411921233044424399254778039963451705242040243681738122304922341450928111769045686392054615247728349493604512040022465536211201709763799982605530956824576;
R2[27]<=640'd50437041368511615697915021551010812245921995037212893506249780680367187327081958552987147078193624927195854073857411427244602682892551544729529701728433503079497728;
R2[28]<=640'd871664547692744299169541835864158985156003816670996352358609556791047219713160491014883026461528714787728993251610533679549661678044242802508428631184999408730112;
R2[29]<=640'd924951194029166771482584704364471680051987223379039927820531011645006535290622063026300158989692382902260711333646902939288922234941929238535402165896937391234482176;
R2[30]<=640'd25049277061110573417941901390308981307605351623826361723378217471807248648170541523923376376781129089389761655822315072083811828659074538680727066782344747714707718144;
R2[31]<=640'd25287267963587666565442167951347366502949603199806303469244615029493715557750925047584255075177447892121116566399851902521301916751389879528945348799797315308017942528;
R2[32]<=640'd1395833526563721953865028027627768931288569993180928831919106393248852199571625813793090183920961559972127984026816609662101328491677117333824122864567761409641599968739328;
R2[33]<=640'd248521086618135689101309743846381524125560890237268543077811474452350596834851678246399286120733962357391996934869265880056869814900613100356008631818799957471229170707070976;
R2[34]<=640'd247570048087080660573282408649346543963228478836268384312830081652123098784942063525429952820048100605709000642326553407719874085201644508428633072282276763336203869043556352;
R2[35]<=640'd12559732207764928253728604805732418590106442500093301390526151736197937104476846044087128551152680845576808222142521057415949801356546523789195827507550372759316701684695040;
R2[36]<=640'd31670851120765145727361874192567798546397376701459596614377642977456622294420198795957665100614945908102881475633784723943298748071605463314081662762777687803773520611198894080;
R2[37]<=640'd138157216447866985779924977152246490791844374692335858694206462606169880242060774005452258532382451943470027804629634714843146270755756056582195484960289378788839589614190592;
R2[38]<=640'd3709956022096568010904841296447712983903289457261282529911452066766188923238486108184588649884179222601318647197235661862421583504596284337915076065409696981285126610414993408;
R2[39]<=640'd531138090995342870943036450103599460841834921578707263018504401760911194677957874260608725001656762866663189378193666470974507066514449892234474813417536698077797674223083081254830080;
R2[40]<=640'd1087783059355290978147379546044834761545939656988062289545451026108080786999676050409484130971577284812185217289576942809494716357137179366334684283351352711152288443202124019903903301632;
R2[41]<=640'd785274024677106895642095504237378258341496046839431756560654650014436080126167533802862057100380631053359240838080895308933227659202072788083121161212610215395792822073789775872;
R2[42]<=640'd506285331815444981221848660527217785759926371745982435339083934493652027384282538220852869150822338538316456132898709241086143744360246459099231241914369268236407037002355081216;
R2[43]<=640'd3643489439326291790842254609805971943265546264348788434291215168800604668961433052587578856882532245712577553373555272240447134206633585775459038506058980029169170200666682681196544;
R2[44]<=640'd3893985669938252062938731563094670617333270203204531252949696035073545087590761101000334428028415346661717837596985063656682672338574748786652625337155006433303960769694080679542784;
R2[45]<=640'd117325627885993651613212459838673748514722626242479280198242283653916641766661940538065950406432691684074195517259933895469308051745161732426760807379368976588650872405605142757376;
R2[46]<=640'd12570114545575039216118641790205060439883406451656899114378056951251551150891107823541919144681476083513789429946311458012604443042882731641234682246237665181725142721755470678720512;
R2[47]<=640'd32701748672724231616401495566394209461592227625316024307282333385458932527316062706557631182231705843647996640300819756782975543819356155339725936165953582812169160446659464483569664;
R2[48]<=640'd51039040737437220064325488089537537585096920678110608340154833840991047783173382066464481219381219864123182374264028450081411534170594928300636581596214338704988687618677866861206503424;
R2[49]<=640'd54306784754463664236072095038103490039756667468487398018892948066319939083475399971754022132804286818596757780007585475654327528640071364328280984613942646693609528561981917542658080768;
R2[50]<=640'd4102314765968388886494568504753028811889999007334340105759077545158984945536966063872776336205475361089251648171738849452552127926087480387370314333346685687306194198020505310038851584;
R2[51]<=640'd276054303561499708426835143896798916498261133936415872047604042862132814525447115506242095986384368228381535551595730393200718590964466069816972702741595297015920534430657174384845783040;
R2[52]<=640'd1671088258291787703334576566284977402617985586806063759791015517143461213419318365991431625641039581519268629832012700044682658399908731675428551983552055193097910667121953144852205401014272;
R2[53]<=640'd1670815722258232635935837511763142121681700002904784546549739858415759513991204888455347159698302577239787411679579791009545796546529073649972912718744787315244391242875713564491362747809792;
R2[54]<=640'd15004647790541008321062781079198075673823560383839603443708241755243189115842646148024563587073890015562783648942061777351878585840585840810235110596149354775967069814642864042241163264;
R2[55]<=640'd8980649227544544340060424063254504837078701761946874811416292965132364858513122451951353790821920244889537297190774271164997362143988470692456531539518574291483894976054775549203334116147200;
R2[56]<=640'd235642544892315650962140610786140475671530392478369298687184739777181757133198197961215639002138877317548682576528636294981247659459639101241371346433272385985171225407194392891661523877888;
R2[57]<=640'd8705418094515914843409686903920779860510447398685768191681014631926500164320699069945704997994333653900532966408946620365754883284474535187411690231562383379801378821593461782178745548800;
R2[58]<=640'd19492850447122437940273762229963585941972273230866283075561600181881578270463481511951202455317003191761321048319318544381240395502214310281614304096905868320507502996938201818663156992442368;
R2[59]<=640'd3383239585292981673546871465775247824633214235195379768708410191448896348697237616955118524550817762575262473022012981283581851759058376238879750784027809940082324527151920589260800942669824;
R2[60]<=640'd15844739687371429126931962523914242267790675825260969255312240207913774842214855050997047230709473020096655393616439722344635722202964020857857178689507176775432586874331553533064470727753728;
R2[61]<=640'd13610185929545502451116207994426836109591944939411067412404107869222537236789102453317553084809946734140141140322048891411790140171675184640965178179070951646478854321620205391223517769367552;
R2[62]<=640'd67321052301078788330841290810408232333743486935419861747681175083128513291785877508487837095761578592662898411840325874549332363255174975291678088438401016429092651779816103894612783226945536;
R2[63]<=640'd2334775081149757950832451885721639836246591457993193745350101552014955543709000706758097610350095785681649793833542255211476101063448057710490539070240721892593045891238464480769149083724021760;
R2[64]<=640'd242836771659631907716062915475100844589783490868561934500917854196581302502604830083529569887823499510744562939631994267743936884388879618133007122589326479858911808781983696601146507132928;
R2[65]<=640'd138958927576499865622748012390395240331170987275979938918910544040186395066467465025024003879699808864785475059823461273690600781112655093185643566534523738401679337930374694516312908021760;
R2[66]<=640'd855527029166166841153813220972342552437448794974474497331256854949324084433664299746594904916846821602709371668941857407285490135353027164045776790315378104581475412832644355178004281600048128;
R2[67]<=640'd904787197107448951412529234803651677032433920930586155009826921413591805471582272215835991982835131774146804572919563876467151631403910029171050670689262821866897400307750367736399767075840;
R2[68]<=640'd3441357883244777074922441889706995227765913449148747472893273872027880317868974785214653584499133554506483769967697419288634102286659679764035559378770540822342652038190724004708970426968895616;
R2[69]<=640'd4013333810096242416134913786793626652219062656148695148240824691478708347448317844185787319632614765437381626674444679817256250402712286680152156534212740610802312125724107001270973393774985344;
R2[70]<=640'd2003968516900798884928243031712812277293236722394539874000138125141250035142894330546813467507480763178159671844751171503034997707054447875074197623521050766061736719309153174264730536666488832;
R2[71]<=640'd1006108670844325936559248557712691010472897328869989241190278547214712706918312032995933879026719578689493552560182551281685755952534334235179651434427488719507949994236622551054118947250108464;
R2[72]<=640'd1994394948976782028911121324678987628489138409078591211678151679128717755887482725574400078669662894197149322793584858920710407911192868581693428933078110589546591734008768783070829350104135616;
R2[73]<=640'd1825086695707297954287693265816822137461432435265394578884416241268628847889696413775835640675486863488894391466525862344889358075354386943863158313732661410711830572353122663408431506344705984;
R2[74]<=640'd4355789358677226578555941376422409883750802072127045291763835227769556469668202092060046627842515263586176364206474805073911973415649149528828070218140021810227792323094686665450530703898639552;
R2[75]<=640'd4278305282636371120817482758301920011854345722509008682835389160659394507769322383678210187855372808197321855808267321466286449680378261912227483615408492531168712424059143201461475492112399552;
R2[76]<=640'd4421594343372528765380597587869953181074884445961260799323177974790773986287599873338336413629631730572917588941177050900518816779028932400886693892660694627329328986922645629745367128944409792;
R2[77]<=640'd3869181463161192158057005108344269109556765295662482236146658527397064907318681714647401877500718024419609482046674736303024233724805379378412111683564777819159880786935209651390503173512232704;
R2[78]<=640'd4555757253020230585294582253580068130698802994770516444278253895407104575191755767839271408446959387406650479221203586697492982281773764614032200377616290403441208984663891680840053099295014656;
R2[79]<=640'd4559934292159899343124148755904622840774083660518119495972509747932036772915640665348889858896280462377224308723835614766232826154117228807964846663917937440277915139148419913385044457373171456;
R2[80]<=640'd4544614496321615800728763014044686934106808404843486216112686604204143533280971801346013968768551608934182210399665187391883740567746874428568030035733910040471448992973850684909211426471541760;
R2[81]<=640'd1140610154405548804660292901425072831223307126812139982644798129474818791802169346626478202759352962738640116723560925581614462041157040415502724017075841183552324913935817334918319845410864128;
R2[82]<=640'd4562440481650869057548794341165710447461259910872721792459020178841575787905366062127738669951786906993022160234966065984913313007055446651026659390433902503869129516712261819951743225779179264;
R2[83]<=640'd4535707431156989007439568726288560302979463650088062261615782722682009722472502718066180586932990137561331414792468143719049478995225793866840051771764336344872848536657123056205008055333542976;
R2[84]<=640'd4562440617622195218641171605693093062821959188449150075458028071100727600094447306352823724569659604554503640040402123140661574150980601271194199189050490940223729324950703281789086508091702336;
R2[85]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811177387486891719291470634414464017572935779757090119712679271017068115491614333067153812407297901591616;
R2[86]<=640'd4562440617622195218641171605700291324893225233857952034437322504709578339609525169863866768112597886788560168412067878811713133518306163850558995413138533029206554619435267639639274588634869696;
R2[87]<=640'd4553529600790901868604763067372816415801859488534417886604829374013569507874967988747207556611426799611581389632979753155672450192495012673155992891521530488008970006533951111598996859134134209;
R2[88]<=640'd3974313506756834116238208069365570115815337876196240497788368124291374156440793684578837193580848181086523974826834255306699835451525247920524357787125749698083939266194578309751657426797432768;
R2[89]<=640'd4562440617622195218641171605694892628339775034893883336299034333073783116867138978225168882957858615242523689553848447503397319795470218046611402118435890108347858702673043100090147263041503168;
R2[90]<=640'd4562440617622195218641171590943945462977986210134695776006999352744086427103649687690906262773776508276121403186005079942418876134357052526212753028545268942792368062823246117941602532856953824;
R2[91]<=640'd4562440617622195218641171576216976102230560010823538498022322036827076395198240685067237933607556671358947766231426224393441333374380127944325127108124853261374965667060047669438632976453728736;
R2[92]<=640'd4562440617622195218641171576216526210851115511357081132597163478210279908283867143327864228573313406246093324790880873874612415786096888507597003621492560206057799247009647176542943312921754081;
R2[93]<=640'd4562440617622195218641167772769816967054099386211210387195967103436160458192789870821971100654556947067513560628106179324335990322575116719243281444137363067012081867814562911387054664629352929;
R2[94]<=640'd4562440617622195218641171546732255847700850385135951795581314008646626953678391595736994846530680798116128155690008948202925072508353285644483880370019661667959813333046871736192052547905650625;
R2[95]<=640'd4562440617622195218641170662209819559699453208682567388038034870658171992891300890781920600704950302547408061702673036896186212711016866518488880446494384344321639372138328484748131319362354785;
R2[96]<=640'd4559098986310460212377516516859446568230507072523673325114981660518978603211793400220299047281537259864350834096810074261079608225401085246433986966817089375166632909171000417442567328746170360;
R2[97]<=640'd4562440617622195218641167831737867045670891423201533337258194837279937335267282399123017120686678350978434495194465829618834274659053546632989031996103204005657421508273940381537570579816642303;
R2[98]<=640'd4562440617622195218641167831737866503351876266070149642623378664859537216958310620483247484719883186219479849359307385430701199404632625607957682482848316892888153756940573212511745136574594247;
R2[99]<=640'd4562440617622195218641167831737866503351876470466635974562970014569615837665854326624416886242992588819746578663713943083683296414404266533988241803728086149939667239828545098440193014486761199;
R2[100]<=640'd4562440617622195218641164057775441681810524024151884948242674652982360723085547272867009788492609071322666359541072148658751417004845168166272003138653637026219269548430550360337745679745023998;
R2[101]<=640'd4562440617622195218641164057775441681810524024151884948242674652982360723246865242796315210014747286119334495802525461604506023044198732180007429995286167760039884576427636921745057963319491580;
R2[102]<=640'd4562440617622195218641164057775441681810524024141153937600963429686986482759354469532771881944000375878607951265147790025797048717215161526948033421930733360697537070687730749773557203854162431;
R2[103]<=640'd4562440617622195218641164057775441681810524024139751589619376167551795530727542413760079771597862997122996459659470416585563209356863139058851702873933901376949014984441617713456905791964446719;
R2[104]<=640'd4562440617622195218641133866076043109479706091752710219025613896233830392845115407367820290852566872245416558688938790442997084211153836626891974055531659653231496132786411520566545586761760752;
R2[105]<=640'd4562440617622195218641133866076043109479706091702762242220558020531724837161322534858728169091829480811675128077971912956752659947194940510733670248263920129501557780184522023307418735986343920;
R2[106]<=640'd4562440617622195218641111222301494180231592642375282409772349854926729254414760850804967396875116170732136598962503203404374162275790536057345609794413518730028812896712176587432214960038477774;
R2[107]<=640'd4562440617622195218640903654368128995457219356873358540809036103871240937392929289759974721413272782905300324242493653876405575487385934498767518484085573429380826439308690965160528860541878222;
R2[108]<=640'd4562440617622195218640786661532959527675299868681305605390277411352265039450834925740137053486741662518901978655936595715396171959898583421957559964030540057571067217344282187807727285333655502;
R2[109]<=640'd4562440617622195218640909315311766227769247719205182603463198901825911826752639579348964167182685667598576937672760774051593671886084847797494077734539665819542402112577247764343786485791588303;
R2[110]<=640'd4562440617622195218641135753057255520250382212480040966265955404007511085712057861045035081849371498236190988398693833263982878880998064554543910408587966427534245225132329472101144822366076927;
R2[111]<=640'd4562440617622195218641133866076043109479706091702750226704238944995095787619450656590153377964362291699293327724287226866600739043100284991549135739486684137701897421453078888769807835618869247;
R2[112]<=640'd4562440617622195218641158396831804449498495661807526567208644488855762533888684621783014519761387531518141677109155845688614035231640915660396096814943821831273521454762598695137652136787050492;
R2[113]<=640'd4562440617622195218641158396831804449498495661807526471847403861272138494139079005464184140852687092719584631282312704592819341350963242616392340557195082146029076642337330672788657682625069052;
R2[114]<=640'd4562440617622195218641167831737866503351876265693978942356819279332973591513754622744089435602842056639268642235899374395947784122364561954649288584345895796477932349320146933176764779741577214;
R2[115]<=640'd4562440617622195218146507028791657435230871223654684562426109616195306434908141150950301042926748168793064888338819114110555311742481617674517502430102217002473900272816876561680254021597659135;
R2[116]<=640'd4562440617622195218641141414000892752562410574811912024800206609368862563608993456595201623703046993084395747081480056242619971519661690627994526458978921726824335158482352952295468724635303923;
R2[117]<=640'd4562440617622195218641156509850592038727819541030235977875770277053744227431497824458651917288171324111135994557576318937162172989083452511266761103049134696804887953447826388123058520167809019;
R2[118]<=640'd4562440617622195218641167831737866503351876265693978942496372314397730114708528250773833779774367458903196586342529067630969011658776165746234305528170859590870735199981473379208222844026617855;
R2[119]<=640'd4562440617622195218641057443336940473267323200222485035631312994452032933543564666323795968274001329111443643381006050019562156674521555016341828812203804488872673479073574486273426739708297182;
R2[120]<=640'd4562440617622195218641158396831804449498495661807526471824145022094679073072850890185402871761759462452317818918394221064385973938912244451379943093371110176746070041082857528632994342778174719;
R2[121]<=640'd4562440617622195218641062160789971500194013502165711270804614766361342510611051603614758259608988654503549505536358717480098116130199419048561758600849940510011535786613563313958776695594942463;
R2[122]<=640'd4562440617622195218641122544188768644855649367039007083827893451602111209082834840340462687674399158687002399363199837604039259303133882550495082236773038552729811713417317540273237702217826303;
R2[123]<=640'd4562440617622195218641167831737866503351876265693978943798867308335457661160748612430359770368011980065723431592901649107447721531287078133194525560388543640032523545256407177065962557285597183;
R2[124]<=640'd4562440617622195218641164057775441681810524024139651135251180860573692580433532683917302856089359539645812107982753220345004684489042978203420850396074038932877877250328566660801560925200973819;
R2[125]<=640'd4562440617622195218641167949674192279025043523242559764913063666160969015262319537794555733416309883148521004119818706660250041955241338511586868914024930857128552592943000977585028729350914047;
R2[126]<=640'd4562440617622195218641137993847445258040560105903073027626434106788102422725659389102467937000547727579872495738515834512565247063774533592720881130203193618139230903792656023520032499360071679;
R2[127]<=640'd4562440617622195218641152735888167217186467299875238828236519110307165575661072637036141636769055921377470560122124647233160734058883703185736585118443683897686263448427551524270213151183585278;
R2[128]<=640'd4562440617622195218640985739893623954226523849084642831317081420696791801504266060266129500448367701909907310222708888175039676533791420037879330334048352332413190929759536487914930729715236863;
R2[129]<=640'd4562440617622195092006979887500195753687629814988911791156153287117507968927153343744416574087632353321566354580128380991119262804919844797253929005278256101520395249773289007784842259943391231;
R2[130]<=640'd4562440617622195091015726020217289349252845008561643328289673426265000309563666607094979340912456697766398266470172739160627680731955121549674167312322383238133274398001603429300427208332935167;
R2[131]<=640'd4562440617622195217651608488325745692943393824467146794254304149607575271592183974131047124231208164170575760685948562069274742347711331559618283611227517293997824551220982991063587477593784319;
R2[132]<=640'd4562440617622195217776964424228618011357549008945579348154255883105020750014964178822751242782166759923649799772172054954813025403518712931645678017374315773670025409975576307321048763568488447;
R2[133]<=640'd4562440617622195217652333066999150128703213981432899812655960087199435652617973312947871190000140549828741707042188408394833780474237403103832089820700009699290083681142985205768627356574941183;
R2[134]<=640'd4562440617622195218146510979658570920281974351532136581061041988943509461124875925524281241365240213421231036716211520813069080456502326736385909957142383320219629453084249827666342323622510591;
R2[135]<=640'd4562440617622195216167869684339028502486948305664257984237704115204295572796630797655632235802333840230571228544798786024131400559048568458510596647829220177513875984620203889780778427188510719;
R2[136]<=640'd4562440617622195183041051958407348175518792795176665097092228863615971392604344375248759864298908293997367608549084405517438570272674792105388882288709695817685036192156093640003682524452618239;
R2[137]<=640'd4562440604076101640195548869803415575935643853963897759882128700939113955783943291758267333892884484680305626986997262662012426702654238191921660415083724139211463394384648202420127361893662719;
R2[138]<=640'd4562431900718241598294188828720999438596537264222620960475536313527013441864238912797062669566176594041403447239501393335041458712397448192136912906937508119906356711793288182552327397536956415;
R2[139]<=640'd4562370930458554658340442133847713642813671743444454063310491725408594848402845451005359819683004332295805137343432143253756933323426377373371921663606328841298158710882974554528465949214900223;
R2[140]<=640'd4562440532670200298514004359904629875759225927332555532930603445850849284780711751674707663928784751766915783911713783542098239936278511311788609514383182484223541844978206296135551573540470783;
R2[141]<=640'd4562404585234248249908654711052693795367333706869458632390776361870831789869203640218154745828457940095439728373469321630501384006956771531716543529454052204117322285948013144120925562509197311;
R2[142]<=640'd4562398874433362598230069217245341013029669971169540905799276263782546412814576976245140007009766799818871267111854536740885497959420031252652452042267006303279307627127080891158805844504608767;
R2[143]<=640'd4562294329475811101410436104516224286578207455203097513244764019494447890490808396327968504121484776903847112760839534057164646227578547025495528695895375027247659956051635784726619259809038335;
R2[144]<=640'd4562438102158885463925964866815445392635182958953014492381964588737262803191891816463242839119333765048268852259550144423417377283564668328696818519127465087262554274713577317980486671093727231;
R2[145]<=640'd4562440579386224632798160075571494856114656112880809792594949139672062758626342576705791037952364683008685651806541009388620170521224562312124731557379877528585662112893390971474002174250319871;
R2[146]<=640'd4562440613912528300061552682097209283843295063934698108045768593890848311542955555696056740029605017138896899821151152627038057249288512834067936752254988002935140379916846876527632716335677439;
R2[147]<=640'd4562440617198944630615299179870617466804870850704016720282988800266063881094988932448594421646795914209886048466632904688096345643544131338986704382051275462952558316067177378874225427147128831;
R2[148]<=640'd4562440617489410720436979108207210124695738588331305990674550430866343998365741292852534816313772418317926000243527887361485115485871897321452621337626127649694414033359489566061458024824831999;
R2[149]<=640'd4562440617622195218641170175715143032784806395259522616380636909654799902367934383540538395121575376420421793964173756971628538813309659462088440465708151865044887120029640196177528674456698879;
R2[150]<=640'd4562440617622195218641170662202486857436621332647417821899682153935705936313295256232547029269411200009660048452875479876577072422908973417646060639178295802285261081496334621152179864905711615;
R2[151]<=640'd4562440617622195218641171605696692193857593950142311499773045150979328107843162042439488097957786103257497381595892349347937161528892273250929373999309681335064565190841625738109602864889331711;
R2[152]<=640'd4562440617622195218641171605698491814293792509740313435031325224543865641317655365364415567451976615268581026372546264988891036028623442241458980180967935049691188236937973942439844653343703039;
R2[153]<=640'd4562440617622195218641171605699504014979183447881568086340347821522950358218045878622160092651154758873920003251979609483131330119455859546457530889733848371018019568084167896374338352584851455;
R2[154]<=640'd4562440617622195218641171605699392036399751397375897301574832621545255609565275212959844410961994862362342462847874602548231871100571113925371821555568656759926012037115366803238405396007747583;
R2[155]<=640'd4562440617622195218641171605698718417832154591101700130086821812526093239323765613087213268890692187166605253376174793157674556654592279027002642579514189085682017224512408727590840051890651135;
R2[156]<=640'd4562440617622195218641171605700235925118011545711833812267352695519397631835805729200016929119192360147133716092257746919224669829313825310842589152644604085314329688767310608911914541871267839;
R2[157]<=640'd4562440617622195218641171605239547152556788236112034669080109419471516147584719375477935913625036354417326856006215233480507421603683402315833401938492919744091261176389911253863694944912277503;
R2[158]<=640'd4562440617622195218641171605700180564386331276167950447914663440987449078148838385222100140602327743363696893905572599027414929745795552839574674680177451427217575404531261054652202311133167615;
R2[159]<=640'd4562440617622195218641171605700264932749574281361347575475841881154025055595866052000691032677252053858011144785079221916204278288437221148468368710710818940210762486986432825511964554871963647;
R2[160]<=640'd4562440617622195218641171605700278032821496615915958520077745682586800971922815601847971781038935000820542519183025174358824225781108248840043733875714814825800899677992096712123793820056813567;
R2[161]<=640'd4562440617622195218641171605700200707740652904728128963946578121302702527010617400130898852375089343175568961884485513251103659471980285289104220778077488664536153801298257887904767515335589887;
R2[162]<=640'd4562440617622195218641171605700228896316044816044271108376734686152995212382576222373899017651883320843916571895692900010296377762210493224317763607654639176208206486564166982712033039548940287;
R2[163]<=640'd4562440617622195218641171605700278103185672632254708098641683740229433203621657121062799799719528632634682362053034452569539043669492439459924348165268829377415304506443211330100332951010017279;
R2[164]<=640'd4562440617622195218641171605700224544034328293237711809851644701101895786527034854336961618353536310029483631504652343221800144606481670641960606917844276805632122851149404773583995550023286783;
R2[165]<=640'd4562440617622195218641171605700234206250442735000828243976576312616832540737856512341027148809206709202088733328515868033699906056279336916523132274328671909482340928827074868688595515036663807;
R2[166]<=640'd4562440617622195218641171605700291324799373851738961750882175063804435768646510904279524443388429807021899016990049256788621482021870429282871713573051722783949315877267353171659087860394360831;
R2[167]<=640'd4562440617622195218641171605700291324799373851738961750882174360929935863667084834966436393381120304789271164958613938525240850682773683318270250958999667668471089838744015732563181554074910719;
R2[168]<=640'd4562440617622195218641171605700291324889876555266074281304299033826898592345493394092875646550171525776910842586604019639897947312350422392032446874754598972418189067505741045869194683476869119;
R2[169]<=640'd4562440617622195218641171605700291324876468747339253432755040981655367860618303655030525080705263242367342741963316192837196847005897213305184487444749645168224795398910366560891620941937770495;
R2[170]<=640'd4562440617622195218641171605700291324889929134102713613083086176143779142979812472810259382583540739197504383427769234556991475368050758761823269093012325901383403907781837724297637466172555263;
R2[171]<=640'd4562440617622195218641171605700291324889876555266074281304299099851204902438201168661019202538420650148695282354756456819016712295907281994849660239007301273908614914534209275962105078908715007;
R2[172]<=640'd4562440617622195218641171605700291324890722010684019956696663400159759696570655944101595813728518485511958545664083523705022899621864726062886753787774734289295267158080699266935242722061058047;
R2[173]<=640'd4562440617622195218641171605700291324892850123753161350884025797206851413614255171962367838193346974391089880699175682840593181433003583002330919011541289109811503836811215948411390615256825855;
R2[174]<=640'd4562440617622195218641171605700291324893039366647808387053770127749719088759517206125636108912823397992822610138670215557046057765679151314713114371722294993208980412111788413556798316863291391;
R2[175]<=640'd4562440617622195218641171605700291324892397072517837037431267785063820854587827143706482063047422136866974809451488477602399345784913481711878662790127014027332739838377821113408776363663425535;
R2[176]<=640'd4562440617622195218641171605700291324892861887540277856706280119053909773811364936761664828086050424795283025962454293756558913891331776674806904816903170476635796302656157134741789821517168639;
R2[177]<=640'd4562440617622195218641171605700291324892809513272981774947484192118151821913330290274591867680137000198029703838851052753727488800629652267989892766010565579147164934067693538555947060746518527;
R2[178]<=640'd4562440617622195218641171605700291324893019010253519418050940570249073294893137359035700790160876796549261978741751161487420142110112143147067265167141695138277654236880597134994345700236460031;
R2[179]<=640'd4562440617622195218641171605700291324893176133001918329161840919531219829488236871557825420618646229089900278798043744063505608615716104060127465566344769421486887101995415479437591359361384447;
R2[180]<=640'd4562440617622195218641171605700291324879768325070646934112280516576241823397137746045419028168889777835590820743607814936822551544693769696810781722216444876653411087588602812706348277742698495;
R2[181]<=640'd4562440617622195218641171605700291324879768325072402890877649864333599580617830608562833059170025745481587893226637634539018259301487249081769740341691790359514970972944752091944972281232490495;
R2[182]<=640'd4562440617622195218641171605700291324893149945874750788860737290595525454885815903747628284336889603031079009540677516512912505447909015643406821553365421740887637175943758635100646273806499839;
R2[183]<=640'd4562440617622195218641171605700291324893045197376075548696080691586901136780844757676211306448114723041420931150014871616959068743693388511282241061637254834710914984923955385366707572054163455;
R2[184]<=640'd4562440617622195218641171605700291324893181043089232947086025167054831679252676188326257126716996907912758079653477080459354848523453277120954972145564038978537921282882391826542524842901503999;
R2[185]<=640'd4562440617622195218641171605700291324892704764752857422108630741944525938715167633046552179036280884963849221090122664535777488133375793081278766529694839827382073963148498927568512536251727871;
R2[186]<=640'd4562440617622195218641171605700291324893176133001955340766552953432888153732834973553422299930830357909933012520279011129872628675519698741777023321064364547077804311141980768462164109429833727;
R2[187]<=640'd4562440617622195218641171605700291324893177360532798547517219907786540713813331507704852539582150697531688674353121141955529765398213591677110268629438403273629179093620762279672355401777545215;
R2[188]<=640'd4562440617622195218641171605700291324893020237783619532748163032110851758891334953498772332404522930450519224410016122700410848126067034721315123706534892598254827740581596978769544453579341823;
R2[189]<=640'd4562440617622195218641171605700291324893058700123262312409683725671167993609036945224757396980093862134548266255561631533246101294583445065094040419281262672423712556696754657638187095056973823;
R2[190]<=640'd4562440617622195218641171605700291324893222577449727622744931909947907497072672311152319116905834404409164760309864958353367229911010198654710336205157050023925792798450160320577561275077230591;
R2[191]<=640'd4562440617622195218641171605700291324893188469275014847011602105502731406613749751457562714879752545259193255721089679841533373627083807352600948737437733047491728653459830173947080698566279167;
R2[192]<=640'd4562440617622195218641171605700291324893228482674155342491327176284412115552151120853685075978997955248504441853588016144419962203522511632137378230240640137859758066403318084511081328917086207;
R2[193]<=640'd4562440617622195218641171605700291324893228507248559930579120116865148185225120770431918426504807202645270132101129477670928962753390897767519689704130729887969853840366033135915897422279081983;
R2[194]<=640'd4562440617622195218641171605700291324893228507248559930579124375685798354796745082876105270421086120548607573468548075709056850647705643322521188157476161220074861014646598665667854520725536767;
R2[195]<=640'd4562440617622195218641171605700291324893228507248559930579192240553793459825911183064173319765803436660263960950470167482220502250796641646011449345696991735344414403104404927283146317740638207;
R2[196]<=640'd4562440617622195218641171605700291324893228507248559930393121804414615357272093893415214568124513990023721182269177995642862528068604270781263773095871268727021293863742406252294743780656939007;
R2[197]<=640'd4562440617622195218641171605700291324893228507248559930579192517185800104317237234651506427034567695080977362649659573727002590731732303912264902870579651304307619010858180656162715407730343935;
R2[198]<=640'd4562414502645962466111987207861401184570524610418197312802562395186547795114571027187580723140393464437211346910894971870310784217689699452495357781358736956473935866645596374660784867199942655;
R2[199]<=640'd4526666013591206781012459385105529174144052741519419095451675078674258994844238770025665271145442244844941429312788327614223161521813740656626932242887165226352934719670916976981942021008654335;
R2[200]<=640'd4495330032005027655210818368360412830384817167953195322304753782398598670415395055102549325225054510751216710837744167014470908256140177094465694227640910988487452513454752481568119157436710911;
R2[201]<=640'd4419864450301033613812851766093048436062174017652319107334681029607122891517865273593728451535474682513051945045402325671460876067935049269314185756914219194621527576803686578625386407266353151;
R2[202]<=640'd3421830463216881382066894978625353050093432902600955553313273474376143230681077019144578083062304658955769394447641470242118080501213648508336712418445485161046673508123639983530428643904847871;
R2[203]<=640'd4115825210913932551300822452287948889374527745036556051867276982387210395036761822708294861205231803214415454631272966735942945985260687084924893435617098280676942453808937566207;
R2[204]<=640'd4052323130335712962180788430016154473333100806511529918922975614535800566195870595047918488005347813700091087396903893644550627797109424691556177618347284343564521153394812911615;
R2[205]<=640'd123665200736552267030251260509823595017565674550469171750257380631364401281280309605379394107853205174865095208798122494380878140982179056143381355257775243822930815904382975;
R2[206]<=640'd123665200736552267030251260509823594972138254282125869652666892573981434716764635153957645919365013565147877029505243543548453315445853675161034707775145575808672910716960767;
R2[207]<=640'd57968062845258875170430278363979786202428266730171072347275570235191685508207585746677234860240441190817497207666759148581004511044720632242225073084465293706149019837792255;
R2[208]<=640'd57968062845258875170430278363979810013892011755071668885136352836352749921228872362648732566474008424050363224228995493098238370571992809209156736026419984606542165799075839;
R2[209]<=640'd27051762661120808412841276111648523930515110001274924927775908728487603327053326950251037915154136983523851529926772392722120333887470338246860194287584171625988670258937855;
R2[210]<=640'd3864537523017258344695351890931962038727329674115162696542623707394896682034558052120870231133554131979577523305769810594993180036333963431593983668287456849995150737276927;
R2[211]<=640'd3864537523016791531698184794773582898787919078251155977852512103762164404776977176304390389702026758038186379705116895534156987947165019707895211157491396819279530302636031;
R2[212]<=640'd1479393270529290811576678243171012679619177855926561107246834283908314320500406499931817337582571575936448705759578523060119322014538973272908463880374075373681115421212671;
R2[213]<=640'd513258889772269785629237742535339486707045356261739359510886048296288332595377605024438048991576512131756343773780279061165469362843268149984139043366350822429238027616255;
R2[214]<=640'd1879602993787719886427217732917653713265041044110570468845082813898353258972030164654748177630220086344513962287062493520824379442874316302208394161542800746472854781951;
R2[215]<=640'd885947699207660042319079326171589467035999453975098485078714454600786391482715183930953985906965346328603244968292204197899703252842502077651790562088269872900022992895;
R2[216]<=640'd99588373653143831025892574942399302000024775927499371320283687851007379003587315179422889169375466522529711663703860519574273337628366667500806322287381525992425117044000487404208127;
R2[217]<=640'd119306677127924018246603820627732928280704691328604486652142892908678800120584259116650177060975062623001413870914546489300194097082115509076832656589339562778419600281198912751009791;
R2[218]<=640'd1178588041662431795902791298760727366459881035729573011397810016024783814717263649172694577872937550051538222496599898618570419531173385602708526476470895977466077493684613587247562751;
R2[219]<=640'd4245472609878703703759921539629857022315258030606532853855735745086527716002016792585434641640729493697124984542422946930698078313932436767542572790960294944823937562434973743548727295;
R2[220]<=640'd1062227105231630264783900967870703866372247204775386489467663683977514068775049714543501957358806229008918361827710626084704189308690576961087919426058732743778403468628316266180902911;
R2[221]<=640'd9560467408390285726574800650896637041567521567228644422416624498166018536882745982377351949555958607650229527575612431094384156532943634684544409845111851813702858591929434698615357439;
R2[222]<=640'd9560483744068642222183066278967145284287556484663270482371845392342721470361182664745583581300490727103265801783903411510674343200231334593724944148461564241795489794758243370026008575;
R2[223]<=640'd281749584221490225656496603639929229282425011470376194077272943228753053414955196100111019243158148398707539271067099881725568857953612876138811169573624440918663409420424384056987700166655;
R2[224]<=640'd3263311827661180151527626282322210656387732594775760247732480169814521198284064379778330491772655106832745508338782006418782236757726932569674775896793180406797127208747360147879506214909;
R2[225]<=640'd8702164874246348231751625310902096842266004313000662272980681317417497719344328558186549691413096695997402752239210418264791318010408734182428112886900866692476970588418953837813274734077;
R2[226]<=640'd278469275977916955799381059847165403790426287854632618940018553516104512493902628869740697136892910645495341717401317347568268958326969243567457333057876529460888291830153997618927345856381;
R2[227]<=640'd2227754207823337508981367775501556050211291985463336299093779867577179359030573461088935512101692544726173447240714305394509062068683028957702766507437424577634963436447666319769723999345532;
R2[228]<=640'd4455508415646675018083502348597401423694313717518297202696901214207684811769185410445336424309807666409236265363510195530931271733079596896170428262457309896344026284567051781873487619871613;
R2[229]<=640'd432184316317727476765693340382999713132434486272070790694496199767264731737582690849198407625732786684136526624893137204087498006046485987684011431834392078494723422192354440141561528228296057;
R2[230]<=640'd1109421595496022079532861130420518585223868701786080035859908972161381507243614744966823922514682539621767645630996975080469252154906000283537134189744130350103662885928266910609336448133699005;
R2[231]<=640'd4562440617622195218641171133954988222200559477054237307045581153284122615153624035780708519182427620674382000847699856272392929990836632350980613396558290627001977324261507555461662562037864892;
R2[232]<=640'd4553529600790901868604762831535256392052961905223178775197974350205176869370203555253569113731514536932993301469657725614049186856562850082451268776734789812704327150205760001352142860008880624;
R2[233]<=640'd4562440617622195218641171487763965549220061249699979274695789676745487029194918927405148082711923085262831330946140996508959957313441759427823993766094923371787616667286669386675296872416672052;
R2[234]<=640'd4562440617622195218641171590958250602934082600054987396227869798191944829239528118096810301709521687458084074680445482774656224436746036290427894080622953333928599722879517013072031860774908776;
R2[235]<=640'd4562440617622195218641171603857536234648335268849363405473840468241571079741749151736255148371770364062007478324088462910539663751821495882533258104284162734518612094093005296184398205526178742;
R2[236]<=640'd4562440617622195218641171605239827498021732357467901458708396660877963595251684677096967954344673180945102726742552581221149786147080380949811169292521413379936024210864502700029309342978427888;
R2[237]<=640'd4562440617622195218641171605297863485971339590806157262555246827737391695867717123099420910253537362623185757553229792501442663924554702534372526086403494550085615069846355948234909303368841151;
R2[238]<=640'd4562440617622195218641171605320554882422566837561957915036964038463395025932505602048493531544233668413727233129553010586139825943840325145518357771719692540254756243353853133280001761555168445;
R2[239]<=640'd4562440617622195218641171605698709785349096976859983921604388747119086336980990178908667291653943704716273996926552899076807493387583689108492332606905339419967964578534445891001883132137387718;
R2[240]<=640'd4562440617622195218641171605697588461840100602546699539718503213825347976568816518690882427476908045685326084769751688277539725257831381484752648527104739729318286897682228463104217219800446671;
R2[241]<=640'd4562440617622195218641171605700290446306390473970058624669824328002574729571349772539317329398240621757240104380012452497435426074692164071103129889104084715741640352375989027789208067706693627;
R2[242]<=640'd4562440617622195218641171605700291307677603125202268291400187429304869239997967709401246766167150182537378001921715193000419621674806795456892174774600441160359895478287273261135781042282151803;
R2[243]<=640'd4562440617622195218641171605700291324866412891388677767099824647575191991404581472098099045902207892900559642931012562445782502627537666214830108203273940633732179161779906276342168290962143921;
R2[244]<=640'd4562440617622195218641171605700291324889902742401915396269032445316912712822061598369750930451936611211785372218098589634304231993171169254598722351135465479317700178220403200001835150005362647;
R2[245]<=640'd4562440617622195218641171605700291324891633548872909756201007309041270321231005394724264305630720751723976724024242238208124167524142076659015259249916789571019622156150538903213344320948882925;
R2[246]<=640'd4562440617622195218641171605700291324892599811664924780666145773730801299264415337915003749955493872608478324085385666199814054304541296558212323263195793142480476790074305487245021780933992177;
R2[247]<=640'd4562440617622195218641171605700291324893019010249502148371078275700505271310699526966443174402159656086608612237205300534741616567296643310756357503033761916677778739485475153556202983553287063;
R2[248]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251926201250212286846565195916635918;
R2[249]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214181605715253614862809170801460772157135;
R2[250]<=640'd1140610154405548804660292901425072831223307126812139982644798129474818791802169346626478202829342849944660577393398601827672176180343859499563165329930553542742962046778666038278840658715696157;
R2[251]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542336656619550707335712486165144348349650456918044045085964874890791332482638373077871074612033813724391833891476576;
R2[252]<=640'd285152538601387201165073225356268207805826781703034995661199532368704697950542336656619550707335712486165144348349650456918044045085964874890791332482638376069236832980670857836710027193289729;
R2[253]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214140188953990849816233393596340969515972;
R2[254]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214170222817216214621972827107554298389635;
R2[255]<=640'd4544618583959608518568354529115524561905364333392120243350367547126231123586768490464874089398162917748256988051822554157131326968557565193571986861442049170973876590840296590485099384474021173;
R2[256]<=640'd2281220308811097609320585802850145662446614253624279965289596258949637583604338693252956405658685699889321154786797203655344352360687718999126330659861106713190881496479517968866441882729134714;
R2[257]<=640'd2352508443461444409611854109189212714398070949050038714204896142041813758091974277417111293335519628010862440873884616269573863371959210217849028492981766483871260788150005553671625855754000625;
R2[258]<=640'd3493118597866993214272147010614285545621378075862178696849694271516632549894143624043589496164862477955523018267283218097246039552303069717412193822912320049879788893906774577958008782476471736;
R2[259]<=640'd4419864348321501618058634993022157220990315116397042432748592751714922818233406218177603035963703543535559737399419582082229682698832455560807265653480894517981240852245554405786024053989996904;
R2[260]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213962622498739062327112928955572164048080;
R2[261]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722211288722709686634988216749181972222948741;
R2[262]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722212529359878081667405927908724519740437435;
R2[263]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722202554515023087886536257769107524566852931;
R2[264]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722116011581182449933425046269758947528902699;
R2[265]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722125712078677430040314811323142284224480238;
R2[266]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722114825618951828584160893888243940874968191;
R2[267]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721517220512023417128868598522636694050286147;
R2[268]<=640'd1140610154405548804660292901425072831223307126812139982644798129474818791802169346626478202829342849944660577393398601827672176180343859499563165329930507236362162543899061541355554280836013420;
R2[269]<=640'd1140610154405548804660292901425072831223307126812139982644798129474818791802169346626478202829342849944660577393398601827672176180343859499563165329930550824394598677777509638816349688168418645;
R2[270]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722081426890709547950127605291036279578248874;
R2[271]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722154277014279668333912494187060163248651034;
R2[272]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722202599433507129365769153405493255794582460;
R2[273]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721835451146245600721138697291297018651597755;
R2[274]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721865213086238228873015307305560773927631271;
R2[275]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722170099502501670220932064721583215713884489;
R2[276]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319714478717512379962777938614963043945753258303;
R2[277]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721494575861827064671946500046036021850403621;
R2[278]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719182948201419711797000160255695683227556382;
R2[279]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719339048656123586237642565764322384593920979;
R2[280]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722189102548537403907679091300985866606558280;
R2[281]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720785426738045058934857267955981476232892175;
R2[282]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319709810624023325821214416859459408186099661289;
R2[283]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722038555952182663531723024957589008728118368;
R2[284]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319693553713660398313698826367770402983397086880;
R2[285]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319699529061565720733777949501494039269860340212;
R2[286]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319711056228207186011707078327801272511956673469;
R2[287]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319331947401421150192404911269300961136282252595;
R2[288]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319542317513304727948596126776204231045447714417;
R2[289]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319443437688304376223756102587288527956481242245;
R2[290]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661316861074342173258118062450320503233374491738107;
R2[291]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719055574376270873564984188417955115470358781;
R2[292]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661318974956815980080285016091108257692791421844084;
R2[293]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319709448408607430441824799664305004973684981340;
R2[294]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319519345898416896271879875280888988734517201615;
R2[295]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319704428030666309393636420842002802578164301023;
R2[296]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319612583214975755697489469736333892991743195514;
R2[297]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319682717941421512166618168206384403683296967597;
R2[298]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319698912380580527649602960826531286060065683805;
R2[299]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319715295681101156930027484720710787028438522247;
R2[300]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319519703194647450217145644279428625676616165859;
R2[301]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720836366992679695234960368429691694351251900;
R2[302]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375400335642248999439088224212119213183717638644613140504654316;
R2[303]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167191025172294363056130819572590027677199425114547971540672396229668960449801420589118940658996009858585330699971707059836;
R2[304]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167169588138543517422804650275276949847927654720536080437700593066827231578889385263881306113919254726255832131591328299515;
R2[305]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166564356113848078556644251551564637700397963595348187509233424146951112503775690437725667156749423573676033372478136670695;
R2[306]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275162046659995200990160362390241040177706380400701749463883514050153744076226809458042949918601770045396623668047089369152315;
R2[307]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275149142975789956154952091551956724345908582447047543275685120998828724877222698838320689369226366221446825316345822745582084;
R2[308]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275094944767628697817300496698997214902391032969165971914949871430276259269816674541549772917102185878585851957619127888703106;
R2[309]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274837316168720470411038844529967963864038903819314478468752170254701723264824242899497435493346627539865126534055523845203190;
R2[310]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275131037162883761054579736286140800915637593857264282958798513304301192061357616867899749011289618800955484237710669654027519;
R2[311]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167048232422084009701485781599208513776383871941066739187997621734472539562526300476838734437034468548951285424972535553276;
R2[312]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167131765209109560686402926464719538274591195757627359781514063395544958764437446748312767180962997418167371853940812971032;
R2[313]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208046954857764067498262597180191832604915507518860282401934296233940447605251499800334171965941116188985794926988768935;
R2[314]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274826351693479334885995153938077704414599516063560471949509803585123089384565818868722117648732886222116511565261443627241719;
R2[315]<=640'd4562440617622195218641171605700291324893228507248559930579192517897921981120365596698623783904026676499248363773831875094084271279031221979125247665373275793644201973149110303494302648819936489;
R2[316]<=640'd4562440617622195218641171605700291324893228507248218489331501706248967805011668758340141441116839476796053149040364436832791540495451606096010996116407212878859845080058073121417601802290097430;
R2[317]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677385904759295923675190790201560390877943434573019237515345107938635646482306860434693554110324286671205561839406249;
R2[318]<=640'd268690453286029085356456317902602772097047425399352240060724661718425129403641287550937335935853465073069932237380149980367813186328123390007604241383071158602989011813367640954292160714;
R2[319]<=640'd4419864348321501618058634993022157220990315116397042432748592751714922818233406218175254458183435796127359583226631121170069297959102767023371580574759539317077345214631063424033450196127226684;
R2[320]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912809287568683843723491742477746407845696897297575351282952485479164199724029506256909175572739936310687353;
R2[321]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811247366568485596508829389093769793726585330798466065179319349238446976682015664187544684335425573648629;
R2[322]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317354320193588667493732077152707911591876912375157031750160932933167206339694926931107915632710921451;
R2[323]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317369493243275092249915682824621408625008905427900156078811086706634073807369643605112460840527091413;
R2[324]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371383091243591016525568425200479202234587016892322680323463918104144590368496566014755667768311511;
R2[325]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310686644657745579162337937441562221968564358044001940010696331976506761890;
R2[326]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310686646380891269211331239846219394518258250399599400915122223390729188930;
R2[327]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399763275052108682567696236875508772488857473592234076759247585049085136149173516750679822587084;
R2[328]<=640'd4063423675069767616602293461326821961233031639268248688172093336254041945795228297356828597579533902927852832952772815933184132222682941277865199126788819135557925819180004592404578259011509577;
R2[329]<=640'd4562440617622195218634352055195536123678657622220889878404641666699257797493125113704380303661903720858132753409467620223824580279741457122181567170215074020483242007501461644023285659373170665;
R2[330]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310687841483051152612203443478337994184960013670013505065091933750113235701;
R2[331]<=640'd1140597101156162582007635009626052393822476294156172499992132361485680550019436879916054191098487326145262426872093048890352718790789303659229321582475666797689537128004856465985421531218467743;
R2[332]<=640'd71288134650346800291268306339067051951456695425758748915299883092176174487635584164154887676833928121541286087087412614221421241506803291304026386246241561107483678287714300094175007115868855;
R2[333]<=640'd4455508415646675018204269146191690746966043464109921807206242693261010905477224010259680479802120507596330380442963288378019495639930251722020726354966957749755654455496193256943516613635771;
R2[334]<=640'd2227754207823337509102134573095845373483021732054960903603121346630505452738612005129840239901060253798165190221481644184718663651325665072140133812980314499532207876581463118718318376402643;
R2[335]<=640'd556938551955834377275533643273961343370755433013740225900780336657626363184653001282460059975265063449541297555370411040633508445518879876798746564545831084319828033166352492872990387497525;
R2[336]<=640'd1113877103911668754551067286547922686741510866027480451801560673315252726369306002564920119950530126899082595110740822093425653331152828096868605881910146710947664387524819355809929481181623;
R2[337]<=640'd4215111110993863695200572007200391026487650982281725342510788680758402651055723398377993617976859611068305718802852226446849255249540513902535116039929599526239630994011254435636750207771;
R2[338]<=640'd33992831540273094316133645219357992149093959534530043084764424844825827831094543535306400144974674282808917087119775523100943529856092609784432775306167648261113432129506057279500073561;
R2[339]<=640'd16996415770136547158066822609678996074546979767265021542382212422412913915547271767653200072487337141404458543559663830734844627178094246046624643126079741031564022689947310696386280627;
R2[340]<=640'd2281220852696402253690094860988469172174488639127632517770285615180435100817583990765652970561088019484109679729470597571532095166693111363629398240465199955572846383542376325852004318945093246;
R2[341]<=640'd1087770609288739018116276647019455748771006705104961378712461595034426490595025393129804804639189577018802644512221057770022814677893703473033586383020243114827919686342225039075682254140;
R2[342]<=640'd2281220852696402253690094860988469172174488639127632517770285615180435100817583990765652970561088019484109679729470597571649548262286516165132154664836607101746705645952982529089694221460798316;
R2[343]<=640'd374262740907152241802252924413747242103139800079192966335367470998349760885914647956356695504790232823181462396245896440823464986916598168066901775062647349223426974192875250544953654078807838;
R2[344]<=640'd71288678535651444660777364477390561679331080929111301395989239322973691700880881676851452544240236119801620239800770891104960033125943521416864798512661929830498210374587673287124975004890750;
R2[345]<=640'd53466372930412422403205758823462043827529714320995337926819590434530889472349336879464448173830594292022036246692220784828886866156805141166286036486473776924990965789770343919907679369960047;
R2[346]<=640'd35644611210478044515143211307857035703602733216231926938339297776885604457063089594774008688325266260766881801277046771493807725894211022217485922863326629638761760291096901558359733321609262;
R2[347]<=640'd53467188758369388957469346030947308419341292576024166647853624780727165292217283148509295544931870889984942404307095587223122071046042380902193392161128674834676557727000642841060372744637214;
R2[348]<=640'd53466101792766120581363863705707414519677784865733630741507670918289652825713333274128532055563832405727458060612859610956507195348427081186943608348945842150018423496338336153067308207446395;
R2[349]<=640'd53466100987776309263642171133044478056810065167565204054569609338272491006182435476178197860213079446282051102862911850394511274268564568276784193229385333892980832009777900521147237502036221;
R2[350]<=640'd142576269300709809627727554056878292996130934449763640198694463203407722098279754965636922449479299590120081704034190731893840431166039962911028766526925483469562394077534546737134239955957243;
R2[351]<=640'd213864403951170073235332450047154668600110435063245385690657225429653387754430948185195663065619175050110600231633797954978955686566245599115726995324592936893837946537538939550255924033363439;
R2[352]<=640'd56731658168294825604661826261402593861498288331439566992128124969293434199911500681092848557355010665143396134013700937391438008216291377043592241761348837655300126055181385754959;
R2[353]<=640'd1013065324433836171511818326096474890383898005918563696288002096935811459197662914988502155836875715422229543064019609271044623414736634004729428215361800650726188572496545582737;
R2[354]<=640'd31410960987084275825683820169495193134461681335853903669085850407928086608772124902770760633704779215691224835351944825845882334774743423714779912166941335739598813337431061037;
R2[355]<=640'd3864537523017258344695351890931987344298927329706434998637504168063963383340965377494669888979739835394544651323289719030922088105622072078265438245006838805307202830351900;
R2[356]<=640'd867588673917374443467401194460596263577349545992724649809000579818170100953890508136936583421810936548297152331106732178429396255931722443518153303104033347242020092899768190;
R2[357]<=640'd35644067325173400640294956115740836715445797279963370790775931551548035505987332028787305428739232543486144946649108364904009031948313516122179434410741831308531341679867093393728930018246192;
R2[358]<=640'd14499563636136243664148480838249447307197234946808646093197512525106783932694026840895040720197472306507784217045376784093633844468614908459096640471541790396878029067287601;
R2[359]<=640'd35644067325173400145634154759449660967293960761678624792877151728575664952483922937778067019751781555295146028521403201148961158491664004623460837535440199187327362841075630657746752458990848;
R2[360]<=640'd141478164870616618543748231402967963324529084556702441846727387256942933651148418685918698525849186455493779845049106125838065839081109200576266717207844973726889956532841992862448739311616;
R2[361]<=640'd13523861067724179071655032015472870707560211809009326128564498071230086898849615531330834572784086352578285472805921960490827275331157341790832182756961491076821680173121404885714411905761280;
R2[362]<=640'd36758012414748149446373852723371887592979083670875726055882439424971271121379941440766289155513614736730944013342609723856690686564115305169548918212023629069139962212636627168700062408916480;
R2[363]<=640'd17822042691932577957857754307766274383182790442009862154545505393727583856146473750456028359801212961893345132568666561132906620866539786326678442067147061664068850488623064938492132050801152;
R2[364]<=640'd124755055715167809598119912817558257926609813886875969799613559042365355504808550721700004762890667404804274530849839040455709275725936173935287726079697371069124165114821654477983316651147272;
R2[365]<=640'd53466114798125947623560981863314736234620730595228101379662022304875116164137104089665696186539086255964030075724445353534701623151372568647451431269534513033725762588240759430475021759283200;
R2[366]<=640'd178220343003737266279020708596215272750692518032861540110531717580884077010011328372540430581205600936308623145530487418356619052884254796459848296795237486238356692338556436929888016698311171;
R2[367]<=640'd427728809263219162611721176698937225776623170537678934932637096120744448128437963895212365247193335865439647320243338134341417037642056300532686766617648705527295614961455286549818386233299041;
R2[368]<=640'd10180040178904511228479384408551892032852298569760408358752784629941372996007452197638651232092941614835776236686040717495196465313889001968426271568791853713764886363339132512370920;
R2[369]<=640'd71533894074056033636469645694120026249085771273287047376091222643073593082282398436649247788038580758835300245033616852829117420484542220233566350552760268471813006265212747200652;
R2[370]<=640'd554670790819934227891277900793812680103689046329018842765934006504899251850234589799369057897504521503235627023745048435592070852849126866805196038084902608090620730283851718880;
R2[371]<=640'd49794551501783389663021107033134397273008169951949519124036180009215621598830953177596645704056895262071091923727631174385724697445740942831062827549091303246875207166112660531052776;
R2[372]<=640'd16598063020179652693450132242407424513309711268794108671288295153794207437122598803838520282763007609508941742815306894600693372045124097508329299975173056755363573783263048935669768;
R2[373]<=640'd7261652253274586685856053708506640882821849149955496711175753647499167091736869971155975056039558432295708717811891979878906040619572140540189321706374920240891179317804687436152834;
R2[374]<=640'd1004960802099004762103988938317526019873565252665351147776442091611385818030872514079736453790241551185768828417989791808326614981043320200785699580477657415248510043098176638943244;
R2[375]<=640'd63823115449002457518849754259196901707970990537256506701997428051326335981056607448261808356281457079777712830552542195853099418355655126323154869278715231923895517305396244119565;
R2[376]<=640'd16707663280547663583468684316485003866434452730208260254970887845011805849383961177013864097903529842119952715891640779639438721734244452548405742491982905232005995726419387219977;
R2[377]<=640'd3926370123731163557935449223818759146879573237588170576393873110804941160181834888865137138946250434795789056767661675380193824778757821907359416635247728960170346663842414600;
R2[378]<=640'd30674766710757990986293128284654282025328605203036131127003451333509758988467359292189675913086340889168379064549905720164640092017332670528886176751216276770613784198774784;
R2[379]<=640'd945791695823256601843923843063042800537944327667589969519013233695578409010447726035717273849131364712157784079150898834862985818747335241275898030600812498265275987772567453696;
R2[380]<=640'd221546211350499102171987527546186265589391598502118820961833358454266434618626051070976753993379656690151689867412607802108765105312136464467076253159197695721610265769573089280;
R2[381]<=640'd23805430382244566229181502343829902458181142748965521873358241604279193014458458168222387178623278701989254095648542231828696301366674209008268969622617740985859836717790396416;
R2[382]<=640'd6183739330098755259692017136297814908565494341196150771039722848190127864181142967633762692572646197665012201817987822490557552973374418502914389997692288505264529777488822272;
R2[383]<=640'd3833645484546968831184162096216522188120609704354000923001160992558713395705651726571667748714436189321836008165510696644369016416281444253292923275409694216198854516414611456;
R2[384]<=640'd1221193860728625581991700486565447530201239103238857078888123752416687779541907959559815017419296486006052730868579691020464263197208786786834414222642586734744384421620613120;
R2[385]<=640'd749705183615736756175820571516261996358695176007238532457350913052806620894110528888219244475077671336949706008676476033994224392203732459840642561667994022800773999895773184;
R2[386]<=640'd479323301715409372168047328109491022288531350160125315550712582224493523284622104208988082031203017374260380878197443659824469044841448425845183183568176020206988703458918400;
R2[387]<=640'd54107298823977677840091622227828764649064246668219947051964799800595781872085347180949062149036561329209561308102625582916409395838727175568460236773014221402416712981151744;
R2[388]<=640'd15337385079642861513693013699698281333172085726447617115000681019931821955489886224554271163180141242062021200630098565954815819504862961065227384930169131755414523547222016;
R2[389]<=640'd6755392740444591082571837831607910726050966829141203085334386066223681227520067921903146976347250155331196455808428739764095153406796771048541200375799265172841787144798208;
R2[390]<=640'd3019162568836926591676157382008221160609587112048522329359793938615973582652114171887688323991276604261062351863136319501262801323320799781019112128901091783237589994045440;
R2[391]<=640'd1691206828752856148909825763688122745707934481960687741956890175582689549398601010152332425431981427384387315954245007334860913794722872888431509001938956754168771657072640;
R2[392]<=640'd467985909622883137722516648571123019420215884307945372725134515450828688055314225739475900338544951392122960438001797077435351880083093325541456540976115986122442195075072;
R2[393]<=640'd58496475170885366092370812261603197452692579379892530672861552186564894234930113950303693964469315245205088559296321058174024485650624486480760320678745824439194284457984;
R2[394]<=640'd14977913373510921199504510692714128996893858255318109533882886257090594459967212853329103081826544538864721910650520204848880202371416547757383277513662667359708453535744;
R2[395]<=640'd235685507951153722972665826584409974411370742158553277039930946734939332770205644925027659591329248585500699821007132072420722794580369980235664354492541596831525634048;
R2[396]<=640'd3685510180476565248936625222244191770180274992855786866373703244561709680071542406144003981487937983314097085123139664063073617036083632836836749592638660593953275904;
R2[397]<=640'd884983132086248398172813995178195404761384888366586678244623813784182419488154263116209441816193544063949770144508835154583066491537955544841348022719060564573885038592;
R2[398]<=640'd234058689495670328738359877855387020965687533758766996095806061823019610488243396576197893210683873131438508228548151436922584395583411808660207429333619149522673336320;
R2[399]<=640'd29304799780691819542873671826396929803252024388807047437804237452141172083575650726571882338610954648120230048288641391195750739112511341260368632672501535609098076160;
R2[400]<=640'd14742037921121281989049606664725111470989493069782606603132460892342510641975451191601736985101541958088461206948667803834501230223210051854458421536137772464921903104;
R2[401]<=640'd2994477021647944965965553601792282632683324837865389782540999629905807679328003308772963898478238430389169976819999891809511879319368678402266099654443555919245606912;
R2[402]<=640'd3232019669999832275039199659827605052288573929762341453842593588955810092613442093239988401890186325698989792637936269657398730475136318744491782603891235147862769664;
R2[403]<=640'd894159116652065566703596521669230953285407377612462766353372556367377206276772206892519921129286904160267956765096881709648359343474148557822887461105577840087138304;
R2[404]<=640'd229895274055691811132354307281316338167999345930509186707535258071038292910963274999378878059791722575290621917315247908280279918712418287036075883873731854982971392;
R2[405]<=640'd57586041745992907915898420597381151646090137594934402827328113601502181177498338818704443776143798460148280463804417671439631755097715924943200287135395086898036736;
R2[406]<=640'd14396524142538225228420667168046557606909466293138172499546817032171368286660297684175921001299630694537384917971277857773904786167114660113179573472666472293597184;
R2[407]<=640'd899782758908639276418595104949708334502382009802800812072098759487982831704577488283391568109443905483236768406843511480702707341110422890684048805510946414919680;
R2[408]<=640'd253063900943054796531473234475086522375760648609270601148380030206705168064490770613827754518783825193969165800114128133471577072432138593161228309895818571153408;
R2[409]<=640'd197706152592318562429556858574176790738493823230194411951945075320888658013911810633045613131962082404230123569116186929530527078045504889678092707142236752576512;
R2[410]<=640'd106735637245472775411438926566694911909689984872820733045091429350809793294432200416543568049207363160337837809775007861821403293009977876921901343281700822581248;
R2[411]<=640'd56236422379415701854685722367059470954979005976279993494338023247059185636521617639178910765278401246488542828428682407338258266063648971215581401701558677143552;
R2[412]<=640'd7029552803973744348135529599825476428038703526633796518262467287213676576934991026233348348592662247181741582747304315122492653191929481983495016851443038552064;
R2[413]<=640'd1757388200993436087035340449727617088891995252887437132246670023896644618625779893590962615012625545789853403307291308173316217791961392758254762439671879303168;
R2[414]<=640'd386144868290361548793405206690360332626354384071034665322380463300981254187931173875747725894827104255359858370431614838075016020484062565215334028443335524352;
R2[415]<=640'd217758133356611213591959113667267720480462237089570636297003797626667067015603894451287537532558599338527370588170046506611123261087950654950085534834329911296;
R2[416]<=640'd109836762562089755439709118371739264491458657814770040876515107273642578518515723267753369812750038827108752739220910676649216494612928222689338502082197454848;
R2[417]<=640'd13729595320261219429963801581180184558049214502421493293985843606663760500835778759109730806355031160139071770298176204976586081416078642269498035467681005568;
R2[418]<=640'd1716199415032652428745475193878425204310762692827996317066855204194301254348258752397113026332214431915946723556514123199460630083224004557676189719925358592;
R2[419]<=640'd26815615760378315939361405142356717573070896203270309055409922843094264081192168809906445549944974500019000042387237903904168802259956056930371096859901952;
R2[420]<=640'd167599081580234037803064719926319682666740871335777591713010228124291078754734258466512071289194618833969000728408570789811735084533973835103348242354536448;
R2[421]<=640'd107255916658324984512852173259669402056429655579928898603806944561516333868313129199860746456444052726071753383414373387115151077768474078719847334666043392;
R2[422]<=640'd53631231719770388398296099949500420539280005275015050066497253182436557198330303812100878400642501886859825685892354037656741462624518043181733140349583360;
R2[423]<=640'd6703903964971298549787012314980326188529390282510766634760357606843751956443539983580517359830749115023891307328641994146433654674600629658128142900920320;
R2[424]<=640'd1675975991224533142034745355087293971501757712196612238227716173886554417731458533615429380496261739847036333458449050960322959328113673950421122967142400;
R2[425]<=640'd160396139786910951630646294806091702438010338251905688898472162966716404536182254543485046997754589295095848092056673174085406331860197690007927780278272;
R2[426]<=640'd67104507461870908335270388615735454610138051382816216214327589872514018377608023142492998582723932512857038772606219484630063634180935236914140306997248;
R2[427]<=640'd52374249726338269920211035149222058170763388448662478494487746149516120070649246543317120839982482426103891113675156663495233275420830511543503550414848;
R2[428]<=640'd13093562431584567480052758787310083599329353420599727908571521489438854789518043144754945821340296129753680091505243667539514075209684543435371240751104;
R2[429]<=640'd3273386315491885185523871544487174263786483078616092327438684240428989292901802100352791267945898176134794373606156047727517662702921378519804379398144;
R2[430]<=640'd408574151504265333783029426493407213696755870967064998921119265772109300259891415009602382705706458375712653465555278472621460544756793147343580954624;
R2[431]<=640'd25673260077798720110882255617818369266377328813609326280024104538138175904225425012722710218899690039270072726172665438432085993336213952311085498368;
R2[432]<=640'd51146728248377213879742322192021865458733693812550589475904313633999829868023243017552263452319095367561392905778137111243220766926308923210983276544;
R2[433]<=640'd12786682062094304179739022232574810163650989275108368457895011911987876299571971877367498945822882137735921552836118701138652256895139440832584613888;
R2[434]<=640'd3196670515479965721477017827763305288116086322197095911296457986230125320038163068418799025325861842802145313156253751117993061237155078009207652352;
R2[435]<=640'd399571644531953470104412903178616048975559395763114851974104801109405882437918445184525562123874688820870058513338513593619250759778112041067216896;
R2[436]<=640'd8976551373442800511802080877280542578942990268278143577222200900643701156194105840938890257556533367876320799282262367815417081148610347014291456;
R2[437]<=640'd20315754237603248830572944788975586844502602560972627584707401388246786791364716115753075485465689674799689420232302967609973755749567409139220480;
R2[438]<=640'd6243497100543968835993023312683875431635758236248056043197583997888531773832500701445630426349202994772284055475689659190137156374437614946615296;
R2[439]<=640'd3121748381689408194800798622350042875749894161548096043494253541482062224437823297725334140377068916281775104033209488706254843524141712960126976;
R2[440]<=640'd768052363929141175456530771642564437159245870476695895827862943096777811966462375506203344776437409803219690077797473664299217262644528364388352;
R2[441]<=640'd192203604133987863977428357272574249934337887221443870702066697271526636270926545997007587979073238359308895440482071344068365957109384392736768;
R2[442]<=640'd91457477060038834903757731341596669113728461210887826685326864051524562660735320901962092863188241342573054622697459655140077412479148983582720;
R2[443]<=640'd0;
R2[444]<=640'd0;
R2[445]<=640'd21778071482940061661655974875633165533184;
R2[446]<=640'd65334214448820184984967924626899496599552;
R2[447]<=640'd0;
R2[448]<=640'd45319992531426404797412790468393612409231638528;
R2[449]<=640'd46624053413417497702067085763764453759452062683366688608435179768437036024921201836032;
R2[450]<=640'd15541351137805832567355695254588151253139332765025311027195494652925188550906938916864;
R2[451]<=640'd803469022129495137770981046170581301261101496891396417650688;
R2[452]<=640'd678469272874899582559986240285280710077753816400237679918696781296365993984;
R2[453]<=640'd355713524293459643974404252608769348018815418810786612808440337637902899709214720;
R2[454]<=640'd44464162267129419042701475057219250061766360426991637922480531102594354057838592;
R2[455]<=640'd11116040566783934444654939712775920397735190429570609922836692619316169004810240;
R2[456]<=640'd3242178891717664676772703452897075966278014122757027664704575195608880252977152;
R2[457]<=640'd4697085165547666455779458516860474227386151661001933510370332413379123606907022556448096753022106007809032192;
R2[458]<=640'd923500966924488829278022197228215698066556395550363133734219840601958530374065073796839186134776681109304419287040;
R2[459]<=640'd1047775431747339879783085894401810730942240901044108145917452877824;
R2[460]<=640'd421243369770776117191986708383149396995645111076943482481371250688;
R2[461]<=640'd3451083797812275812103026726952231647375189116249281956525473819262976;
R2[462]<=640'd1763396612854104999380915335294456793213082997036555954013003923559809024;
R2[463]<=640'd35835915874844867368919076489097841541710281551729842608263778485520615045155134942352815619283076775936;
R2[464]<=640'd363148590109069717659969773082973616634517417042783895340709839919758156954869649142083435796302002488475514173650894848;
R2[465]<=640'd452312848586557221318397203873964462218103800933031801144126796120044077056;
R2[466]<=640'd411300375794051806414273529149521056864092852907821166514667520;
R2[467]<=640'd1496577676626844588240573268701473812127674924007424;
R2[468]<=640'd14059105607947488696282932836518693308967803494693489478439861164411992439598399594747002144074658941410553812617265953811549610338989507167729172124686146863104;
R2[469]<=640'd899782758908639276562107701537196371773939423660383331317236280070033971913258767642482191972143269246809666598313998403260662951701816310520112444211076452581376;
R2[470]<=640'd29484081443918291814387145163970850710288447034503440846700267297937114476521137939757614391330493613525036201168021768995954654580570062585473556792185340236214042624;
R2[471]<=640'd29484081443918291814387145163970850710288447034503440846689662160336776385851449503937737541316250297015122067400604549221140694297362454646438796363297256941511770112;
R2[472]<=640'd58968162887836583628774290327941701420576894069006881693378223441337877537377325813845730080900918242835443359855697048449577589100606156471145007514246146632752037888;
R2[473]<=640'd29584878800134287930722386670093179833839425207399327632747302561383142559580160;
R2[474]<=640'd531137992816767098689588206552468627329593117727031923199444138200403559862026514030549418879174025967298819387356718762814956359087467335008708378441200426944177632620777891654795264;
R2[475]<=640'd88452244331754875443161435491912552130865341103510322540067848905696798082084589544649172431600960547756767168927407058847087928182299714412623384405371510984139603968;
R2[476]<=640'd176904488663509750886322870983825104261730682207020645080134670324013632612131977441537190242702754728506330079567055229676746154527766187941064587990629622446234271744;
R2[477]<=640'd4925250775552716605480106115619086735260396705504526859196102756065684232401866968266670655410341330804081038458880;
R2[478]<=640'd4925250774549310721753901806147423365323302577916192840932073260485378881101130256542321251256160099296799751405572;
R2[479]<=640'd141083529341953760589421867365499479134423171896242854599852349209482195588038876977863446004799405496345290923173929502870581315425651915021375070161120152958842242806470868040811520;
R3[0]<=640'd4562440617555802969539075718364092799074169928832360790863313527499344649933626941523306280974976086995488648864983241124907892094457115581046072914796024190906171255367286041228450039867637759;
R3[1]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
R3[2]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
R3[3]<=640'd2281220308279959616503818704160557455894145626294686847562564335750193445403935133392104162919523197624091869117907874169097851345341139661473623420451587115359409985236301204206043877091573759;
R3[4]<=640'd2281220308811097609320585802850145662446614253624279965289596258949637583604338693252956405658685699889321154786797203655344352360687718999126330659861107094125997337180132475041437096123301887;
R3[5]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
R3[6]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
R3[7]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573579585923266328248361220912171549267516995630214792682163214379329861311652691967;
R3[8]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309569800132130560326787237530613030482371842041861364826120753951170008879411130007551;
R3[9]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594378362666395392326582105506409147745250870755828264219255085686872213964193791;
R3[10]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594378362666395392326582105506409147745250870755828264219255085686872213964193791;
R3[11]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594059482108144189522778911973475065811514326462120152509693298127605327909093375;
R3[12]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778626395229998840359290081487658414870654811609972474940181023171096377389966779635053101055;
R3[13]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573564388190351765720371265265389588970696231754797620595625608073969548297876013055;
R3[14]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594305978475845551475760798930139721583952488303199901259256556730234865081909247;
R3[15]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371387246796484867605105803548872564030266032400453759989942736265474793931889569167873019490598911;
R3[16]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371349704223814961832723894157034570063743756381000379202542436027421475442626050865800790050603007;
R3[17]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399766420093704148998205791938233432942613563651103485571377357479647437246027015537230985822207;
R3[18]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399774568225949757357539305044428552119521518461418787246166272833962692411027903981006792687615;
R3[19]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642185713297761151957855437529246393074081395151850507260970814444796097981995214805401599;
R3[20]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371324685347959954397802122066373880421417186681143452577526403205904622519525942177820731670265855;
R3[21]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912793399413454012508970754755806357124447186848688372490820743067871944960818731674825577043622421269053439;
R3[22]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371349699067393569240749173275557250543433790461562439074608862111696438301066772294215604543422463;
R3[23]<=640'd4562440617622195218641171605700290006852077762171494654054239094271777451477099757786466377464371911974310560577143501026943050191202448660411484268834096775185635538140468495675059706584367103;
R3[24]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386496518067595893676915788334041687995441666214086284678547427685751509471453813287981677145070978155014340476927;
R3[25]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386496508606437918483871184164450525958861326492606102445612453836211903000701028318978997269218606199323590918143;
R3[26]<=640'd4562440617622195218641171605700270236234816586015515506179937739859311715503435346262231073195066477437191381461825361624296650106127709648759056807682191722715783472650501150100268661289779199;
R3[27]<=640'd4562440617622195218641171605649854283524716891550644909028181705653353172171464492999663030637004212451560351020607260232495079794179583924395249892477611505359443129630735248354440689167106047;
R3[28]<=640'd4562440617622195218641171605699419660345535762949390388743328358914119163392006390153554201760580352558929149082579524284227176006587709005001050786042664526573950431557756521451689192837873663;
R3[29]<=640'd4562440617622195218641171604775340130864061735765975226214720837847287943829637458685381799672364864488020246547294248320996321819114726664605758380433291953310065435824862784185936801012121599;
R3[30]<=640'd4562440617622195218641171580651014263782655089306658540270211210293923543382315663127695339510122751608100785650218030529559615331613782175937589235910385529177455993633198167738126477538885631;
R3[31]<=640'd4562440617622195218641171580413023361305561941806391979231826014949671967402373917261297781823655842027717261989339332133240812600258871598400758798420297436862115145414916150285558884228661247;
R3[32]<=640'd4562440617622195218639775772173727602939363479220932161647903947906094238376758280112663959117799773964849219389673445750716576737348621388590559991230537070918170551495697188673232592277864447;
R3[33]<=640'd4562440617622195218392650519082155635791918763402178406453631627662006624130865912053562214482519721532243023452860444953296707786506172118195791504821601087895986042541464992611645021539532799;
R3[34]<=640'd4562440617622195218393601557613210664319946098599213386615964039063006782895847304853789712532429336253212356753546306704979704079048884590532787234520569679823361602077988186746670323203047423;
R3[35]<=640'd4562440617622195218628611873492526396639499902442827511989086075399181865818151234769714874212894553734555181022441726465111896499232916940836711518365667664462798846852714577323557490561908735;
R3[36]<=640'd4562440617622195186970320484935145597531354314680761384181815816439678552831034409049290516897172603820977208958648499207807229087590714054953913248116750874170331911582577146309353581047709695;
R3[37]<=640'd4562440617622195218503014389252424339113303530096313439787348143206939308514470923899742931075310625773190051041211955367218676916745803283409515048966458131669799189399975571294034602632413183;
R3[38]<=640'd4562440617622195214931215583603723313988387210800846946675903060637992637297225319739723888078885291594053659689415184709370057524139776135831077815125929850336918608950567968797747581831610367;
R3[39]<=640'd4562440617091057127645828734757254874789629046406725009000485254880770765447766191827954937056762674776985546706931217932495038250400930931738211427487739374834457976282467275859791110991773695;
R3[40]<=640'd4562439529839135863350193458320745280058466961308902942516902972448249059127890386829862401833240428201357497388377117733745895226659080861073294985037930836899283522071821747958854288343302143;
R3[41]<=640'd4562440617622194433367146928593395682797724269870301589083145678467518606554027372069832685149837596916585209192963353951447866640480129065025002117649426105130833461750049554290052118456827903;
R3[42]<=640'd4562440617622194712355839790255310103044567980030774170652820771916839828124742892853885427034833178925773158751255868994232571822666196912108916959475755089020752759990996713675837189891522559;
R3[43]<=640'd4562440617618551729201845313909449070283422535305294384314843729464983952039876781836951378264783820921759777327881829757315149449134990864046027733946755149745935694331095779882207509565407231;
R3[44]<=640'd4562440617618301232971233353637352593330133836631226660375987986646325471173603841418322050216371065350613894226932689473091719657718755325914086570935561562914839667926960989313180111567060991;
R3[45]<=640'd4562440617622077893013285612048678112433389833500045207952950038619076924925023469864146149376833333828235876881910333115171444787479968690200916157989787427444615305383676299210468587103846399;
R3[46]<=640'd4562440617609625104095596566484172683103023446808676524127535618784897110257425835355021703493829480633960833490080617880742393263362833555209778588080979506005757009178539807361118721567883263;
R3[47]<=640'd4562440617589493469968447374083889829326834297786967702953876493591992833823218453978596748610813768596410603729946410670387884964592462454433305164382488252086041091548095789636214727763034111;
R3[48]<=640'd4562440566583154481203951541374803235355690922151639252468584177744441326217629603332530748212507293664128761286575453899326671822432149679632035369069284037725462739612995402721247238450774015;
R3[49]<=640'd4562440563315410464177507369628196286789738467491892462091794499006327100888738303030512858601179575485691280715096012134879593101034635852702343641348587766540253012118772125559649458249007103;
R3[50]<=640'd4562440613519880452672782719205722820140199695358560923244852412140197622049692440970121036653939917609545373242275672200191921516441447884715105618030812077797582650073483298274699406580645887;
R3[51]<=640'd4562440341567891657141463178865147428094312008987425994163320470295232305075862862881266367225727935658944708760122633506042194446677044579840664611656522645927819227557716313026159533039288319;
R3[52]<=640'd4560769529363903430937837029134006347490610521661753866819401502382131705995258068196286454312303798844869523366600076626100939095444391177816286234255551384918472140604135408793562742379249663;
R3[53]<=640'd4560769801899936986005235768188528182771546807245655146032642778040859407694686196051453517352885505471207740324390783671228395513326797985301286245642339307877226033721654649941415269119295487;
R3[54]<=640'd4562440602617547428100163284637735522611367094546058821541686928961199630071656606834657558139224524953230415630340483542751307159995966876006632576858937457862821548072194235457170275435544575;
R3[55]<=640'd4553459968394650674301111181637262975666464563325715848253176362122640830944051010751485344545582886070697098961515647728887600088771071623504257321309545180858142064318999219702576442455883775;
R3[56]<=640'd4562204975077302902990209472637109666432327332486208327355100163902092982430483374426362262008900992124233007019910827242656865524045617918948387618672751653223655478167772613453479276831571967;
R3[57]<=640'd4562431912204100702726328196042201936533559076471037164694887245901010130102261631123805957970147592796795302731752012347744570145084674523685821794492606684016118201516010607771724290304507903;
R3[58]<=640'd4542947767175072780700897844391951713335416702798731856055691376701806334104844447256030629858516574589541857457972636465726469920927369280236933649833513254306300993172576774743717223845593087;
R3[59]<=640'd4559057378036902236967624736083570523798163303018054624351073096825240061500878360337825196648322044000010415703313189758550858679975677418517383741305946919517591977540494132759493624016666623;
R3[60]<=640'd4546595877934823789514239643290650371499399403317780494449434436070701885055375494146709656205476510259149785965285032521874652292525447674358921267845285383786772584628132264287111379941326847;
R3[61]<=640'd4548830431692649716190055397749529431221020090326276668837011476223373222274103995821813653819799841154091981869907622062938433324191338704481704880188910964244813305647127866605681660068364287;
R3[62]<=640'd4495119565321116430310330316503924646754195845619411377053946238023248765480056506915621640543946205979415684155880273381442500055729121398408258643531904905776436603979935749349677292090032127;
R3[63]<=640'd2227665536472437267808719731748435166023796555582449549738629794632581066412893453630879456733835160773080162105394497513958968414089537276535651016701036759519560844710829394931358654765465599;
R3[64]<=640'd4562197780850535586733457324527801806625627656128168851721345342555107386192329462136743326909221757809796600802175142567648850862569295170518448790413688494965698449795902806936278297704923135;
R3[65]<=640'd4562301658694618718775566837435818828998494285782404997219703787655856800634890788740424657424287550182656224717251613606878692100991482807808735188985294767259203971594845799040489474602516479;
R3[66]<=640'd3706913588456028377487358498978764367639160486680879889392885951150277770536152116162311757253805264948119781120363481437244649511065509393327902479829876394863760656343549092163757826747859967;
R3[67]<=640'd4561535830425087769689760005214053156628980386626054257170645590718181683052129521021414358525902108267735787376192260527775523738408484361807749320345777402089859668662870890861360085042398207;
R3[68]<=640'd1121082734377418143718733489955720918668667294459803858228998489773637475404341627498827719443858718560848500899613758944703479707269391416429561449301574212775870346793917992554767439973519231;
R3[69]<=640'd549106807525952802506392797031514930614092113452506368690684498846868549444968651400676297260070433530288227225426926756158914347555367327656514625839020449058284732956115980954597784483381119;
R3[70]<=640'd2558472100721396333713124466224592440730806571847738035589832532349589036687492863214390799269726090470224698910860441968952907139444306489818772766693042565005341438147514656769821040836845567;
R3[71]<=640'd3556331946777869282082116463561759945569769976942524631385540296500103724205133386887792106205708872537097591020151042048577891902712995476661749014110905353481567342065980671963969067519182799;
R3[72]<=640'd2568045668645413189730805073506268004674538404192971852022202462459833054084108212098235016235434616027901716218291399953655478013530817875604413371690475025745303050467611870579698148458039359;
R3[73]<=640'd2737353921914897264360301649205505812237502895373721063519998975298376917220162309726779382600729634230437118369983380586100661078612400753268228843817084750758810701710773246786152349827268671;
R3[74]<=640'd206651258944968640096884225245730360838148355563808273852502001164926558983803101921294725139705175600646426693787678904550351691035326918654715742107270126999614983989910680317904875034968895;
R3[75]<=640'd284135334985824097947731444377405734204358199902647871522118976759460190215423264433230577098642825741322518709379408208464301389887579663790088612614319107316366939489369175919206270781063999;
R3[76]<=640'd140846274249666453264347980255159685163881711095466109560684087202595742745551096584930001710669643705690627710416646638717229760708458643272400103817734960729865796522311442436903622415483711;
R3[77]<=640'd693259154461003060611610752109324464049963796479513457367806890170943637163439910836785553645751356124556909583085032298797169051391509000168436332038775903550086548456788074226576616431550719;
R3[78]<=640'd6683364601964633374124181971721159900379894700336373945609559328291062702089077768840963424053324204653828835188407056821305340010592237361210607286179859935785593546077678400082335453020415;
R3[79]<=640'd2506325462295875523298949308146707387922551842902328164718153727326113199008996927536495875708667642329018840194691185318509555387635648365826431577246619166342786688579580870235638062252287;
R3[80]<=640'd17826121300579417916273129178621649131115454295979812676022481073395265587224994403051232902403632840512858524980042763928193963874230585702551359706239091453393674975071936356882104023254015;
R3[81]<=640'd3421830463216646414035948363978214425081830144882191645659999416707729293048981775593657144361502260902995447954157398103482027160995848515565300453385608403713131305761391585094566120515437567;
R3[82]<=640'd135971326161366759428668806219905338580631997140503326778495988798253765807519514855150837788130486121385245912134800063550959657538390373629295420215031723479789687549948290474461638911;
R3[83]<=640'd26733186465206211209331954457765538603155560942349498444401320826320591912809516384920598651380776192552456906798143610101559540376302241053609661959411639868960309693598969269930330100343743;
R3[84]<=640'd6183260036820415089441293706691767610483134738633846882330979899568689669917234164961908114913601787182383993215710175168610865598523910727230753104603251183771771019976508351;
R3[85]<=640'd61832600368276133515125630254911506959363832452222124887618528336008442721990343338480387635267503172770725225840335806738365788080613696466521768393654433567028242739626943;
R3[86]<=640'd309163001841380667575624877883951091122938103057304936651485773592716105610269726480930722335758212569550082450013664556375171312418022439802851970623126425022791582876700735;
R3[87]<=640'd8911016831293350283738939730396387956997676161944833080263623391415450053056810051119745049623725167740698600154237941008716040993206969717156488034377354449125403598171223045243610379335742;
R3[88]<=640'd588127110865361102650293919732989682181647364492347114271163799187474612233035841549293499712343136996243203119796563039397339966092581422399373018902517052310837942318437497572386409185046591;
R3[89]<=640'd3957286423564273848414586863959678446247055142027708298853100995817524890190729056924142519341923915733176877351073936221939449358743344729048490158519992807112577645082050623;
R3[90]<=640'd3957286408813326683052798039200490885979005839599766677793737440334103854135023866908611718238662410012735735488638271878729428916435542841415685029480823998357623283690505247;
R3[91]<=640'd1978643182301521049821351671732156087712550892148766319685274665159369719582195451268219554733857704347796182032418834652574709507383798481263762762695016843932602493013329439;
R3[92]<=640'd65295225959415831877930552553295379371286832413236566284319410765132313761020833841316522179307881386505483137875636186463851116459515510094001651415177710196578980872660715038;
R3[93]<=640'd1978639378854361914644891047119827976894918023449398243790388428076283023967333951979693015708013135414925384504429910930266398742433715001170392242771731935227918520093247006;
R3[94]<=640'd7914572788171309612743702550516101946123417307088949723533464487031588862294357656079701021745602689395382686726399394950180128819691181515023957403227493942132422990433878078;
R3[95]<=640'd7914571903648873324742305374062717538489283328563544066691700503652663787653248998617826127324251244261363558240033631594513112034801404141224197747301504375668674958515503518;
R3[96]<=640'd3341631311735105195811904120256403658736038330154291270064598172507303420550124821744569837778287317210550584521464036037197773565257951749193225468152451945947486905979336281635705491298311;
R3[97]<=640'd2034045217940849263834350395781531464255597036811573949444865405510174615379545553766883971872721560803286730598178714264003120241596047561388773614622393115369587410347799611648;
R3[98]<=640'd3055025115221824779893785787393503681025983702890231728554390195564082403502850298623444913575435069103817994887063962584634305615443573853291060625237998827377017602655578489656;
R3[99]<=640'd3055025115221824779893785787597900167357923294239941837914200288016783424168435231549898532325557233500547673687437530481419656208917347853190526402524649084553449571758182007056;
R3[100]<=640'd569849237446107996832315103946170450858604656786826655475037182467606797651054148412840576181131577987853926826265446961673737623489270578811905416078154917282065354007450222593;
R3[101]<=640'd253266323560534193234871877041022047613636529937275503029421663799622050743876728780716410272620665571239540014213842852020307839607169095009963345497628417376285485200132015107;
R3[102]<=640'd4052261290187419836404190599902792155542613226743289225139840551601650748557661705106943941697662427006061315548025360643852529440468715791779894509763671229015577290038900164096;
R3[103]<=640'd16209045183393482687594295589517339425247856368435233969124104170986711620092322987042870998569661925517633482945440441044334415043941757899950153324382512270289774443248597598208;
R3[104]<=640'd8104522557731065123879133086356303273359628287500867966244382418353061816306457786294970847045136393744020627975351019984081969467263666616849523455642302581087085609042065752079;
R3[105]<=640'd8104522557731065123879133086356253325382825412141339255200354304362900383269256678995777755783502787905108336072466439707205601318980296032406534684708169504392664111523523723279;
R3[106]<=640'd4052261237351974681950896744977876271461234370940277527721904539542226434301159214269812418003983808999720309408938171519762698917007083797849116072658181216857588839155782123569;
R3[107]<=640'd12156783625254732488426186797742726594878858179107925848781152391509268130313601139684491457051677447240521835957516752105662566885223188393774460900190932329264677649618909003825;
R3[108]<=640'd15955778474888786561258759249585331712872466039040338040554214909837756295583577995338022089566541833250195429340308175560172547429314084025803559691700586601711712258361636421681;
R3[109]<=640'd16209044928651017212574736596590612924852660719833991630078992536124634380064779019641020358391159459862413551701123275213279545943308220325617251173034409032140922750961700569136;
R3[110]<=640'd531146097339326716757519282670135830767856534095814752450020956955283076674793356600555365694592283102190472623371212613979607183271737782812657590415489016560376068372218769225809920;
R3[111]<=640'd232380976379893336763413505714310893188718046600286725117126429437585010229854031775627067584558544186684772178807381300428075512245997844470010051448912585602996895338945233496834048;
R3[112]<=640'd142743343674028740034653226899688696825923541809343296854252187350614524186433124149559081593700497986721265014399523102238213702471986474045636614775245342795394637142981529822933549059;
R3[113]<=640'd1078890256954235901723595831165061288999759981966929652588548793593145714677461414137595391445414725448681220434337981880090801746071122432483323588834837464141597643825409241462603779;
R3[114]<=640'd52068137567363886810830801429770108788956574938244908777994222765945396216968913758546155337101114092824576065625990487247257841746344112416202781669384107937563853801099304400458874881;
R3[115]<=640'd52051539504593702036051329161417635616947823080756805650185665600132128160766039952326104157625765230535128811333218048095842458202718408775829196976094945076993804072909689557125955584;
R3[116]<=640'd16398893632740249451032626196688285381257292488909675513270993819578264347615378271709548126355386289314665938728419703940620095752209326869789500102860874731494301244806053005325500428;
R3[117]<=640'd152905507302218289903063502650388783537110634742299442889813254521173477849493162373590201970467140806568843638796958330299451154083806312605256265492407049060077853877285627285431386116;
R3[118]<=640'd17822305543012497769543878692674240293581825293819916181859360713925093811596373842892090564464233690317629971200191246769892665498823353500158285770977997759976046289122023723648875340234752;
R3[119]<=640'd1087741578888801927944632401989326643933733232771815796369538088394301315713075643182943579196758356349027775815630715173530977936735209085175102177242508358364293528775332662072427151393;
R3[120]<=640'd509882107419696794521443243130433367927047352492157779033874666612456791969316035567019950675918516584298826726319881942385578970699838164290789556926672687659240364370308214745666159360;
R3[121]<=640'd17822577545832795702967134713846442794240510376656085238417750831484609785401948330588511615982251510440977936401095448676465959098585387770303312893317821632950138455585799706253869893812224;
R3[122]<=640'd1087768615576180483265180291145927965563423830780014464727029625324916653583851687647931238626242288605860748568969477996081980351517596789551643029276692549457439755433168743380132298752;
R3[123]<=640'd8702162815761172891601155807603768287362655424159450657253582238525212805871473924735167422529756413150687724443441429745267789159404036930132888700250503362958554524083715556729677676544;
R3[124]<=640'd303252225711881388555920343984920510793883906307010872610489164625154686904661384067478309394531776581169681788549179378387446306049913440640905421253164558655279697765542253958760767953043460;
R3[125]<=640'd18363743425890924264903265988726836468033611537903123563897552087701236822340054560728662866427089225819344552186832267931111792248854021553730280438373200437506531393290029633545514677960704;
R3[126]<=640'd2282303728337937036598702796504095912599012278278265556131402888689101535046271403282904994047079877692002022993310062121248631759792864414204208901989040078644549566737265169913341676231852032;
R3[127]<=640'd267329689110843534537973691751892096566476653642436300536981143763614652647765130761474475715870017607417044545767938182536963504624354459900660298610574424915247282494002039774401637765890049;
R3[128]<=640'd4127610843182653215015326435839362384121652903653232467904747774233227156548447792534276637991771631888213515919352906048253896790651050750008098858953481261143331695360305624008197472285360128;
R3[129]<=640'd552483043540171366577946714548929926632620688430160959831700982681533340158430147176780022691802514140684447026280029151065778688609235716608268776678523827211307849610462872639712796952494080;
R3[130]<=640'd4562414511127572161279291229577760937233255785445592431906653383915538304301285306800913872050005204174443789387213158647109851953780378772616099152666411067633539219575433271760824312608587776;
R3[131]<=640'd4562440617622195217651608488325745747861775105512000125448961198569413341019308769532603021343531916582864706993925313925497283880911370914309047404215276161820928032002447388194417288060862464;
R3[132]<=640'd4562440617622195217776964424228618394070018535652511789839699231638572338631311337968223729645961083134758742540807952884422813549677880972120542664993250113823298901570538667533806004013629440;
R3[133]<=640'd4562440617622195217652333066999150568050264140279269469645090141112297621698460483841122290544409308516574589701982464280313466758992710877114716962012651586348452430144183073158556216209702912;
R3[134]<=640'd4562440617622195218146510979658571030118736816917950692018354770311680420249226195047872890698170439934420912188823560282662153433663848990180758814411391128744664355467564216842482522047643648;
R3[135]<=640'd4562440617622195216167869684339028557405277211658723542822899640927200800206237054789688700784917073278329485910015386384619154788844235971388943284893755600771556426749766778543513311025037312;
R3[136]<=640'd4562440617622195183041051958407348202977983332602672151756238327302517564778967217654459500241117662223662409234618746713807817731845396843694598122941479746350638120960475867272433340499623936;
R3[137]<=640'd4562440604076101640195548869803415602536734767785387001199418074375320278967939416936901402831814517610886453148133669933093100778350650523652797833947595692271178171529203419072963730491834368;
R3[138]<=640'd4562431900718241598294188828720999442457985934853753701796707500473129805486120300739311242637689287496950309501079928642786044343534969262466910135331058979467797350055653785089598716431564800;
R3[139]<=640'd4562370930458554658340442133847713646581265771752455326846106924664779822473705981325309507092411801049019476003005726753950069352471651333826981383945184770158838970373254209770205263777759232;
R3[140]<=640'd4562440532670200298514004359904629881256427178406103639402845532114278918530053337916830956419052360859927350451705845094807146719037172323614328147067639718794808187321743442135585157573246976;
R3[141]<=640'd4562404585234248249908654711052693795581858633420750109962823158129585269356577173769592463911145705664106547857876573073792681022980046855235063469731133819820623512195790829332407279316631552;
R3[142]<=640'd4562398874433362598230069217245341013244194897805906128579088862623694174910365142813422785849703603852789430603650498208248503520875043714224982597012675108601060181122752661370698874056867840;
R3[143]<=640'd4562294329475811101410436104516224286631838686482749770159571307034770912874167101497577410782044885682821414376605904774481432166541486603274441429786468352554491879209792997804991069879795712;
R3[144]<=640'd4562438102158885463925964866815445392661998573690326212763191689996096501462326580084720089936638966379323861950655735969111797419054951835262261988793407815350253172786034681043425840796270592;
R3[145]<=640'd4562440579386224632798160075571494856116332087759130957315443416460173306492787901592375744296944310195713000484700537353585989131081402062051848239184044505660355151571190893504814734695727104;
R3[146]<=640'd4562440613912528300061552682097209283843714057895047827972959463711793479855327268793806480865652220431737349360623756175559823956285472194543431703474394291222516981632756820596253228009521152;
R3[147]<=640'd3956491472670996828139518575988547525217541313809429482173163656454070564422858438500769076520672788294295292341600464384034230111004417779415544844725501297516297423894327392573135486525112320;
R3[148]<=640'd4562440617489410720436979108207210124695948084131459896711475989762900348858684615597780924429903586297593527801495577927323482742096054047173735288850309822957567764380685748868304162481242112;
R3[149]<=640'd4562440617622195218641170175715143032785015840712115902921239760828956130765517422646299317014667905361037654990492479356139719433920487886323285478655790380461224634893146477527981000558116864;
R3[150]<=640'd3876292321612607265837713213688966482403899576989949462972395017346775421180217216643327260857078787152470974725091951789720166288032275605288561938891820276778042538643501468724132206985871360;
R3[151]<=640'd3733437583035935748066539777683400734250410703360242263460778219871451420926890618209195189502542161060945154025108946267350439774641742027433875817196942028945602729239769988402054524208939008;
R3[152]<=640'd3486017631329556325961883956660743027893968653525162950063488159118330906920429849299172829911581730421783072249159385447007046659141329592075198306017382147859120804194009562235371067155677184;
R3[153]<=640'd10860301763138770356872906043054936281710883379046354270358510408675513484937896255339083900037352442774395655116248431545810480135988649737685492367192064250886653433325954082068131929391104;
R3[154]<=640'd583358324514239270547541770475870596103454879355497974969573367408459901410457894455466289151215291749323959784172888347820709858536407043340948129244033717141521680589699215913833549922041856;
R3[155]<=640'd4000437405709512472497288578356234488495124804878446189817510429982712162857624402015815391217273954515966940147835460829829659205667902773328620496260486938711866628082707511028857326268055552;
R3[156]<=640'd4048351525507462848272613529159455914481841840576485555508867966617484990153223359795798295401084401549674413280591829205958588076714749764925328293351879271868177587876934119112622399713968128;
R3[157]<=640'd3994417683157708590152707099249696219954826129349800517914959829982879398776411449920045574258118483142741308746772765165871623807001585396407592502055189232207942427781584319025653968110878720;
R3[158]<=640'd950732857625456353257082979896185531387794600246406394697698812962963546838129903108756955969731440788304794288633916153017644629921594438884721242368187676050260909870280126708361986048;
R3[159]<=640'd1141657616952562678235900288092161120914636730164977707934633869683638812998672355764912969106956577580027332995552506060058004672910915440725297062423724188806111683397250219962752468845985792;
R3[160]<=640'd4010460270164372179649334257410022459681003958468499253028276959934299726850719625784042715590175037071955391118614227369888343935169683239799966222443914321622289601537866717466380085298987264;
R3[161]<=640'd998569915131706262314568373423187406413986556723253023722115381081814725922611191349294915065737983030003815514455338053755964032771678101962884488172572615237369243923179064980991762745917440;
R3[162]<=640'd998561315144503320527994053619570674874540482917375039914613473464948466213701951909295100182930013340619655991751222061463551250998633404048978624506400972668488807254016066805651931811151872;
R3[163]<=640'd4491217646582586199431603860563198913089821424972072091829921931971169314919183355956719409837149710013296456136995577285227204238155140586288201773362230116549907457945651668938995565264896;
R3[164]<=640'd2306840110597479468412906697434420570855804614590305193991689517403969654635301155813438638738396160444103464081283439860469129531211181247298743812858707736599068268820115084623999376583229440;
R3[165]<=640'd146893204994146334219834801068973316474657262003724018297195777708632257860526713610093542867923110262725913266815277558963212311225750311112865185878837942108906244858757846350002143239274496;
R3[166]<=640'd428016639150766024138333612034300883465421091234337502626706679839740986961322405994492480762640527544112174388581773826063270763453429893315877532611149945821885919091765786244162016545538048;
R3[167]<=640'd2423797361951902584611072604030030530732879336345416569072356761672927529888984770825055298534031712185556523940180902901001336746256467292147243836079768027803047041844752748186072093267197952;
R3[168]<=640'd1158432254164108586382489482667990683935734242599561238948563123079250754806444841936176384397671499772435618009682118527219038130570929903988874246909602132693921349355853717804493848616632320;
R3[169]<=640'd1924779696241909929283410649311356134365336262593743738461270120772796260006606558636715593614553617828577745525191123348112530879223732899181676676134175352058023815252730871109828995964469248;
R3[170]<=640'd427728860484858664598353950261554643958258421563567070032024571692079908596182017466416768147415589178779740027062267035437357920652180264699197647224957744909968867744770086057049640543322112;
R3[171]<=640'd2436049244844748658508410846366069228306675164512956737326665204855704631146790196417015440845481913185500491357582755627617211764133806369650192126357744715865001838486984149823316490966728704;
R3[172]<=640'd2311295156331766424524800306317433878374454139285069050054259642627783728146214907685560501246212904718585547420772725637910832536481547586055155068955343267845406475224479695339722043985690624;
R3[173]<=640'd231689866640508757653302583108972669160220235780616052436168180500514613302728768921105790832757000505550178942966369302981531929109753864945865967161934079394067098509974188111550743366729728;
R3[174]<=640'd1354616205423341537884578981446808082644127906746004001071596465849678384143121816668985020415314506149405536562325057501547151113461948065526913123639498480379517953043908735720163459595141120;
R3[175]<=640'd1720244160028538624165740130134191951595715933260572833620770672391475092680003673423064155532997760565795310920451321568819903020032212682136451097552414476449216689279575255803305146692108288;
R3[176]<=640'd44840225326490950759471646493276948135235579281673650087425175500451994421571383749575945993737961740832477358374705248821705186236391033244508868322315815163284373685603898032819840579532800;
R3[177]<=640'd1149939837141302395298017653787405582269523272654365750457138324653281548817099185627685679594456899071679278782907111868360647464743998755234266750129630674234334073104287895248178784518092800;
R3[178]<=640'd3431282944541799310630577356816757943349990272464969225994715718265918718396190537696104559007690338994134011185473028295650590573967972377715593730354102722699669951286229402082305661049176064;
R3[179]<=640'd1274275196399070854855815142625611897879291836183858119870021128263170125203676321281483099928128676554738818852968454200404563286396754013954907841770310153583047986513887414605633836606783552;
R3[180]<=640'd828724413267881594017531068395204259225632442322902849275888897028688257993167835852396918612309606876183900644847218785969365461637399219974814355038209275153374905179602078703369245907533824;
R3[181]<=640'd2218827809351958621419215787169147218185351788715367355348532977719491844728376254258093130976281289848592643466854180247111659136808264944788623394928346051812442403306840554206240546133670912;
R3[182]<=640'd695059285337892112296644657789151094172379087313523200246303495614375223008622614188123519100164856141080693873507046262990418014210846022823714583526668834590093158595446147302276583036763136;
R3[183]<=640'd138676822822792224849678440724923247671387139125741027466259548136673943302846061750529432233464137709972313768648601645718857073541393613937700596984703097800963894097389707372320417650295040;
R3[184]<=640'd463303117393214013702685196129523844217824495363905262982661371256752949988644940349158347700850563820102138729890898033249690769485404054529136145081668578678980629967660228475021195848147968;
R3[185]<=640'd4562440587874318105333333086124881517110397825414804659488258963333495619669208758280890882988579098261066139940332178241954893469388903064244471518624327163435548530037390085523049057340964864;
R3[186]<=640'd4562440604870733875469880244191665450519848092355748137382100692634684161101309006952356243129199592344191810380749409894922579867660605442210980367944310075653859481690464435885881966479327232;
R3[187]<=640'd4562440480584443556346379150828043813518617890477360549214123916492835615594412473956644167637725493729154609209746396730079820470735414033314806352607537896486811262143386893048874736236937216;
R3[188]<=640'd4562440617621676529195061481580499460936096384770341798472515358561230516540013685060428881792123054744969577660090558077343053348540921949109114500754582758371846439670843345502568024425390080;
R3[189]<=640'd4562440617621676529195061481580477630879575631771090935689494973291115834453461221075212071973893776401675414959390317170521003091572504490617806304372397482827108484453385950513179835875196928;
R3[190]<=640'd4562440617621676742934902804619002159290261892763912284509815908971362243651463874283394513650642278924096751126667585938579807178321673405941872675213743359428107078954482408045190437446877184;
R3[191]<=640'd4544618583959547758562646691376032385553268132133303064652887815821980654950680032302302095534681281095806728887327675148567269526257317545641264471901150205326483352696479720084113937429168128;
R3[192]<=640'd4562440617622134035916891350241008694408560971550913611819329416933133208758255111343511514735376699669062599089466108376106725825722049573075828020045183070910647400110430168700021690537678848;
R3[193]<=640'd4562440617622194787320138661744087677511840654055780288892501321022916045327042145344094164519573393605932381612135538205775019110092264608879790693812030882562039703738323510749363773261283328;
R3[194]<=640'd4562440617622195075707386779383974602989414516821341440354219903630942832201572951665978100999078064728985181505985633249112322324382930540329426237809526787055852448681802806961823983899508736;
R3[195]<=640'd4562440617622195218633442530654256918040600365556451395601007171196672066139561514854156831792639662779882507779803156400107181864725815980530829312022554552466851888277717433166168258753593344;
R3[196]<=640'd4562440617622195216631612093736715737123478640668176877422109163849058532667776263766588795976784447846051676272209526446021785723514899947995005883748203332114291965727051056516543839062196224;
R3[197]<=640'd4562440617622195218625713455608334806406196347894386748928831351786979562525857054939273501895813436833801373090733180152986086993366373547989838957517466155269911214491613282129406823604682752;
R3[198]<=640'd4562414502645962466111021073509777378850903637324147057067896790263835930981202841951790868228571410258858624164593109356785035596657803645702594904167121406092721885331698007827324852729020416;
R3[199]<=640'd4526666013591206781011493250725113208319479918727812358899744158503749014833108054750241297799646927282450908368240415824999054069767145744263348359838600100689230514749453702015786850992259072;
R3[200]<=640'd4495330032005027655210033398919524715102402503418488847846732522694450870712021976267978961015240686618411026114863334889058080214118176256645725294462375300292608182930007118035235189797945344;
R3[201]<=640'd4419864450301033613812733829768825307249931022797455959362035323479350837559317752134060779984945195364907868116092511686859929196050214244392774812630362123472821835448428079040251872679100416;
R3[202]<=640'd3421830463216881382066785533760022339312858050889078276155643905464571864648649725010097923574270257994997890464361749261879961660244802511211810743622865517717374055612801746066430458455982080;
R3[203]<=640'd4115825162073609140728734724925594566690836600961383175362933633458990533647575814223663602911773454134224432605690398626336159080387582781045299393908825192179125545046603005952;
R3[204]<=640'd4052323107574750706291932086939016717285028617414782023783638515735653426169693198978948318044636529139391909228086300035854155900968924702467878471719550514545346054996862435328;
R3[205]<=640'd123642324774861966925589772482424810418165827769091032364668585484608730586343721906410280568262913932133186005833542196966160751661441694045739257944206310674532765953687680;
R3[206]<=640'd139234637988958717984084147370757366093948968493215588166443749445830829937768755561734969828236907381598256188136076292979403788955698689004000543431318143982720580010609967799682291728512;
R3[207]<=640'd243694609312217871120424947836452616147132117010723495985040418852376662841785535582728935995499619225510392789289049458583422022037734916308545857185339734993687348840670302028239226691584;
R3[208]<=640'd452528640388398196709169290462216974094974371932091366148603120953276349521657517076764936395450183758645764087940588530784232338150669695278498872270984447848916970926144774270564935123712;
R3[209]<=640'd267899986779229498901899569202075664615096096608044120448979515392867425227674827814007955466611241061254743844077543461115691937599909169455713781209353760017588828600121751473554979840;
R3[210]<=640'd7613331470346097347029960555930447038097236781786943160889213881554400713233568323564553220460160616732490649756569749466117975789448153627117947045225351379615177729300236069888130546688;
R3[211]<=640'd8430222076232957702020487854929452084024976878389738507339901675891493138996244190240187285032882755513848279591228690209221720422572919278777889262880638593279423247968158311183265300416;
R3[212]<=640'd78047541216451196883541841262756889389652716842131410135454497812526707911514367486323330160914184740801757222285457475829732730036762624272602378680690330553588751955573724348027741661152;
R3[213]<=640'd106601519710288509715806861835086512928123770925544577617695353796235905571427613187853398481454328213843521028592828571778453257796852912868463098995898468493689615646986442320252481044472;
R3[214]<=640'd1087770609284781733572309968262207594861910082982052990391883249706371987558959703898610781391583755407429532476010436420546118443960651247526188968661615305318317462525109220141227311103;
R3[215]<=640'd14141017920752494249590915140057312514997578080180929299227044736143029598223930322506072705801909132129240799886882995264447228462910586592488245641373916878924857207279268010215040090111;
R3[216]<=640'd8702065285935888005497020816352040459953275597411418195076161434651566718234249601495426644609140482047216656306663497187298571381418304826672312508572077055391703270121025183435597021103;
R3[217]<=640'd2175421911900102781812833585684223268639493005910494195743705230217355240559514167511334553764523867035094761750336067796449455618942422461579584706530253126417335931473293714636541001703;
R3[218]<=640'd1104983490231535982661058662687031284400053614554810707302412926399022743587633964735368140485734481263569790133555772873135715593706042331051799063947716620447564066866018799141071179432853349;
R3[219]<=640'd1131733941988280084389895842702455274338784973738481825029894224768218615027918681121129109357012182914789580515325847486552861221041484583852881997278494741306193378684782502369797572827021303;
R3[220]<=640'd4562022912646001237626101623493557838558673750657985347401455912535627999485089432649472282741494322306250741204305188430699767047128139932113799372207438871384871505987647366438672907961892787;
R3[221]<=640'd4562440608061727810250765112327902727746359331321451761688778360133907132914930961786528922034298716644924207052161002980462748499894451018234825484866578972129592411393052399449906935138090899;
R3[222]<=640'd4562440608061711474572527732466264340461304572265376360087484386993544042423639350765822461816269129279403080972791764019787102145483816321234378382767898354474266237723019613615620627363397593;
R3[223]<=640'd4562158868037973728415514991273823512150470980834880830321660457718178957746216149061793596226192203757282650695846880923359874089295273684580192166297348921187802879166538042165699443127484361;
R3[224]<=640'd4562437354310367557461020070242081616629767323844711491603492912511752662659446197902465969672880704714414008114316294954089708708645673895527618259001497558422993723437123053123107656654258155;
R3[225]<=640'd4562431915457320972292939854074980306094826019023881870492811223708059403882528574890058633238604920523817505477714125788812980171323384120933768742546563669325213787624474226012031754000952803;
R3[226]<=640'd4562162148346217301685372224640444156057039250895401964760586433785644183356988193749875594730689625405669983324901192119545729580704492701706174834552630495991826642378693901120474236809965410;
R3[227]<=640'd4560212863414371881132190237924789767126817800233568962667508198453894739353125874203716579214692509849279009348098631096707558036993632424670125784443651322178820808112349680424341476833237363;
R3[228]<=640'd4557985109206548543623088103351693923040484339819753531765965387591819702221181507646267180791861333350256215475779074353990863272709916349199856285482554632428594175940513471096797107959844946;
R3[229]<=640'd4130256301304467741875478265317291611331744167318221986308439269593634470745136311181712956169763723722902589935598893720098984292861512539727452440489978745713237276350695343008231786546443350;
R3[230]<=640'd3453019022126173139108310475279772739562097342222731025142914848560669113651990358542260022911458522278383366767389564973773225663201591728710967934944235460252244892868066384692794090944075154;
R3[231]<=640'd471745303102585406566954573753957242667437928005741981067728375426243713441225774980368725279402707700459263697997977629008199055018117710290669265229564471901803206923;
R3[232]<=640'd8911016831293350036408774165034932791663304273096457501967411328268786829240437190004705508353562684933249415054839971881510609579330671969418018299245054927581610810001671410647568626653399;
R3[233]<=640'd117936325775672748289124134073912649512350638711787893105611387201023838121188769579781939136625928366574046707507372836943562210471864225345891974989338327704129529991;
R3[234]<=640'd14742040721959067806139537262341392873759407591970626849465285200858888142888623712670559995566011252026999152999827043656743546108644850242727825242877827984487392179;
R3[235]<=640'd1842755090244890681062784106244516101853253440905090565518059191801234260303628759880400010764634309842659918845334581429796295136717089813589362191585797640724753255;
R3[236]<=640'd460463826871490421347094653622523333939342123658476330285364281609316623106078905536949927851792543900583847228395710787472393648877726711763897442216573885646149133;
R3[237]<=640'd402427838921887279747098719953010683567035057541384155085468879531439295542221971339882346338454288168397011339986722445679734008596708334522334327057397326712004416;
R3[238]<=640'd379736442470661669686602015542228479435880141276171784457419279773137731368480087601333625356456481560010802039400548383254290780721558890728681791432594529428835918;
R3[239]<=640'd1581539544131530388576008974803770780188830227687207597245519663428767260328728405426308368846448344863381939974881680748136612566404710566493409176300582595923321;
R3[240]<=640'd2702863053127904701860390860689304073927190639860867815030383840463354111618469777828112875395781338453074185353564526684540811452604687609390838347850012292275358;
R3[241]<=640'd878586838033278501305909368189896700437637327613966595481919130778080300468055356469545164115213538624244732562404856160196760061548804363556053409544237666852;
R3[242]<=640'd17215625382046291639179005088594405927210709677104666045150221217290167181612016897888460754092227597923902409441713225540846495591498261336540739711640570305;
R3[243]<=640'd26815615859882163479367870324083175804095914407813765415163507171423831846758143337104722591734777057375084748565700635377323764485246026716642475118129864;
R3[244]<=640'd3325764846644534310160072582362454386615788136161880865434793651410149504181037076610112082695047064283211914379103688757062255697579061342033255868618251;
R3[245]<=640'd1594958375650174378185208858004845977671991781648505686650652618127979211980897608874737937859022148878485972309489296068640624280755977491805079218143904;
R3[246]<=640'd628695583635149913046744168473867944262048590909061361877590661004097201323358543724906106803562241736552716676792741086301676521696707693425457507555445;
R3[247]<=640'd209496999057782208114242198769895897977859539474797287097784191611150543739565930457422833397502298795898876833484422741702342044274200463518715200826861;
R3[248]<=640'd1075682077132862549738663055125816756194600726479523483054076536798687913727174751005221398724;
R3[249]<=640'd1176564790002906685583417206192786879782052645287335293747296373786517370662806119060851621966562887019305850;
R3[250]<=640'd3421830463216646413980878704275218493669921380436419947934394388424456375406508039889212939837302219723798116670901252734469694320756363513793636314585005011410233407849489701488895149605042096;
R3[251]<=640'd4277288079020808017476098380344023117087401725545524934917992985530739699586165054522473300191728269639606005886417646113318837183225565223547540013393504702862619320803489907098194705319710494;
R3[252]<=640'd4277288079020808017476098380344023117087401725545524934917992985531162775406200510229689819115526472132685089581128548428408691740910192427299808528004387721553221059759874448725962837853586390;
R3[253]<=640'd8715361892688209479147500920655656219926210804045662801831628763788741697771535594258328130421596754478572986932882781576750295;
R3[254]<=640'd13949268845385398940843222423733410478979213862550638564478225650945080925544770143237653096250854228484637010582171974737233078753616930468134956105020098578008;
R3[255]<=640'd17822033662586700072817076585215720754836715731799503541084893908597645546792505319939153463116916052022162851995384445853715659950413639900544870238642583481939655891202970439518695365056210;
R3[256]<=640'd2281220308811097609320585802850369647064668995158060394749232106030187054560896582047980972324792487342005405609735556083430380433303848010173002167657376018602015447979974455108263951088685381;
R3[257]<=640'd2209932174160750809029317496511527610309015768373865536950698693411706522158015143800435032441617083505092739105892272515834822838631916394006488721627558115783224431179103267635637749488503736;
R3[258]<=640'd1069322019755202004369024595433321917342435580026259442266061740694863675912068115476994397730846090802058331248686981820776888942076917075266270316718546195997339707326800425047017885457519303;
R3[259]<=640'd142576269300693600582538500069647452734253045749886279507666087329564416291663880261668510473784709326292179509589157528021711015367637401360218130853779253611691955429639495844926696360167151;
R3[260]<=640'd15220364604047040013055708075522894121337819770528768128042282385730318812380181477508403067890273006064893355032922550368032886072057208573718630517199910693009724605507789;
R3[261]<=640'd15224164365043124983070409968034915698287709520248036816427236241239416022509445598258437132666882019718160358520163836977023235969166361932766292706650574001881762378160682;
R3[262]<=640'd852915501711189033193742149666645947526286657807553028078733150284661305060413391177765746223899052481941346210614743763029968995178593296692354300218220971653343913551973;
R3[263]<=640'd33965655524914559709860641795994246996522331748886736783008639278833914169443301489439317911221172910085440811011176337480091444067305487584807475522337595360613545319072;
R3[264]<=640'd60383398797144661609677748444838150270411567978606229742097861770569966112623228846244615518691156328494575575588720819229952882637834311969865783864128702792107789817707;
R3[265]<=640'd120766740008192753105722484185147511153567212128686400643168378185554701658381505907399088772171886223225286167958179440871301184616000609482253354039553470055515004018147;
R3[266]<=640'd4084679388177375574335039119201169509096119567912951842067823154896768523547524321225897057496117438474402666698943142435838309207781355080173127951202643583501359264354592481435370;
R3[267]<=640'd1013065324433836574614494317165643268730223003118486418791496478328286402758946682742323150330752104268636821347320696857211477967496645732566385590860356412442923131194635216316023;
R3[268]<=640'd3421830464278663054891357862628926509344543164177486745376865084045435201720053991603535826568232541254913084334913145124632238729884987454868016555043902532728169908763994127239560661610646314;
R3[269]<=640'd3421830464278403710168303013407232407138231755045769238180823330753883220911055698812292807277373503864586319770268403396954464110016215508818669560818865129474460508302690864355921872365813619;
R3[270]<=640'd4236138669195691310674125260640264411451553582756493875510761682071160956527641615770959456709141872200123346865280874398062544086167404621643680748030394560939297083880311041307185099;
R3[271]<=640'd7967073881196462972168936565371181625946378271573036403004593566461191549987707443656974263617856504625431963920851300748618067499730641379421360093148416484627274301447659486219587937;
R3[272]<=640'd50989267065183498125662021309397550352047359784509027974802312325954596905776451479521178662576493122174596965758072908162113357684247594099655541328380264921869506430839731282397276659;
R3[273]<=640'd3225536676471225659868121018513047111185087166127766655283337088804914810978754239765598787325983612190396481300110305556987263704899175206340452962414114995828583887365465934791840;
R3[274]<=640'd8282252370854373529094368533295871254050403085106984364152643209886016184161687411302229131748805579583827679471598052389402095847660196857721599038886801083099537955564675396641208;
R3[275]<=640'd32280392369106063028278136030174817937927150424943232174887473782944912478625130165048036524635906458512416136892234586378895168009025365901421746475569557579205094419919239234403938;
R3[276]<=640'd56826630144057355482797300707960220134739675023588134790296933769170590634255957962985326420975827944609663512469858474216921160160761118261892933858199659941848413945435681381932;
R3[277]<=640'd129672358568744488893424325582969994450173735716884552422536432447716818172438882661326025481043416872253427570004344955042045951035234674695702039999199943577569383764903542537116;
R3[278]<=640'd259344722088927679152710905306859599199892445579786675435605258111911713691460972260929316316834885141372315618724511145860824836270116534156923241264347892508397977271558604684221;
R3[279]<=640'd1062267817794355949575043599069683101830380988196953447600710556714043928202590387731939955279461463954328449220190691363163571453481515935812507142586941231254036128629841246321727516;
R3[280]<=640'd531137992816767098689588206552468627329571776253520896823909216979105978330075145774704150341048349929401821610069799704533836969507413087881584486307903663431133235510640906497923326;
R3[281]<=640'd531137992816767098689588206552468627329580923117651181225789741505088978302314143428421840466368077669391615407776673648884664924336202370657333965788077126794363001783488047505391439;
R3[282]<=640'd531137992816767098689588206552468627329593117633996566490124145665648975885241881017499571917818193370204986720976962724630914187162189070746686565000133037396030970483243270775410323;
R3[283]<=640'd531137992816767098689588206552468627329593117633996566490134660587152545777018959920367968182170463932193387319121209169530747704279041647302597503031760123332039985522752011680050695;
R3[284]<=640'd591747474947310671155095576680210787699992579689914363328172739116828547778040423704292412904047489441873376582575940650145980530453409084165547941843606940067159691430584302460880050697187;
R3[285]<=640'd887621082748605468523219303925706683211286978984686974459180743090943964072941467340821132108052618520047787182107408928053847913852363023199724244533933064742562119598464444507441052251135;
R3[286]<=640'd17817682845718539546484949038136515957083235337238305872739933007530476949622467674016576504041498397885010696269135317424000806414675267658576769261201251177910435952486863430120493163077433;
R3[287]<=640'd4277283864175266020020786729116810019972609551534365223560604561388281629029242486398303925024007963989334687285310931927574715119429334873906312832473870106470918238756475792532609406299200595;
R3[288]<=640'd4562438578185087300459704412353975215051816718443386138161847745570595348441033572885451647546314081397943736530378146624756206895069120800121664133706012430140431382433850050522717854317594233;
R3[289]<=640'd4562438442346545637571518922491791389257965278899946279473435860532955412501856722894995836371565653169008542460836333389304221392342868374591740849445839371794193547046087667912607463110502093;
R3[290]<=640'd4562440617091057225824404507010703118340759879918966812805643082737924518896007584063427248822737597537687080770422277780208923912557949121221275910697642543811528392302853104164006081871869791;
R3[291]<=640'd4562440617622195218641171605700291324893228507248364821248280266820757120878625401731886775352260205765018844986324890406351357064657409363641592710194478382103547042604026504298147574185152510;
R3[292]<=640'd4562440617622195218641171605700291324893228507248267266606448430397195781208711371506883927478240087162091541212614054596726741409399355865181410506626069950570201141204111471725599430420919149;
R3[293]<=640'd4562440617622195218641171605700291324893228507248559787630912239727758917992128447430708819476139961634913070489825882616077271685027809592140853187437005819861572708631502718105466327037392439;
R3[294]<=640'd4562440617622195218641171605700291324893228507248559216021771463780238332125996508770684490953884191883208051202827596521499060771043731458224986062978416228525067419467655847910780145441530841;
R3[295]<=640'd4562440617622195218641171605700291324893228507248520394228204163425282800312517901596802978128240900013446295562563284147556246491064801668684429894201542457610536545383583909193818390342745587;
R3[296]<=640'd4562440617622195218641171605700291324893228507248541734351941630400206440937856103200984006114308406330001457660029809148433025263764071652395918158981650187631326409373096515663336640320481105;
R3[297]<=640'd4562440617622195218641171605700291324893228507248556977264807685302492818557880450358091230182245653243234683846461808146845201342036842842802708207106797696387732328359562762428418282130370414;
R3[298]<=640'd4562440617622195218641171605700291324893228507248558501556110615578713016158666002726509506652331449557143984895965668629436729195829994542070823787605130785380189579580168898882866663291624304;
R3[299]<=640'd4562440617622195218641171605700291324893228507248559644774576705277916092310117560908317696823606888487794184210617384835885357368837966903249770484895175183567223209202888990672202969191316487;
R3[300]<=640'd4562440617622195218641171605700291324893228507248559835310987247025488809127707239009382484516890971770489512358111020305935933122082681137297612884958586531174072536505094435111088623658542486;
R3[301]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167127982077815696917890623925653548188500791101284775469945417144793305361530179223303278336839764138067038757122723768799;
R3[302]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167191025287729928084630270389813777970588918684117520184614133646864411365343512196592725134614229575835935634107721055999;
R3[303]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167169590413586111526147993464728361880145590487469268295385683805024804853944160690905774469124774260156955096302962760852;
R3[304]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167129856133330505325547752722139483138020114090351128052670440806515802227653235631407698577573097016518746615330233754379;
R3[305]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166242196010206195883737449044438066437180415390609749924678928209045080651479372831379246201623645166624689145178227595539;
R3[306]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275156978636605530247760675221571929239817503524103231854887947758217717324412757708295262473360532527777749833065804118735053;
R3[307]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275138838001593168989612917837004801485833086524462461773617933272801550427099199630534324314315185160804918709793957556845006;
R3[308]<=640'd4562440617622195218641171605700291324893228507248559930579192517899259028026595736441771465373479112082919510322780759596352508783579576295530383560859264680852916064965942215790850024722778523;
R3[309]<=640'd4562440617622195218641171605700291324893228507248559930579192517899233189579704960553651186040964565199520284260543380792384323341241490061264458017814547032587711258055330552817108418100260003;
R3[310]<=640'd4562440617622195218641171605700291324893228507248559930579192517899190588513750690630183909510565000258383648315537679875621958970694348601544318845827307361541463427198595508839009752832402877;
R3[311]<=640'd4562440617622195218641171605700291324893228507248559930579192517899272525727497070122567882549075701038495371368583849895593103483588051673530940566683936197539954304097108513271310354701654450;
R3[312]<=640'd4562440617622195218641171605700291324893228507248559930579192517899270038937331684499635986506962623190620995331099579090480014702836240975146485902282881793816323701470178118892205318988667151;
R3[313]<=640'd4562423213292446598816881745273939013601248171141278251197133118513753950164989734468108339973158330756657851362897277652723342632993457007302672475516993022100107964242184417010711787026053464;
R3[314]<=640'd4562440617622195218641171605700291324893228507248559930579192517888444767071110564268561984375568527485535912432471910362937866987029049136921426924803869659232482174164543314211658751578914446;
R3[315]<=640'd4562440617621157839748951357460663222927305716960806771387029273238736259924085765790933468632703414427401911404286290723731867694387444573925108813876941686134868279153766960159395002730399868;
R3[316]<=640'd4562440617622195218641171605700291324886524603283930073277096317743647029867106589862860043587178329323344861177631100654387964933738453963799084570292946161409572136625941675047352496012817406;
R3[317]<=640'd4562440617622130382460407840185314568520358333654742989987707741034403795518925433060360455114647136024294534640199682438939119560847007149150136020766726840332004589517665059645039693965114098;
R3[318]<=640'd4562440348931741932612086249243987481396064357689830814159788975563456055219355206317643362028316872755806871434451803533409782241302519992991019174432802934254023907802103387730479693238204910;
R3[319]<=640'd142576286297109370719083770744956713581909465398497265095621308566544112098000968000521523918959750380469011277044230854640474041119351539552627562735054369877848131874200291097244572400861128;
R3[320]<=640'd4562440617622195218641171605700291324893228507248559930579192517888742603773871451308198965602847911879071092519439958104753097029428320839601854902515844109233806371321058205827856402890061050;
R3[321]<=640'd4562440617622195218641171605700291324893228507248559930579192517899232861896152179001549195842722650688285829077925515196030506661064606780179538535085437069904979461662611342638176186967942766;
R3[322]<=640'd4562440617622195218641171605700291324893228507248559930579192517899264590883082934850569390243180616785664596841425098013639025267815759959785839521658591709144023595728254149273864293170083796;
R3[323]<=640'd4562440617622195218641171605700291324893228507248559930579192517899100649047583324523437724218581889572405604377603629613670573235478965571189236396772294088558095624480163267355475693037188026;
R3[324]<=640'd4562440617622195218641171605700291324893228507248559930579192517899273854133974404540222732545216432153720552448063035052592442897861661385841332110349950783847053722184253301836908594040279527;
R3[325]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275149132920852021354190660165958427005165900636488845544521874615511159028239082771233629201443767710984350940421170215301510;
R3[326]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677232591760884165219200747331679668106307012554931400986101423995312441223859023583809169627464812101039234551667006;
R3[327]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677232591826106651432905103721951617677666015989404619475973159315115174139714351244907313966958642650977313406978855;
R3[328]<=640'd499016942552431592962236314388230963928876041007369649286548278799482074734922050224622401444765731629114512365416471603756108690893228076476479852534213249610766341734635393998671973516586551;
R3[329]<=640'd3421830463216646413987698254779973694884492265464090000108945239624473745122060312690352112480110579190347852812423697169660106518934140108665949363674618288149241631944478463741970542965438599;
R3[330]<=640'd4562440617622195218641167831737866503351876265693978942310301612068733527251272036576017543434609786941450549724508267331635582178062909841351489129176005596474033730216948125771191810600385503;
R3[331]<=640'd3484220634285086086888400138083347423069629063144507324156838459971536507012447152268361681480097743620636461277249009407741188028155795684385601491995984989163345981636063121831398169608330844;
R3[332]<=640'd4508957112304686498598430515519638724637655649571959189510658206194622650783093375538656306661698734847013503943900983594974601038062315619395750380737194938129589186580138851148423999967099941;
R3[333]<=640'd4558542047758504378000242870197373595489633219217463748997887055542671782666384815496935590897544544334495520490706814433342092838360466566868549474765358630166139569054912697630219757503392631;
R3[334]<=640'd1138399804527474086975480627278329297141804441187366701123254407513708837173280255027638439466316016724095210368725725508793710090076722690968472449532368190953868524490605272950266642210123830;
R3[335]<=640'd3706562034592238873145940930569090172100973782544579323542032198155882750305190101708912924735968895953828570899338564632661708130609246384445842271863893711351905209004313076321657474960538611;
R3[336]<=640'd141470278533699053577827168495614554060091636180219756871105076171792532840460417023931350865997975637121750374059985514647832082045662085079305167277651967208934010394018276976023335935569615;
R3[337]<=640'd17817835547891476345669034079582172275833760752437172768504002366575707632171755864912111578790577658111394620511593861204131902884029858565471593190286740182463427538291628694797003107748187;
R3[338]<=640'd17822000197764300361975956124995499282191689393122601434534325232077841961633652832726148392460220370580673486075370135808591549122068876890046734563373715058914863074991582815592116235499387;
R3[339]<=640'd4455491950368897698424209768957287620438596246723272269216623510492726692966868323840155565764550285488474644873749214612255418463375740121721420970106742636264484067082370951265389711420389;
R3[340]<=640'd2299059203449266277664950780412529433551053005414241897146823196076848799037255372048440882291528591623380035200333597703519401780174359129021179239989856781921505695510679300178382032650203055;
R3[341]<=640'd2281445511319662901485847595159863370907380954748288809990760094804859961839061195902807850420921184570605770844220062143418997583071899781524177954878321185351716432302944564604194967877597247;
R3[342]<=640'd3136955867002348255771481345669086366486901665493519037170477432375495395837226647758031490561478222772089928318355576457595534367038658614760921451875576594685936887174988167713775177887985406;
R3[343]<=640'd445603029009495513325974207941334382237696804628685652339208532680312063506098908957442326799975320655102754037567856710354522465507414670913326098717973837521822771688998102170729563372199039;
R3[344]<=640'd35678332165751785493366233095206174627536784753921553001776596339062833196612114353533905864957229511403526368589841049816605828152966650207755840936201075859251837100161626509629237823421237;
R3[345]<=640'd34536953345017452904246022976855947245542623008072005462815554076474783332959152018835820375510447258737975681608918121891768599157832672305078680598505705679613187847295670374080789113283;
R3[346]<=640'd17856298486695050017391715141878188407375971366645916059873883756790076285981201013994266174463016666272584207620210551511693681166815080266053202986330803313039932959784960928682841802279282;
R3[347]<=640'd68529548440291814303109549278360705815414502006399269337049459030583492796056403476830500107011811441657360514072405557496532680079618031493095477683942324471401791091907907455909887613588;
R3[348]<=640'd1740432169855969980646255823169093578029020060463450275110351191676335514721547689908136706399389843401865029674030325129962861189822068427429640577742918954810598345216476460744340232359313;
R3[349]<=640'd35776775339490433089799091820415890356022212190076199626164507318590668549367925685632712596831989236287961540734960468368405316112443753159339687810015942755785856309870582881470044359922033;
R3[350]<=640'd178220338750402778659393250292431438181904140923051755403422298765142964127353719941638354695693795557616373120676413136719982547228525081379730338083867088603937074644640395761854178741993275;
R3[351]<=640'd1062146321093830612936153790022589133119559481370335185571254016127296085481004867674446765932428275458576809044986915982811347758048304250959475366561179867500300270670895997125014877;
R3[352]<=640'd66335596565985771575564055992344871777480030185748333326275164651573261391079961460671515292677204342938865056413302745994012247148533509864900618747011280536541734409311715145842224;
R3[353]<=640'd71288134666943853335089067170065449525631945109723257220879412162096792739592382781923912736723038179687278400670555334676904566858029064966131246171937711842139797809921584576571668921085293;
R3[354]<=640'd71288134658645800020001573933324671167366524178056500590252884703117037559923046865077902912604659518632006351864333668522342604659320743881158969067351513920495323706779088775061530279545596;
R3[355]<=640'd71288134651384179179669201813593348940400669219699437215859992487007095517902943136550380141780581460331412850609412669666581393100363249391411622210514106456807182496627507990543742636817265;
R3[356]<=640'd56730790582451840716079064769613337584049624843000234626311662063887816033243371213609728566841090179622857376145977189546622050842476986738123506445857885929196199220922058880395;
R3[357]<=640'd35644067325290661962276570445632652274715949935039466309490241264652882118805569346035670490128610684537043851148188874362775749573341668026324404817408392559040507612510420472399102924427362;
R3[358]<=640'd213864403951040413720486255937416195066955661656020720175798787087015133501295933677170168397512362262275948073245917418918687446452582741669549252022421958222117913308341559794846022879163950;
R3[359]<=640'd106932201975520200759983833182806954937867587079622122938289005742597408807671693069633131114146553618047217584389188444180033140571666474727560096726471201455990039174739718025216906188498071;
R3[360]<=640'd411245275974223895274344472627318854775516890613751695549415981667573579168812299460349554631033055273425827958825055026456315654843779618975260598029237953378237390416744973944811209756430;
R3[361]<=640'd231303219427257832217849180888900013339768806481513530666379633936323893509588448075394271942252393955620847161035036512234943652438252586006529952393959484284078456145345766882762782626011981;
R3[362]<=640'd470060557184393446331195042332930003698552090691392811809220449677808207730540911752331497393020316192766154894140034457194289913554786297820055048272625048291783167601551640528878043804582152;
R3[363]<=640'd458918293647404992133626935389165352214438086499027418705714212129365475830031052879685180822990501290223769410032773776083308032169982109637909098227290513336574340642659952199482767473120008;
R3[364]<=640'd258419517851234748794805137096057630911321544305883236804750947922555562267417294955134757406453142100567221486092460689748488452099515813003730846764874857951020085696494401858315165608934148;
R3[365]<=640'd374263668274865734046772422614476959190057303801967137344097857070365028330008917519917718073490715877472655949615468934760187269188032328207698913940849333391831468188390784159015274423452463;
R3[366]<=640'd499016944647997800504543353937212091630447966582062320792251117739475136277137612222718364870194324680849033832328593885202581553129283570130211956941132887354007577640564770446860556099131004;
R3[367]<=640'd142576329051480944232485304990109246840713213055940830612321565020753285304418272803125591575664216847261325578250724275011139749012444747637721868715765770446207715424394766247183976687600270;
R3[368]<=640'd8526645388524124685744876700146187841185754251975785695759493931016432796324854940266769623866988175169520687703583342178299701500922852788956710415774747694606974185138456011341111877;
R3[369]<=640'd531287279474491451649388210394964980656205536865553805724417114062469549830970439463278449992660858981391694354521390484087425098526651960547845954786749817934836115332554532867289202;
R3[370]<=640'd464762396628565381477039131596685529821144278454743555327336103312236025120161933172044395065312507331777303110870908336294348086879818816798294976238648759617462712985949341986850077;
R3[371]<=640'd74691350962887196629356823997491366849415173977484943523209284336557883634868102105654569338580415551678126101718617254859708534087466789364307368450008880022140074679942032771385108;
R3[372]<=640'd45644675831197537731182858687191762847733938774619198709127088680003785036271673802784848777430161805136831717243123303433218902906229696113540284753661329829218339717486108798227447;
R3[373]<=640'd9077065313467448978961680858355153310873317661489553347095883871646001310411451481260565727154241419010422201125582677242978289510476041408798518988442344417076186249364172591924153;
R3[374]<=640'd3128345722466222807164152595328348451780681988753549653352898770110385384022017398008338612596155691396982334599273778200513191474731842068566458025368285626336823592838547918750354;
R3[375]<=640'd454803014094291750085653260554969284630533305981053127286938108545696177591855546575586375249726605009336872822734107764506102487959473533008596116625661008312500260483751164314189;
R3[376]<=640'd48128022823254395307350860674686545968995665680258597830381552014041463270986259923013636715727086825179758429773828167637156672933142195819312458922885498608548688628656036053446;
R3[377]<=640'd16205117854683949986486109895364879774070812354375379863633219495633881654958007074339137061971122047674017629885258173003588066974581937596918977097435099736227195719816270839909;
R3[378]<=640'd16209014501079269023045936948692784696018091442143927696157722258947373111094753383040235447053594768383800464904531665590198820881406525362924945577132778553683271145113664880680;
R3[379]<=640'd3106469601794152930646795325957835934167271308483352991759210317734725237913218818724218903988625819301132387912800107042727306372359155018806073392238478758698813431939814391808;
R3[380]<=640'd1804584437516712589437316977264940690319801198253536924235258604601146371358878572704912504270114057585547541874266654209708491133312706087080365550463297319306235190839856857088;
R3[381]<=640'd229460889404312808392196162456181655365638289713273497210800701492168545017391134237592054039335308913223586089409025500764475075786566309643553014948487889703226914818848980992;
R3[382]<=640'd57132843447015892986951974161821200830045119727953050562086048828240626512328868132133048971605264487637794424281710987259922076768427283563753565456353216182105802781220667392;
R3[383]<=640'd11995500209710123047698053171741527716092147263825591377233010638887802944254883282946563065975452893662071947824144582357822729151353483433983433220176305086820078466568814592;
R3[384]<=640'd6693378986410719298568317425559783370841799008020547857531491370239626478080956294593807866947852648802361817473958370568605579713546397480185807203482859448547632425881042944;
R3[385]<=640'd3207581239953935788684968812768870575024376018947567594926060718978366231763845107020742461826068153121502732069596347819392532878578339622694327204580879979088640368567123968;
R3[386]<=640'd509998304177008764063906912009155223242904177135202192451228170183026121657874032396516652966249436405942668959439187913160837866474543790965200423100000960444488854330671104;
R3[387]<=640'd193223102649126856220410811882338784588844368082080256855861655208800868945697063569734814018263405691719497979686517418021826638345228750608237187555812157315894146439839744;
R3[388]<=640'd46495215288633272001432614114006149830774603042923258714052763411096635268581867055159239946648348264829898325391882174315395470516892903284057998956605465339320867148005376;
R3[389]<=640'd24160907443693475674990976671498277965775926614417220967247687131004861437852281899551051726682121749029801195292124862548092176839587603376604369370813178078470931551879168;
R3[390]<=640'd522129892458594741134800313801006199464966823652683684171214811739944075138382356426180125051138403210550730050026020642152548578931397605471349268712681651229622922028542075628414660771840;
R3[391]<=640'd469916903212735257999562205776807079254597814693219598673871163566869001349308359887557998969180320492093831826579721523910495060825722155462311020916869028611625084278470767613189292032000;
R3[392]<=640'd469916903212735256324379982643836331920396218247843396929599644768695554062902821191533875293569569248750054288735590900214184429158085722764292171866635569765895606179792371141773499564032;
R3[393]<=640'd261064946229297364530943515302362660156130281209135913466236683030484118648730362680800715951269909867563988465256616893361952106086695277939226922071606685050382988851810683144094644961280;
R3[394]<=640'd45405485423633740436360351093174408326335552007209148790142007922252403097372771600729200944845281902606350066609283442294385168581084038559000948478957484386805109227520;
R3[395]<=640'd14860164191335011685993552402861117394842160677650147201684088463860645469396325677491329950340966401105922429006197672644459994946689136962529424508481304043252399210496;
R3[396]<=640'd7544239339462606139234171341734304843033334667214307631475034636065383957723039807865529192553123214725432755716209862731984177901357148336083905410735864498106092486656;
R3[397]<=640'd2888979292735292954068738726472050505754780710796886803840710777455792227602284107950437378187208900324099030461935030534009817920407300052832287604824830743489877639168;
R3[398]<=640'd709431916709715009322028764354822640494197501151113226025314281695251440681195915982459351550411662962073008155433887173444123330645070500817977960778213885993770024960;
R3[399]<=640'd29663363107144764085900618320500534113384935207806039256376398194794970492335761136324047435756942235027600244180429855919665197060317602317008644808827061299998359552;
R3[400]<=640'd14742043522797009825337538451613453704831825621954287411892209321731793522204517665928569867177736032307910882273329227986138574179868667622471896544456004947582910464;
R3[401]<=640'd4376543339331627987631232683434781868572910429657338187590096932831211664100232294973304342833547300944726338026470238693376078900573840135446218066307731101478551552;
R3[402]<=640'd4139000690979740678557586628190872208610867940888148299937806959396574591603947050278081976621871306739408554081608949387781813418755888096928302653692534437219139584;
R3[403]<=640'd948595973592827671695600049592566283743763283230086720412383243522669654432403753566140244794533088184835482197979807201092450668387571584857559198969038284213190656;
R3[404]<=640'd288379595075684412167419728059830886919180180973071225541612128371173194855752460787139286974721180063829452660083783572426189310107358575879923792400937379206004736;
R3[405]<=640'd61185282429947476590299795912493412718232194586227876018805946310719988461207952603655906689247059370680298699989991356977468523762921510437680058120492758247407616;
R3[406]<=640'd43189572427614688471554225683816331831703819537954764743577099245427903923934569887355292847065069229942335919101090710487422188380617897443921170122190969821462528;
R3[407]<=640'd13496741383629589148575128113830723819515793644369670245081720314457755048604248554996405655764904230634702005717380524026473253032507019389710987600244814804680704;
R3[408]<=640'd3346067134691502309716957570220021516128783749106390715371803915266864715665136957846817107871610473954081105552436469414955173151470811098658554919790333772431360;
R3[409]<=640'd702076606316320714132550842599600218887766143497329527444453969518651384893755095569726240183729704597221493927968369215130620062144350536503969207017649993678848;
R3[410]<=640'd118210052481687043729087998726749340496880161537118888915356799052217278620616961885959714651310471257561383606801165559747151809119552222597223425556343643176960;
R3[411]<=640'd52374252930446008956922670158157567637928333741739163835190276847303529488745142994907369497303433609178443289462311579203877192854196630571777808924672;
R3[412]<=640'd7029552803973744348147403231680230073964275045596893218037097096976451721870298932914097318780413779163323557703103513220930784801441604992983153123640639225856;
R3[413]<=640'd5272164602980308261106125965825603944130747746969126946370310882836911866876318399672398888982214380523493995808946977321430571809663032942403056938978792964096;
R3[414]<=640'd1371243332703074538241961397164672889299781979306500898878699117527797459227384358957171158487330848343583550747509918713936351177661000261672318798712147017728;
R3[415]<=640'd221588916891747808166882537296490585001090449808682999196129014634839874820895080706857796475995998892292053458308126195779537612913867592368069459456169082880;
R3[416]<=640'd13729595320261219429965095972569977045683338883705095091665785949445551752766280086154918744717751607191680780711391096113002037377057423275322224486440239104;
R3[417]<=640'd13729595320261219429963801616710430384468789972840561175736403179862160933258261388209226383122431197914340832386577336580035033965850358017606542244565745664;
R3[418]<=640'd12013395905228567001218326403937777518463353289209321972903764055383718485292787730276638271970576612414852285367157121881317599843601391785821362020887298048;
R3[419]<=640'd1689383799272274112806113794281407874979228862056572497463020615237600536358659911888530151321833995198745427568622745334968524445036908867560053605933252608;
R3[420]<=640'd690500625936092176569672879785562613609398310051160892100517343570127032614829212115657727010817881545345781109292215084805089453162389562673356479693586432;
R3[421]<=640'd120676818150699166179906251623184054169446734876295781112554890184796957775540880309996936579726719038096558888298354466513957049352387425901361346746777600;
R3[422]<=640'd55307207711013213035742853225906525202447144943035221446508070578963049576030323127388757346004462509691841254335931630598548601663930712157825471304695808;
R3[423]<=640'd6730091089834467684747118217046252221156957446492345175288372215223173461719458754162579690851136850348041028489092182938445045847580671578298784218611712;
R3[424]<=640'd5047568317394142258972346286258122559398532057804413553249522628059844768657140147733278547514964703348639886713983382146311405598860322904840030503567360;
R3[425]<=640'd1515579851455913685816106829800408735486612262368437517421002715802873761747495403522503985417916877330149708717647808978711211516688309769102238240735232;
R3[426]<=640'd351889490348835251026417892535889654871016978757027733073568966997005970808336164193811347724748067419789529216854022296484520059601049068414675611287552;
R3[427]<=640'd157122749179014809760633105542275250760453087878049717292550645047043728940440234297855820754693010293580902714674268406771588148078897067282243002564608;
R3[428]<=640'd13093562431584567480052764207969025726198118635350042592867560455090604635529442477476148739106370621294016013812279906857920480104875447514549255667712;
R3[429]<=640'd3273394900300398554502507849498531929249194718238266971119007940478510093592196024051994405480111764046559217928710842170451674237350250823276633784320;
R3[430]<=640'd409773500469770133720267997754808414721813349047946088874108865471151225494541352292091192763909817945234899453589159220684770803533513003521221328896;
R3[431]<=640'd383500565909219013640766456488203668255071590404510643638052142098046238625204340761329858511130319864475490954746629457961297262689799034099550126080;
R3[432]<=640'd153440184745131652996082034185064182372382034495794432657254834348916254979525216119791785370420557962323839794287691277021803990719059010194820300800;
R3[433]<=640'd38360046186282912539217066772599590041887039938668417927506743326390996477510158349844623414035940548384157654182452214582388176638846832597845147648;
R3[434]<=640'd9590011546614338458262004404811504875534902952911272546598553925757750979533808808948699920497020586503352887194997131655783322556446784181919285248;
R3[435]<=640'd399595984348940541129274665536496944798883826048374068192661829024044494421725123329508213942210072988404531874110074963385751076971010139898249216;
R3[436]<=640'd390607263067004205104365443224203529991550810717412606187965603536048457444188413168104120218477233093283158519044540398925557013668014631793197056;
R3[437]<=640'd79580199372508502486992238623130270577627094749835083510460620088531293566986185761665050781016118244253082898946370548712757612263217017548439552;
R3[438]<=640'd18730491301983957924380978042402016701870561624123816031872110474242809968495143075491371394164792566339208356817749225249280013116205478046597120;
R3[439]<=640'd3121748718941866464520700908632237664062410578511609686710633944619472550863956583379631415173970175282738200716130783590263968351705217613430784;
R3[440]<=640'd792821910411161375401710091386029434152926061052325721791137985555663177908032447544965700834321793673141516410437209764189354221685682003247104;
R3[441]<=640'd588233370633135951652027467127184360695257806646864236041471596232056450546202403120051145062452415153904050419972061744027951695055959829250048;
R3[442]<=640'd103627990283392961111002575277939351819357186474456977330041225626062400362362244433589775950365164318342817667495904467123108142599527267827712;
R3[443]<=640'd48586784688145631042621294775223231608812637823402348275084242849567172875980030670993484258608795315121817225404018573099358554275966944804864;
R3[444]<=640'd571081155381527806391094402930219648258344682302901999810659621007343796146032717209434619724421295952101376;
R3[445]<=640'd165131900351285148835979104461750259737352679220116240909106396435912892257078256335195475761118132345765888;
R3[446]<=640'd10889035741470030830827987437816582766592;
R3[447]<=640'd10705681053419654637621553834719515669444952064;
R3[448]<=640'd63461373003863865499383869571146019823526849564570997051326284384909469020901713220445338839850804645665695462538254405861376;
R3[449]<=640'd338460656020607282663380637712778772392143197677711984273740183199779021644099438080675751477411619920270347574559030957309952;
R3[450]<=640'd1163458505070837534155370942137677030098031095394983079025188935057018463680147558743138138901862431422158165571929932109447168;
R3[451]<=640'd1163458505070837534155370942137677030098003898030488300315407396456403806244693486316850124782145682848434403476265944664244224;
R3[452]<=640'd5546354770209691541004818510199305743190050580345496285459450222163196021940436015848736747254064472635858127143822660325022367744;
R3[453]<=640'd174678190729611336153440093601014273316495535748920789628898590324979341869980958584951918336040515891998104029680519681407295946752;
R3[454]<=640'd1402970865225132318946677577176400353938837160140895667424254002194632395786773893409459445097816426171774398253060115325735642595328;
R3[455]<=640'd1073023171624755350656846289263373393229901148172869398412642478560590179420966499750071187930454501845137527762852575753974228975616;
R3[456]<=640'd1219974665413158538214502241022956829512602711088834192295282414474086658176702336621160810652260393942675010696128487402258372231168;
R3[457]<=640'd1064705162542392907156124701167464459122748287728628411299250760507139766362796510947812699420547888067955640381838785516357038374912;
R3[458]<=640'd1401931883190940351505720810237563696595019244626009980214269261077823904892516486606360838325633411219894405431296;
R3[459]<=640'd214524926879081553593184399971293538039670483515886484243540299264981597830038453502756058014645682709327195053105412205001223251702251252622696209407016960;
R3[460]<=640'd80695308690215893426747474125094121072803306146062350612546095913931595261107541378962009056710733025324155366782533632;
R3[461]<=640'd1716199415032652440654000858629571599077480093472892643198675918297404895501351303555393262215153032460717108935221912092361365476108262553930690508001116160;
R3[462]<=640'd1716199415032652488288103494066464778117965167221166980593380092587527737393441559690584160333627591770726891963151354974694903637894755759148314372746511104;
R3[463]<=640'd53588365464909827791036745909669456058868634893121448231660204344346409628518241867115975594341354798173066729643171151645694029861759221760;
R3[464]<=640'd339392981277487863901329194949383054071841639425493222622460898235483065511860176677856654132772994164893258495825227743205583366813418258432;
R3[465]<=640'd7198262071269114212496861612297570974191515773237147306420848927707430104926954804397048082178988335188486962784373377238773490864088855067695820683930757404557312;
R3[466]<=640'd69617318994479297160149380949995777077803420585545727035212258343154492874598479367223886330726055041430859851797464709449696817295921854057917151896664329094100618773458357004066178990080;
R3[467]<=640'd482835233594231822758482976194186673946812262130367920790159686006231917958257019115808187878012311577954789791083957830083480234146287835807512482869317455587754551279616;
R3[468]<=640'd30914721637584206457085304206284713755024124682316348496196636151225429795767701085217347729582777089688197578208059348032971824887586041190329666158977963081740879197634560;
R3[469]<=640'd1013096237055811767763593764210089830803740551477237824103440997960691907929217102142802011094347063169061264181140223954726963759269335669717208950676978593773259137090920120320;
R3[470]<=640'd61832194950571576617664451745928656252294167522566765476596388007617661640109938029287938499763820724138468678519501749110506289043519779620703085143083606351840348741828608;
R3[471]<=640'd16462311521643510289668048840000694124447369309825497403985786469377359636906687895424763940799314907966521807144673943217875086988085518501643324076871473000698649098883383168512;
R3[472]<=640'd1122788120747111620156354503341614700940841369990798539610220263803827289325552888781502945262304136321462558785192170055829599984373999450673328623899126904578484227784599531669970571682646016;
R3[473]<=640'd4517885534295631582049829336335397375136659531693378048079718077353640320589089731542212140442953831254865188703142480897834156027435027551322828627616260356907585707584017310080300687057485824;
R3[474]<=640'd4259466265548115464256960884237544649968162668154570375731074448420287197134583731089066696845676103844354236566548954419561263288811729540057678585697833159520201418816931130892065240749441024;
R3[475]<=640'd4562440617389822346783835661878037424588614236539291842282921967878891429784663618674431864408778590011048051971713766547751747132544926983698972384085681332690312543324541310505750790032850944;
R3[476]<=640'd4562440430429200248146243994891093552003536816173169614991334339911054368543007670697502471801336970573907158754941956239081857228827430590047311822647676890254286357193576596989193451355504640;
R3[477]<=640'd17822041911823651008230252553153166293721739229118205742969639887893848950592828410301346630969846477379361920249545943070996069294316424088901660623114150062801266100091575864628780151603212;
R3[478]<=640'd1087654422852810333330607387902336311171782742163248581353116224755213234473880203966309404919433608180168274379537081546529924909599579842441879776749584028385359012772501273814139273227;
R3[479]<=640'd4277349401831636704867562760956837875914081350402813747628289820661427560811942579126848387114610217189390027188376928881740806508564570139255516675056981165905327941095732327218944494119684608;
R4[0]<=640'd66392249102095887336240703135882420882580652441344090113697248871102450621428757177690276346494428904551249654578286751713208453402189090262826364165889787769896304005817099146493952;
R4[1]<=640'd230428741772359047248403483563278983219156451436705705083707148028259375077303942979117676605204448209270685309948297988643650694286992444885360039824491323234189312;
R4[2]<=640'd8062250350303268159946115414623899031592965841607467990114811232193001541694499364607194866158535851322920998431889148877361443354870535123642088291444208380808265728;
R4[3]<=640'd2281220309342235602137352901539902579553527812092717799769772806296550563684698925693018620177469159657051561776075592346727521476188999133063698820823794984047454474876072075859617051351973888;
R4[4]<=640'd2281220308811097609322035004421277134406321858163327707067744630959204598234004615254374293077320225207020527829530562089219587002824449062633238567792311539069609517740475276841850257432117248;
R4[5]<=640'd483067197361028394885979702059607148745528582156210070757080991885686903515645874327414289915278816511327028927022497299829406896944781823369855608454018375750889492185088;
R4[6]<=640'd2823416369033517116424485121890535254668606740118493083372770227916012155455598142186085928155723802319463091402309069673688420344025682445854214516954255419137589248;
R4[7]<=640'd1900515169614565774039411043183154337359382263093164807196588958786671170526389885470797814565777654541613398231409120383169162208686762790892505215300458899098828800;
R4[8]<=640'd966134381648615815004712651352486385720727206937891191148737171616709594613359575380838818676874916669595607805131860017767927286868772868998064257776973201467053988380672;
R4[9]<=640'd966134388087782320151291225480869393332858377412085183757652698127511916400488873069936463108176095917132532636007090546303564370637277071477842000990997591866827253743616;
R4[10]<=640'd23413663082584750992272996485510330025482604840376497101826606159405639336262707663210815783029087939601985382432557297902122651208503522290873078300303286038311144299429888;
R4[11]<=640'd23413663770468892864968617055022439684376704035568609805739988803474300255289499555039442014890350669075742158482751892915443344993259911963042844121262875707234286108147712;
R4[12]<=640'd23662745290811139318683540842756596480892459219665599864766817033877055333882909958485515256322358130886953094552215874846168467951603133483391303174351826379367768154177536;
R4[13]<=640'd148780921589713159942457677477921902147164019287603686397150041182124529806887523021743420186616488185379701550816272927800518837419630075978740208197367463402584033178157056;
R4[14]<=640'd463742638122914342768748082404873646802088428523677435211882082742082694272481555000926988573034813236352223144443496589371249821607129131834759991499022675447200574376837120;
R4[15]<=640'd142576269300693601540941030220215762924429247890174724299836794095128103590809235819436494676917796708419551696677883485432218552095397564420385846975565070716042029721211946674632403928055808;
R4[16]<=640'd17822169899878665565593893169715702788478881105133194859937277034107126381184009868557494990113044747502560955938205126043362205969350794766807911628234153583804813468489256260963055319416832;
R4[17]<=640'd17822034193732034150555496022759222875623235494488232845972366151242190954855604485343587684627872043619725945174844516962048375977776750196275859453810611839199485655724171575409564892250112;
R4[18]<=640'd1064471547995284019493955488386415652983031520529208725512877269310537908884041790641456036311229857775002409075536573519745959064021853065543591941309161322863415994845170707551141888;
R4[19]<=640'd1746594107593114607337154878287229626383957358742849926242539976624845525642902006995211946637026896423588442581984219228322817846936441992744369153340328729697188124125061351890335237657124864;
R4[20]<=640'd1817882293237207503706689911084095368858721615838638487210438942860012403881168074640043507713716245207916922487862913847777021830997963235553086937448166769233266993227779792347692581415546880;
R4[21]<=640'd71323062816362484538517056303695270888065236043558434481448641607563526996754516970231850545980440880387486043250889396084589033653785595631384243688413789132122475709951597045363928871153664;
R4[22]<=640'd2423805485031382919041547721409589099188776849672842469496622910046438581288939111106040730031948155573308108880278954810110678219488885433798601058359383227798790792094423053834754103130725376;
R4[23]<=640'd2708962310052284996927586116842314203329662620074924100528069844794611554324702530631936492203204482483018844265286463975209660330910009196723066919807084752850084580078850759924160310129138688;
R4[24]<=640'd214756087709326351207458438152582574091719725785406217489621219479872287256304900541170353375255853435817192885117094573500542049044269128781477897372229684195762796358736350904230322827689920;
R4[25]<=640'd4433290939931890545645610910562540150964671451554709489910504516304873215089240556575639830530080766446459684746523675140102007947299950941228096259319454535408288311547640116544532337941020544;
R4[26]<=640'd4504657360105433277215334191000236737168596707026897646412942486933306122709911813085358655785261753354268148401843758299544451199261613016561122380178133802595863195604960977825000695711923846;
R4[27]<=640'd3698348483740635159730717488708103436880642095653391042307010286260151092222739295737004520951094071826680798958654071912461293513114503501201421215657755639063557340988044248317846146370239686;
R4[28]<=640'd2407990150457660988591314680815099584063388507309974428413552342996493592066233401682199995053642909584750185941279554854057957569334324764991149898696281374919830534113966925584212329058271200;
R4[29]<=640'd3439158649022616026539470990337287229718676745766157278332082627505901915907681707310581400569187841855380859223374830172322771426669578818905406041634324822394562644522433609421953164275351548;
R4[30]<=640'd4507921554684643619053183795102399141654252233246797875969142011991253570084429656479461352717267550032774982168370307414570409796878219520254170417831952147989811211800069617078127961074302972;
R4[31]<=640'd4560482358582815061701212282689854491547228165186403701325385221221313436566632366254921478283030026818559112044929200679691910558301390504432550408776742416421354663943184389241883054338735932;
R4[32]<=640'd4562005509378412860721116628327600040630332709196124839828026901821223905048091078872618251679742363405026928408527442262510689275914685353624368145409059217246410025027738761847969405504323580;
R4[33]<=640'd4562440617622195218392650519082155635791918763402178406453631627660652781506783482922908691931668606442674450662150292236951643117228577823227715692892139899106675654596858838114088005054496764;
R4[34]<=640'd4562440617622195218393601557613210664319946098599213386615964036982150669681153731039325587710181318431183347321383969850905244206687502781449856588999320017299237308563867216152234868187594751;
R4[35]<=640'd4562440617622195218628611873492526396639499902442827511989086075399181865818151234769714875192782878437344897105084477852171361975600240114631649278433861034865392634001993523301013935250997247;
R4[36]<=640'd4562440617622195186970320484935145597531354314680761384181815816439678552831034409049290543774126597867211390739305837783954889397944095112278164651604063108784081025785792938253821126803193855;
R4[37]<=640'd4562440617622195218503014389252424339113303530096313439787348143206939308514470923899747580785685881131616412070180733684858555328555992062643628206326229996139316746959949182353003454547361791;
R4[38]<=640'd4562440617622195214931215598345876508792396697903989792124020565328687896976903291000114255727603961372074106449244358643168713462751035579674656812494979236036762087619470347024675255766482943;
R4[39]<=640'd4562440617091057127645830636480508007519451074377588085120356068485604490919700803275672359770039663051485902671278952833408139644808336442616032130286695014170493601931503338991743777105772543;
R4[40]<=640'd4562439529839135863350206195717547366102404801562672216788736626236499356228060848759047394891773743747356155338847315737272221277573399709752174713762315768073876769936842268265699754972545023;
R4[41]<=640'd4562440617622194433367150791062136485772405682381488548085077976627244727678263855869497089330893385901369354461559766425931344864893412821192487723096377990508078983311732082525885166828650495;
R4[42]<=640'd4562440617622194712355841293970590787147985193214655452074269815367291964643237162079337410142826935730463862791856228622103845239626598440512825870511133102894267680740861679938785287019134975;
R4[43]<=640'd4562440617618551729201848616301038159462423584751948466713906686051199236188674791089669883201477474545497990798051455522103412160904477872560829957381364130888119979149134519280310901238923263;
R4[44]<=640'd4562440617618301232971261407920713271846618336008617258731242111816280127269699757059868897201353460702961048109670864571487132001133812595995701497300835419623653255399210926330658621526900735;
R4[45]<=640'd4562440617622077893013345980906311030967266496693655899240275950511534964023704057825715545543153381356056045312692084327098951963989683776958325119931945141535606934359802064250448712797519871;
R4[46]<=640'd4562440617609625104095653066850903042400895295345268119533469286897652803817759138670046824393225599547440106609024250817183670423677105637598264338019120656591689612841249555603281285090902015;
R4[47]<=640'd4562440617589493469971461349175564475139229344110559332988103283835057805471180026492033802079548957050478484036580595008810645809073148460506271972492246520049261793328127797844790142711365631;
R4[48]<=640'd4562440566583154481207151861510939429558727461573417298745284814600535006772011978736154980560883970713338018997933187483878658247711031873311929919330341507361184742431025178213467435395121151;
R4[49]<=640'd4562440563315410464178292353812559167385636350297736326159339463219482013565230838930100207452487837574433083271371035597915330079805615281287690873033317838371396555861383949855887347272384511;
R4[50]<=640'd4562440613519880452673567703390085700741282629686479904915392280066816342610994690444959827894913919707597861351996278468778148740581641128125003558790454661833408093558520630174874797437616127;
R4[51]<=640'd4562440341567891688800048936491663868064057167309024694244598475304079945675050583095779497191323735481551977375540693677721216941603261340772656755575397741642973408748468272859888215733043199;
R4[52]<=640'd4560769529363903430939278682780288176285867259446600114313968514441453423835211712634253810981944914199858182187210994729708054095732731311949666424015906544973491275536446818946829011675774975;
R4[53]<=640'd4560769801899936988974083693073190832173960788518031024416021148469960552848444247336561344501437635619865596063478548084362572740708661685147279785714833497156381530647369577929557823505563647;
R4[54]<=640'd4562440602617547430079749987028326626601009635993893290521535300353754111452480557685911424484183992968830856999254869621765111383697098076669259489613680778117130325904150460750205189852495871;
R4[55]<=640'd4553459968394650706207208490932823072461030010489535286226501803345536747889944484156038210098446727499805563578919736222416306128759756359967742627491534339999543205114737373910129463201366015;
R4[56]<=640'd4562204975077302935522852460681935762634380293168374420103725893597233462925277149477299375522740658041690600136983892730375558683367868823197965911042720779436405630784784871337630164378976255;
R4[57]<=640'd4562431912204100702858748989546711114660628584212892541595273534436793044888189702750768134579131719985333796607808631851853477904312503036494221775459802972252284267936009793598492457199206399;
R4[58]<=640'd4542947767175072780704279312881343865618704197335904307955934731246089105446918655730416324069029227161659076836542619130041689569252346101344676155924763890600937639968936888114313858572615679;
R4[59]<=640'd4559057378036902236971489269908478888683722634897887254581875857571500986050631277477818239966491713862554851919412460216183878534906435300860213393142474522176854246584449261270040309879799807;
R4[60]<=640'd4546595877934823789517621113394743894803084692431739540583665107910837133576417248046281629608311002259295489986104666178459707919384696440812372514040070872859919423848423135574184271357673471;
R4[61]<=640'd4548830431692649716193919935185216804690948386182872257402794570195606820020775100856526734998818451206723163696643708316645085457286351967233532904765067691869295623735082306615304114543788031;
R4[62]<=640'd4495119565321116430378925854309397873983116691070910011679098073730752034360021928745084943982142676849679209637132200411889552925764210146514492751154667964832963113288079520698168297190850559;
R4[63]<=640'd2227665536472437270019235171374739584435218824541378771878793767300954956210847524664728046496452072948347656163080684692850773347412822616486497305240447985730628703530424425571615844405870591;
R4[64]<=640'd4562197780850535593658705002288757595165720379937330609860811312708789526447495067837039645644739729434142605837688768149979231934410437786944172565722699302236071282134391063687700034614460415;
R4[65]<=640'd4562301658694618725577116918450357716971119714780459081918619875638910439974690812457838692466199359938000104645453640186398866933938231348247714509150541249589393266639938955661473551085420543;
R4[66]<=640'd3706913588456028383917948708777851062845464484378117322590117508419967495176926637369416931773811954583156091900263546769375503084641377136805372265226222477517732924810072432748473475799122943;
R4[67]<=640'd4561535830425087772163062162447967530408436970225675617517493750696262202591198036377364458675361069894646697106781331075926825133091919890018105070213550307469090947484693913603822327889331199;
R4[68]<=640'd1121082734377418144213386744977080343921492790658196800269875358395296797929478301370464762706323463801723981690182675264960067433770760818766415024627749588403162113441965629492147169602506623;
R4[69]<=640'd549106807525953847477069064648470822113813735579081219191993110505468251635862311087901350797029063369537117631369919136486845978787749903338131145929399326017294215585474745932216623223127935;
R4[70]<=640'd2558472100721396369328310493877418560897739439722149013958818285647237297973778873052695596694577961957040816622798455714066572843887773433186683923086913422684261195440596841635388975387746303;
R4[71]<=640'd3556331946777869381013890221655254307693129669664271099187062561440438293003329819343480060928776924119692003310345885530217964113056083722904186475292761625124983186945879892316384787507840975;
R4[72]<=640'd2568045668645413250077913447973845702328655955593097745809117376845909042580623686281628580864986885547496678698365177203567611675607291737392731375368259541441769189298212774014973349493671999;
R4[73]<=640'd2737353921914897343368718301218331194956644714369886771990057150106834219981581796777971459852946755225688607066621636238103796375988720608905599384970278094478748601915410932430835633858215999;
R4[74]<=640'd206651258944968845852470266304025224196774605035426199097468750017177525481835765113962144696601095580549541980691594032581132420544070763390775344334895851252318238901463387348538664024212287;
R4[75]<=640'd284135334985824345030047730894891316787905978039391987227447357483349433394418801172116698784860601549718546768283416846260695546903662003411050813908822664964889540634498287460309520394453823;
R4[76]<=640'd140846274249668473451519305279912659503349251103240643925137329223586373431893372831765164723762739482926493618752102327400297365027356184462744618041415383946119865914724305410779603499221823;
R4[77]<=640'd693259154461005055029079842430738439527635552290909340659278104867221707172525789207180406862548558471798444666239626880887773140892590460124068255688379566203831432608188405545590997279834367;
R4[78]<=640'd6683364601966611962266314201584383517141653437050804297484104099163545601802767986816082652268000133218137077282568136150357311372358506731399459873919488514828399129151160119866122038018303;
R4[79]<=640'd2506325462296382043408981899228730789571572747560125721168818264341790379406428486988618020666514894622532488120175712309528932963338882748631446580641387270651478313037384411953729318027519;
R4[80]<=640'd17826121300786589767390884173316545823223366659989637845472149577839697506185105663626239071246840228537466278075323929545026634867626764058582514019703243808836162366225646898678402713125887;
R4[81]<=640'd3421830463216855105382642650696106695091619504931766594848966827214278678942905996405859459488385162225028531050644735801039975302614273142505985287292630927113532009561709689833595221395375103;
R4[82]<=640'd135971524721621584604006481244152992331741207335640226136353094130807764186576154288422290321113675342871593316836931018464994663562893640893483309894436580967837829752668196725258727679;
R4[83]<=640'd26733186465408824258764345533629757433286526395395657776004089284100182312949979407443059344758727943112636964343624033432653826386379714891982441413690039116401217881511303800568810871727039;
R4[84]<=640'd4360226973103665792675707076088647368200612396776681958830792373624743005557319794662798496431792335140876757232385918444730917155608063461084202286446545850051790636441981132211135;
R4[85]<=640'd4360233094531102259213835250548561587302679880027204625971600847574346054107638496084220904818502545868840811145716942503269664612080126254249024844372321538025020305796740526638015;
R4[86]<=640'd1782994662324560501463495356723095082967141512886877885337744466530565725604087451434819661277217083756602017776723568723359771696569265097598429792445876863805451218201235821695039;
R4[87]<=640'd8911016857908601993181296933143463821106753681877366206099651332749229331156345396518724605357625436643463750078577084284197396523255729177683374764943027784653865282099736793538523329214526;
R4[88]<=640'd588144515466901978677054600682063423120829121570602208859288628850633318621244542520626043961815672115853093362230726956988657370191456916505433992296427335536372392524378791060462476294385727;
R4[89]<=640'd2074753827455989898170685718531095773473881769282593766915055458864182823714916569673835515086612602149482906774428857712393462381461998003170940455699673366896503038662651697692735;
R4[90]<=640'd51868940654118465747568131713490002233543818322297438619825745098329248706248768613704630004145227004158782222796306342134301852107769626583084845308447947102733044032699165174662175;
R4[91]<=640'd64317489339932996420447282830471272576059992098443540151667898086546014799705582832938816992242903930199530473206647817416953584350184031905977583820337407621587748735977636361143839;
R4[92]<=640'd861024415249497193419771868708076102684622887902779136166742287122550996104472758159742625503801451053751734160207582463730910552958000657294200369418517325228677533547707430497945118;
R4[93]<=640'd323662212397934943571674441389456632473814855522680737474488821674437946742203112811354590613546100788629829939630846270297397622963747544107536503281076464936201233493878300949349918;
R4[94]<=640'd506240891492531238758961871940014758078583197358919264215475651832742680589346171132868216899298686294706968652796858641286238984167922708322110847460895366584929065717391535208661054;
R4[95]<=640'd1140679772128083665120419655267807192635109730723364643333717671812026148119988368164838431968374053506987640657606692122573594375748018604143233300541198587195889356833565846253265797863440798;
R4[96]<=640'd30074681928025666738163782881964365096186144915654454138431733777436226999692974274051377303707981953224919032646339901744221659599123117025885556445462881070842333379825345554171930762811399;
R4[97]<=640'd39418363890060247330414018533782553522827132973726922153900023168158027955975215610044608150554331795406181235435452207892625626957497498918798520054886555148360786953355632066955520;
R4[98]<=640'd4678575748919113098124266298430475242578750335499540210863517928950404407640394731646648467639537848989483196750698807950821330192868345018242958614666800628420127312984042056013841208;
R4[99]<=640'd7336340470818305388639154169252882630488585527572966200610568345679301799975855748302221231486357762577137635683179339575940190269616375622061655622788334002788392837344031432756986128;
R4[100]<=640'd6805204963238274991099619787828682356867891499248484149067891857951867981861943521532195533991564239315162167856034946613078251725330019601219276421008869154436225094014088847166537729;
R4[101]<=640'd414951303869091055681635916673736993013558375741558807129062198885243452347031722940075571024854822253854141507832081903152246410909366943992076224207517120626773514979364455271367683;
R4[102]<=640'd285152540709337058142642825451937598189164086755300164473302592061316604759273613776439272806727087218515275376012138581819488920169180811067815369302474001433120211410892746666903573117273600;
R4[103]<=640'd2281220336429738337533038631605701742447847874138944395820271383328292791445148736824870319482496684673876818989107768752402462288166698780784332229764424577482396271060011642169953179060404224;
R4[104]<=640'd518390672884765720370429182688289601125698730824708467186664778645571447008759354576238217823474726572772279587162380789143847125422485417966440695012946529128715972544651199011675439119;
R4[105]<=640'd16996407667468892076737798077064998408792039997141744525027878831315631806379448107439347229637842590895630391499007247610477556697144503326642883940976316306866235160139066947984687119;
R4[106]<=640'd3900966358310379224426532317986168627423610495120946398167618157490995042675642358970015189933998245612684974759816661540010380107713085247982846690863888905800413092599562077920617555820593;
R4[107]<=640'd73424516114834784500169248697523093997126646133100439642501736165286096234233255799917873451014803780682237396343196376401805779009519962802881458664028155734460159526395228778390548906033;
R4[108]<=640'd70501132598665546866717391216338703884343992185183654194155711076987088608195439020203791115733532680068469088009751657052952710406753162065161159203860718477371773751303795315536077783089;
R4[109]<=640'd35216573459608839674534114907303496323423218058261872728233831035058173548408141286022586588146854117950815767236875674399244648781061027256838729311550133697751119288642890297478999965744;
R4[110]<=640'd2283222350086347465576348517083810190142440938597245173839821499426116665533402774618703862363752114650645100714439674919536993272962567138768355061486521714665524562083673368843426827423711232;
R4[111]<=640'd4005958895097051652889123981670409059735262633452394874103145043204713033226787715408192809886756046823928549055892862429089047189354773307332496820542270134667293740404454417023058791735754752;
R4[112]<=640'd252886944045321076990920211033389240767254327414296759713665562441188438476144574251731385857828905184346356814530353988162657710697789295855876279609099964490867961221215329236090354906693635;
R4[113]<=640'd2290131324563500955661334173031293262549292092155928269507273586426239477728712208708283841499840334506647168574248542864329876287952090773425503488736468648755697534038339216846480244054425603;
R4[114]<=640'd277146494848884752061164064611526153521006060831449095277272227654053015095973568924827926299099969788285899645460731660522416595840032271169965905852479472412796850921272212723719659923177473;
R4[115]<=640'd516717093855235470818162752902111233406769672292078167050580546066192776524987393019062971781312927358174756367931269379810956734662250342937765314905704988161967646844844092428173969138384896;
R4[116]<=640'd4295110096284503110935390066897507899200703194079779156963747212612515935050760017558617833961976802993081442608015504332850473597268309616217361596519653984808989083184630191140433924590665740;
R4[117]<=640'd3493118444961487938184475809322298609966955157933972975191676846049724843049105352986667216469898670852232653166743960366655877787569575183288270693259006701082919907466255519991779717950734340;
R4[118]<=640'd124753963757683128943634079531524507591797517221693849121233098139315027095598031437389191288611953012606857084781825236576511081684423388830771526489773881841153325280874776632994606457290752;
R4[119]<=640'd2156464985962550319358139342489430033616847453118599993737511487366611860548037753578893483859682889242834861096027179800811819632674809682921515449874376222650233111776796789845855171279585313;
R4[120]<=640'd4562440108271229844022415509768124148720639209292024817079835134656920440269933302899622038156610645102948390012581089334252231368975797201542303149351089644502334809290093077758756961554268928;
R4[121]<=640'd4402041770775671255591938716172729923368245171020330157468597106888541798763835340927870855109249814387878998176363362074969121355032716522225870215852511595656536646967554223477421395553550336;
R4[122]<=640'd4348575128027091454236731944217651220690488765659547053928985785202905376567490340163587841463067089237458627526270598145551795268732357612648373225779899764065026189448678302936404160407666688;
R4[123]<=640'd2281211613553076249414868274059661627238456908053478340560578633224999081184834501240649746116111309828972983953685468040347153452980877457760919891445349295870438389187662007315311974986809344;
R4[124]<=640'd4259188398815107768315125390797001653213792734625808996567614567316019241758058277856465137246388594308249702601270020831280726596028594642812309067180337351568142122068951014660006499083878404;
R4[125]<=640'd4544076880569960303104999796174425947757461633731801363486622162346185398154759476218921942218982037340125115318385427654764059660513844071464685901699665009946152087106592751439129772649611264;
R4[126]<=640'd2280136902031570258953856642096326097434169291808060231104533647628737894516268339368994838012468565088593279627998320087034251915638028198254168612580707847035051872546089654501838545621090304;
R4[127]<=640'd4295111073843985209985529391414497003571022672408622365654077288721006298467614213652455056749226808101024763552965141941335032057416696748862761318352960949667990835526715285007426302698733569;
R4[128]<=640'd434830212827563267980696959212839146689436609045038243554713530309653116377222887775242873429484469823634043337652284707939877153953212322926173537265691120701337563301308791480271889552637952;
R4[129]<=640'd4009957607087272966337570531349291403726349179335505133760808167176936517922658260844062370335063694130906396786370219126981045416203656860112065493868025755921703145738941835997072570709966848;
R4[130]<=640'd26174148327169810011372317615121755369650513566084322184230135892363456038050167096110088243701427396001792859160825850339592420450717449895218071341954893644005866042707571857148766846976;
R4[131]<=640'd127408802239998289050910528239029691639749818430333985281926026611566026827382087733103037167921239870891961160194602450756656556949612896694733512268868674346244042613812111546703151232;
R4[132]<=640'd17822143867496378550540823568202814375619135416189752172488950953227321855730579870427194500192769520056055283522269752609019932446431444029695081942879674743447158557564857610372284724019200;
R4[133]<=640'd2027256361228197215350485123392549366336703330762777900749234718656289611570538606400936458429008422245205157591648493522574039351311945452287140336893029474031910544405213265423077794815672320;
R4[134]<=640'd2270082554345210690214613125671383423825728882923453608292753501847192328771309620616717173424659177524827238068874146592197914792937911436755610565561743630678968111458108923077085802125852672;
R4[135]<=640'd2343580294240471442885302035941021219813480509933258748697865781620580260438689514736412421610625323180387901325914085965648729077547675137946388075098040441679899301432878200129837696613613568;
R4[136]<=640'd2415425588397745255193715915581533551859597543657626391145792642725801297595861957006035499522069329640382067197437553870168235391191630206489892966628925947826085412013910507370184134581157888;
R4[137]<=640'd3404004608810707498242983472221959044347512157978033167171102268537319209306412085090813652177568199433201609530063121704401028182181214478154476958959334318072597078665371410519432061102456832;
R4[138]<=640'd552474326636128691458325411978663590431406907125985767590847258409032232602515407568647821220674693531677171545858113914950581594787655543554701607282297562312341694733126163460715887680520192;
R4[139]<=640'd2851455426907481874894102604377250165013708679344059252228243180215572597358454349342793490083869210444361972854865985155088685074625773772150501141787381032968691724078259824498190458212548608;
R4[140]<=640'd2708949031761078132147287276322976986171037945394752844010041500317995135900135478774866692588056863832818247535268747905841589485609594346953335534566624296617049170364874093885595906381643776;
R4[141]<=640'd3279218161527997740143229729220175096601151850089741574274470324358849430390707197775955883639757004310175942472752539557269462150249639851687800433439532417175107575216285619203138687978110976;
R4[142]<=640'd3270301433895826842950831166519747496731063121077235840145438300355123781558471622355197310728076637868572982815321787408344708422325617976452205680222171092719443042309652816315986640633823232;
R4[143]<=640'd2325072166269200094326831047704535769425296496111635357849585216866196880374807091981506021787596174857211061385221916189918477461296672932409178264046230902542454742242928071348237060978753536;
R4[144]<=640'd18863777984168301649228900491078136175218744293280303597885612199353973915561174278384536510729621586050732823705684397644780712571488976190012300144367114852946556882345442574253753876079364;
R4[145]<=640'd1113838867915249745766474342576162894247380690097107332599155386513570427545133111851964237458017339969967078343392198018360752235593248039127226230552430621406957829819632917372711737194496;
R4[146]<=640'd552583759821360967278282723509920410498480648902950986967597525039779570885808859171563013603994425884119209617457728635049725016051181221417405379358229608551495541356510115575978159732736;
R4[147]<=640'd606088378742461019275871641374882118627696600960324318433237498411330982283067000296100854264517235871189803434118273455012656873581060462857257389075316527215674746829088297637110353129103840;
R4[148]<=640'd65266103570336238683107954527524032157735108264126849568788475963021915870859541558213047007975919564390069788515599967488025256246874577987160580080506423722836449065791154877950152605664;
R4[149]<=640'd861514322524512824134125212839273726933240918795506911438588458633922186901510854153685195863866630246700750157811719302727122830495680880223431947818867845442196950745911857176248361942752;
R4[150]<=640'd686165700335641413194983111352438001305084264709576597882711738769074701582480458024653903600390859057030531359716551829594417729537645937978933461618898376170583485016736513928776181662875200;
R4[151]<=640'd829014456175685583368940544296028000605577962684732976603235996041417344553175409709173892244509469585349509551498473909396791259605390824940079164212180654090880988382455231258578541573307904;
R4[152]<=640'd1076424067688759021388719885167223660828019888148701693944749391214403789408088578311594184271101962221226581935832024334353134746610525538528754510051469605896358479556699789113364669481877500;
R4[153]<=640'd4551581193298189361484862868126352832690865656191935043785692075495478214933466537655585149148995743016317454550343330811855858239259680012891310127276009150544632395674013403775458137730973692;
R4[154]<=640'd3979082320726102173562742776603993985445713718170897431371794270564815204692730906040033473904153208536570663826682393291531420455614126359103034364078896549680806127513797879900506800317005823;
R4[155]<=640'd562003213519589124313648304141702102521492984946686465578413852338853930926886191607542831153350343821152446297114721635248555314016283124004178311203408333765129235982344167104773244038938495;
R4[156]<=640'd514089228086064989752382351259242253758648620164941238770011492650924450299829329638692470698347537768058566434147482542602697310440800782458132773575657963724351977314053802223846436430151679;
R4[157]<=640'd568022934464493086779911545139538873079388016503359928590870713776064927495539788161358882741800954668190236489618677877978555189490471804268118716993509929819670493867808527758442937048891391;
R4[158]<=640'd4562439666889338068059189648665512309981678125507501023537586743929651973062935054519197346723591047608347150686744403377215886316704728193772031791772613227537248684429759493736750559231475711;
R4[159]<=640'd3416327492253986848772743333598510285762198405568188589483561331315030530373514533019328942630532908418721394424741143558612519969977362713333958771441570369475121020997963403959754133461925887;
R4[160]<=640'd551980347457824653564698171853604998850561727488147206820246599081546399200633106651808039502742041407790641529376875592525325970346753711139524841719032882695148608071834173673357095517028095;
R4[161]<=640'd3563870702490490064366802060171694272451971583228597364004136788147103027105486283429807695644057721289795232394179789438384408483640898068930317507344572049122566201808703875168947660938936319;
R4[162]<=640'd3563879302477691929771468955207258584857461434155411269139399744068507825099230424410475072538085019780531907923553214232740478248169206708750260991391047543320843268035104791423372384167657471;
R4[163]<=640'd4557949399975612632441740009245363679770333890539809624448465184317560539905175506786603033414115005483631059995512393314417712945408743120495856026751760065337568594221011555156367678516559871;
R4[164]<=640'd2255600507024715750228264959868728307117291684071214249875719351360670107730247794913473954214614732634851236005977418680373034364617478612165298690711289303945939470766504921337900057757810687;
R4[165]<=640'd4415547412628048884421336804634802902169498228212813717565950308407694835980156904857818197845097260524283307341276127354440821598213849674314174221372170132249933236723470751780734307741532159;
R4[166]<=640'd4134423978471429194502837993689272320126884718463880745753368554391999188270123294101338979644884039748557429170887754381170695864527085206195011928727130042481963435369578430818093135099396095;
R4[167]<=640'd2138643255670292634030099001693317500631502348167347872598815136745446448314472292199344882141313878254922569269982801800608727818818491413380427286552946161456965418881949396349144940224315391;
R4[168]<=640'd3404008363458086632258682123033200423709751683500681307333405551059195782542386643163725489854127083552629363663879794361945909665357313716674816055701844364369061021273863297320377940453883900;
R4[169]<=640'd2637660921380285289357760956443147101718618343942110532416414890836283782539815945259025307115846882891123001640624257821841056217612118786443510642037269858953455274431032124668374744664637439;
R4[170]<=640'd4134711757137336554042817655442532584524135880296421184057775161255817496567882531977140860883385069519836123717209645994024060979713776884715417756736706514374830489784714889946049435979087871;
R4[171]<=640'd2126391372777446560132760759334622726171608906651957030439848756722917652593800599530282667830508782387081976369149286137359403084661051361245601377011412082989225758957440013808077792551698431;
R4[172]<=640'd1680840384087654391785258714289573745868737947199956086158037959222471182326852776284454152286352532685435674489888816784099152117586377633934724226365235039421122296195853220669217562058358780;
R4[173]<=640'd4330750750981686460987748255793731395961783748474903235890889383954381773795205209118973242980676794417986054884462413507036492668973530429525552658909596740016503289474495732503901528981110783;
R4[174]<=640'd3207824412198853617440009847138729538583285591754500906716106493388748478201406731932749307379401280134736136740083684621476770921987000571381726683992896731557039306279722233927557374095228927;
R4[175]<=640'd2842196457593656594459973325531622978634389574284981355488547047761679579647741377617291275219858472212646867509836396772351144142260609384660464859519547712738107470760891483661309328881647615;
R4[176]<=640'd4517600392295704267881684863386110829877610365948160917111168980682001248751348859239261620975014494290291073215666035705148831521460828065763336490865125789978391318667325578026842972307589113;
R4[177]<=640'd3412500780480892442454335683331904189595578163306020589636205597328251115534879804041289971698890466952729973683739660186782390903169973887482002194291451470921507677074779400487465332918110207;
R4[178]<=640'd1131157673080395908010408970915739802429456565181176247146409605792081528565243868913626064853430158803648174619972456888859307892684028824732273299562729015894370588498008218063037466627080191;
R4[179]<=640'd3288165421223122337654522671243520151283318974051525926718108189944698523435156622067337087746270123941954565701294926109436382384355400566123117957965718807319725824206011807600976123721187254;
R4[180]<=640'd3733716204354118902387834242605902532830597956178867350103921197046045859045093110210985927591884260910951673268598886686527094569013672285822415217953230397816486236637496155557862530626306039;
R4[181]<=640'd2343612808270042060978614239965326720586069693610259876492525180292735106805034200476350372838599932660207327386567732698098345022614198295456151495532359545484230737246865204844747164276196351;
R4[182]<=640'd3867381332284303106343515437529044604684779693901409173641493186897428550525166525446963403094915591260247369504214823401925711079225223882803841469555723177885955629000758135704969211759608824;
R4[183]<=640'd4423763794799402582232545092029093879379397012808551575919216895197212464397005580531378192323485700741580135860166708093877926514486651792096417804483119027509891298286226561976926945258520319;
R4[184]<=640'd4099137500228981204937229591631059333091969433828762778726040074526843980553240142480192010816942422515442362327763996894194473981521845866384828566618401269546636165198182989849055123904437247;
R4[185]<=640'd29747877049989995710756061796224437448861775698676143875203623893820149925920015280192278677305086993104639577733872086219442988820910512851241836234964198190680618576075910551634624511;
R4[186]<=640'd17822046414048043242746037658032061201136799998700145595780079791023070305367148579128516116719866821493703240775108308326675724466821852110968219859584926893925007671365041130464120662343679;
R4[187]<=640'd17822170700338362366247123650633337195980886882714841350456057110317784115907078710389848101864865305573400101487990067245932841476278574016328496852144630981778512577183219615952861835771903;
R4[188]<=640'd518689444751497646856109089182347848349044334525853119598492785304310693509058285692956840694398562631366361431419920036479417501129848665227609723458454794095709567585591092289535;
R4[189]<=640'd518689444857168594772942296100897044524041401293953986106950744642412432103253382680194525497235509038801190038636562377610525101290401286838631347028392545519794761508423908196351;
R4[190]<=640'd249508471285031307862216859433885745565785425414537731295509468088923915405060465313120992197110041771128051075120425221734258151581651075828409160000735360760091208527753399787052802519072767;
R4[191]<=640'd4009992383168965619631857806932766494214695657701029901052017981223659954556852251389352107234207013335174991067671416324320506151962040244355057356635817040792314099201618435226624376757551103;
R4[192]<=640'd4277707414719384991725235784175305747392467100209793722141719563604516782716238432605832513558393130234937208164333961938760388388942726028900169927599172391499363712725333283480033094689286137;
R4[193]<=640'd4286096573602886075600647342144285556650692239736457519430750481939808052501668045674602045759601667321904447126174323775374253374459311120094909417784315701301086882218216769453287328354074617;
R4[194]<=640'd3176205333014556175297618864364343052762645964765391181586696703626195678926572263747948673097844897645217613388527833685370556473993730915166490298802636017367820918718216525020127665814765561;
R4[195]<=640'd3139177621475275062725638213727406685147017229906769564364182050441514660456623415847022260027480120459832081327071895346457240330592696242433079751248218721024513773932698859741805566036017145;
R4[196]<=640'd2869347419676329041371581296281444097541365661978903189584407411961370153532096845826453311247780727327513911784006898555022918961598795473481813743491572630692014071658968353340924680211005433;
R4[197]<=640'd3187916271394960944880004859640356216884270599513703428088692408271775229455548538583200058362161966903211405276544371430955823754747239817157339068484729584752627686092446126930885179340750841;
R4[198]<=640'd4415382724929614639607804385216933438526258296480859554312603992524791895624549046304031856103513769724192987536849385171220436399462454853340034392678179234457187677610013905354823358872551420;
R4[199]<=640'd4526666013591199665673312472392176114781574583737777077404799639411930004660392383795440542552567159474785468068273293435767841847477686692679420346351855154026975006990887988127642716377186044;
R4[200]<=640'd4495399649324021627960642412496555401548779642926032237530539279112988054610957706236238896063141136581172586921667787576364795522496541046159252740614213102349492108085659323434554115431596030;
R4[201]<=640'd4419864450301033613805240627371237048192515827235353044243672462939566933698638483812438115213711905847737613724499858180426257100282714005498739203638175067800932690862399087914026755079208951;
R4[202]<=640'd3425884584277700512383659249031108014112510742811556602629308844346906811708374710698618485300907834302547599854604266023908557547666662891111732240436451189290647512114626964779458455271309299;
R4[203]<=640'd8075065250843568128988507046376382421707047661896702241273150844976533457249135759393832899760363719286041775119644167257338609775545026328454772706880270797776401877749741798994502020431870;
R4[204]<=640'd16150130700859704239555133811717031235305803985404256971827530222592531135894275252341869240905093510159224983174489921283459838594601331347444300267465838243401274948548721571969251548332031;
R4[205]<=640'd17821475372238914768838936682956001223152703269516748338040372584175036227723050805672339816857262231201031869015921965556748117315969366842095429544083253936940970528878862934476630916071295;
R4[206]<=640'd71148900012100015705983072875368432730829338223385249666350628947996125850258313320544172379767261453112041103697964483900493411170917087858532611281397346650461054934604248678475027577831287;
R4[207]<=640'd2280976614201664832339605116983622509070381507811628454762122775259003567978394740273103026083708337127913493008793680945728801585839123015766193878418352429249687574377124783538498730487029759;
R4[208]<=640'd4561988088981794662787168654337006729064414486053425312988213042173850970825233344763318309429504196565959948242390387771432306186071086171463944926708578010163748725402286220644556126558371071;
R4[209]<=640'd4562440349722208438971107878266301109779162200763756136889126244072890707499609375607336608523839217712966762651103244664243429235749805628812197725407757830553283563017989927557231790205699071;
R4[210]<=640'd4562433004290724872427884701971743230847712115281063237400777031028122137015456018696923563259404298508015480823664080114795597408058491698473573544777534709881267654421504122602857140844495871;
R4[211]<=640'd4562432187400118985567532072157679143350292526971055227905093898392166834803248047771703387379829963630338267806975309679023941402004545370755902934012780250295640539628757894688594891628347455;
R4[212]<=640'd4562362573267806724224184241801064121911552509899077051650629673622366793475331169673324522604155617572087786348710371378249618196534698957295181511723024707388200553315704736193694387174119455;
R4[213]<=640'd4562334020318392748053738562098331033946652804698204987136819304654633942728998149165886908512200808979719383672053254272840314442599628949547086014372409344560763700247900853468991031213031431;
R4[214]<=640'd4561882629535341308920617725073549903385458737211144525960067383742034281372686694754211863723033113147942422009713993985480094878014670164785115540633475649332123361014559285037498244762959872;
R4[215]<=640'd4561869606037007143466002459861538175359008919979944066735412182379666347196765535668782939651057584494622996829072772795938066416059361995222144817772939384325752091319241319786508948856635392;
R4[216]<=640'd4544401097723371561443461071228354868720161946356794804439353286760182367328524140175109494880997220455658985787053417115527580741848771056324698895080941584194098488942920662399175290099531984;
R4[217]<=640'd4560767898248454743762388445982421296927658755828601619131244975611444746341007239920242555533635144504516644708627864516897650149170099336440612796569471439494851755242999874457527759154839560;
R4[218]<=640'd3457458212804092425565120830607387628220412428556722002522124223572505768824559974916976303439794175778781658583521970185766618074350815497802338703532435332341195143238893779814527122511201498;
R4[219]<=640'd3430707754913579187403740670596154576630936983395509392924046871862994720073304057002868369989727593097885555591322667436079529105141352949685786843954002403471268668902101881719688331697554504;
R4[220]<=640'd418790622349043461681845152806946245037893784377900273039871533988680498589360569241378760106956807644639200296317350976334674268813202466984034982480205382429669664492330922369952523995228;
R4[221]<=640'd244738826622544780399924393826367682058344710503978953902962128289714486894348892985049330270403609772707648323265306656401543860207386628562813044901272009947411631547596597230801857805560;
R4[222]<=640'd5008086324681602452329381888409652482526098474501135949850156520905790180793757341835728418304481009050671951111095336901122278223567196217905412218105470084861276466106216341186796932168866;
R4[223]<=640'd8629267250183996486446769849701327088043483257900796679973985522864323969431358089991059634262781259598196765529137329214874309729552537522409382003692035053890857584499587296560183627954552;
R4[224]<=640'd579212830722434599728573998957900840742863354756353429930017744863256852893483144953557965359037922891984400304284878163878769793001596904578756689383463069093146594524537516095453849612632053;
R4[225]<=640'd71279432491891335838588957297658002808581303574118511040987148307457184444168878403648965874269222850851067991301668261361064417821562672486493495137790091847359360181538257128971112848501246;
R4[226]<=640'd4490874013711885038042750226538211113527908675662298844264262220001937740374878611999260514429675813303680181384861011277798965633708417011731956879834043358674841225040238502621509657372503934;
R4[227]<=640'd4453280662517693310513963593126623756312524626920295580348137084754145007940622957789417776093227151122837319039104134374317156612537729390403133616547852932597699321559266621817338298471865883;
R4[228]<=640'd4522341045134579140434961259775512783596642213898498502835027937477055702900942341903966671654168275959614124573558119788523763656665431604607187692206642802675884502106120283698207085542982458;
R4[229]<=640'd4130256307810891945330345063719150938546548550866965218189638469019240911257730582590451829291044959559416873341442127286780818809345549995037780124587442463704918858237511979029042021984003423;
R4[230]<=640'd3453019029562096934762445584027151509435932760703208084885500870221832492730670483240471476059373616708148130597918448118642098034275747946434255749063499528361611677486553202420305924589356778;
R4[231]<=640'd279378580176915299766934507985168973374295022634613481165335071142764614130247057625386439955026702134719721470213676498794747749480956878994259195226045521687411039346934230636506474615;
R4[232]<=640'd8911290898497580077933883122873429466455451014953349169273374401035519717045089477102987779186086933445193445627149332333144373560100021973821408220772857887803035026996584074761680826870101;
R4[233]<=640'd514141576991227575585101528790648222725681721773580164711910748626159156065078228779930533388193375391516311413029756781877509347301892490958210217484693984025627983192976228276243618793;
R4[234]<=640'd106227596731128839505520539342316668787856560741838217108266137606603950372345456427050907760057970258912801070579743488189446599362185165830884417652793023389343322710954908072963333103;
R4[235]<=640'd3421830467465748583650214669231001933144883680137241598286633585959241646458359671810278172635765278856203172774139886074137424845264824633413452123814438697492336593806943681859046461157137198;
R4[236]<=640'd998033889353959146610443877152976734524562853737547595332906655002158931412259686550676509774149839011919369870319672989276548332190698879106023481419146850970242160297400804901859198523529981;
R4[237]<=640'd998312609854058149813250320429447529109318355856619060082792517220116389298440402829851360529092452996018143742105747925122928771606577972016350219258049609203560895371483844959231750174770555;
R4[238]<=640'd998869293198357948334368041793777687441841970399338465863914482148317877358289659720908818263856190158360848002085329724925642194534570056839276995995580912114916504955078462696614856317023915;
R4[239]<=640'd4491709421656588750915912457586407792080236526424849038499858146495306887115443308108768055321964419664426597453004016571837139788329481485524249488278873334088874129822192093204898648794676469;
R4[240]<=640'd3479195134600272710747514385239569180113084444152083939041207387921266166487602326686089794438907994398987356444149084477541276712081259333690856636616764293664640162551936914714447742363580029;
R4[241]<=640'd34530190271055965952422485694310449917024165298315932650934847311998235186887760975291229495626917460291571305822448030274030048049933377240407908949056904226675126888017338268203054000671898;
R4[242]<=640'd33196156209339332225479639869477361769231533533757268771148176838668402679383485417677513350386017823669010845695303508745573877667784478593642216866360772126767225720143521858429974;
R4[243]<=640'd49794192762501550856657711843170054143564079109429491595084504293695381295548891001290974306053766423337926345553138650641505794366669853392329187420826232698997925333270253014049368;
R4[244]<=640'd4157120484065487976725700198533238109456180761124673596811982194344706560450597515253214421432988466971021334359644057991041863638854099272207327494227909212100266571041728488640148;
R4[245]<=640'd4157399225431722127960407924495862335425978691071163860436069038851362082352820711981505536881484875275317163326708912954827421926289676233666310340833211565053116833062407553596930;
R4[246]<=640'd8088940783951846211270276930884699566237152710016244246983593988494638036303889211628379305226810356723491161305538110758635306116887055650126245927375704441218432254034191464245;
R4[247]<=640'd52213122095191879184740268585278699437676954993675976370525146868801038805015103605344874940105836565603816125349210264208449338665181065475833998680984051837338011605975255676208399828467;
R4[248]<=640'd169692746588461259756935373082000170840698459098495579968474229990264181185095513115464499864966723536683627845286110979890245812508852792129320954880650360276734176594062482680355137150562;
R4[249]<=640'd58093470365008606539910958217468517556667998413846679789780127939812137189732527561247602490569281366208041116516939966077343946881847110244749322867891850556264442599656231585061668;
R4[250]<=640'd3421830463481194747071032397041838903558082019767734241615632553675560745283387497675696586501233687020541784610984732802161447290331674884285867497876101272994840921158774051489197488390993564;
R4[251]<=640'd4277288079551621829388080400984402540055111374576927876918326290316338293716483431308000362327310905143542794859814047331527720685053283675149473551978192883941584555331540347256445358961973533;
R4[252]<=640'd4277288079269778951608957943112726866547438875311338188910592689205085903213186195166608355403272156680738256688548961110621768647267972983038001977390775074766445157686100740479336062005562143;
R4[253]<=640'd136220297095225236842045325349253385891386552926362824470064765763398958424431920077490895487260229306709207582498699428206472894369674562056236143543751362670584593370139122534155091325;
R4[254]<=640'd5186894461101241198126560560559078829015609040696047935070727748835297288902411598901381078890306332617758302773271220117298242774000184865199319106462251165016535043399223677774730;
R4[255]<=640'd17822033662846044795872138644224830712168572375668993564115476829333334148229595295789475255182032623151755580738807152384019140368864041551701569023167062193994336030476782692027580382491679;
R4[256]<=640'd2281220308811150257059164973773459932636984341448261828501305894595103593667888803916670426087641577004963583626666431773344533064063124951623889621041758323804342820350558509238375980647047427;
R4[257]<=640'd2209932174161189672093691373195866566354491861896964929516655020488198409605768038239052964933192330219077862210690102398663435021376905102996025502727620387161459160995321273702534766458720687;
R4[258]<=640'd1069530871712671960946632634321777110004024270177845424367859667360905447656905380538617139018497060621661582172142495600105282375790372379006902409004934152284456746446691373741228791154703165;
R4[259]<=640'd142576275676553944529707937070888950378779970226694214293248012568295927525153296502585862392141112477492890461769904998918926237405943545542027329186444163498597066842935262712223743192736387;
R4[260]<=640'd238416770955757079087194068892903882858814107265554592991090808838835139646978848715883370754728514278346839503849942213495283707790552923537871238576275250400400136428178943596135894790;
R4[261]<=640'd835620266727577790627045105073953637864057712359304916000837033022422008909764833223226304849998564755813284611060865157129675175245993383841457433295084626173443218240472053175868808661314;
R4[262]<=640'd974676450584970801967601014043059054861981723111991700147578436690460065671717701146050283269516717993338845866870347324356870771178099799823491954150717050249685838302879074246122580766492;
R4[263]<=640'd3992135675327433677183518391255185212813629099737862145251995580579007450797285830160289832397491644407347940375555261632104577038578352529302824167067946119230886663288642908179538730205678129;
R4[264]<=640'd271942587486065762980523665744732783964301245701493082880582824301185056735153808497054579559461986701261722996131898566076127036930862713499248514924272789463350233462133783553277667709;
R4[265]<=640'd26378437271199907101219097100515836000109548499302245387884827977586346705791052358922753274267555885618252127715256167196100130403130985609825489879663276890616966661251934743207819297100;
R4[266]<=640'd13436142561849587526409459389296580207198126451057929655848236616431095356399135951055722355085422048275607916938009867100048898661990860337562536780990338460615692887513251172504621764108105;
R4[267]<=640'd4455508414633609693770432571577196429800400195379698804087756274469514427148937607500733797093973117247737696116513269157029010594670121346415185826291177496368282251267596327586147480153705;
R4[268]<=640'd3424058216362453110579501680494606323368782618427408111395526814150108054545700700160463230647862321829110746759931801492304359719845881443181385953081228270153628423425252601935633988507361414;
R4[269]<=640'd3422944339258800786548005462429752502888352516693098138139767006768344782628329686949141329818770295038631016961929835068889965518367980640359345107660082878468799022879016036423409115315402762;
R4[270]<=640'd1113872867772999558859756612422662046477099414473897695307685162553570655208349474923304349125707350615098801616483363280492800273552669310328013970963512036680629097379550580605580112250610;
R4[271]<=640'd17396362674738627826888257415745920798710160903407809022996380926984362657970418582633221674976008148656601584419465778469249648720603774000889377993668868519821232288853434792967936709265;
R4[272]<=640'd556887562688769193777407981252651945820403385653955716872805534345300408587747224830980538862826428737496013712869393467085833754600550428524093280201737742607707324691629240568896658299710;
R4[273]<=640'd278469272752380512166541161768859653172330605321782946822623513045476092787411689662475790354473284213842122617140568648952377980758940558970575595897845698963330315991704774394762459063563;
R4[274]<=640'd69617310712226926305068176314876634625473175076314443130613177929560085512065440998620096463821711407780796281724631670126195860131431484921117175017520392586843756406896952196848590896974;
R4[275]<=640'd139234605708566225212820382540354305667870920326284631531962909276932807851250771695484852130902822672928946221543026834923965361587608702396942912988583955549871492553404826210159312095736;
R4[276]<=640'd285709477153286208912204701644059371848489576915913996212076724570572027379957819067267754813720891682482792984143619392409857808007690173720692796141286027842045656056983023858978014235645943;
R4[277]<=640'd1087144053417659032083272927181879117934131635248370747222606332603264124503994941685189598197805080727155617108700797847900524038347875978505239628573176496492014980514350713158937255359463183;
R4[278]<=640'd4562440617621935873919082678021138613987921647649360038133612731223839561950565474792221350362608476260589570083433052812010951133054931835924384367839372433608874401410587393228495810818091884;
R4[279]<=640'd4562440616559927400846815656125247725823545405418178942382239070298564610494633458303322423602929450297444941014245975907438984281037221599597996645572420706294613019882506308808667278674529124;
R4[280]<=640'd4562440617091057225824404507010703118340759879918988154325671621075365950229571408175837665560163386247201624242850507873566977581566679060489446571151990152403777085622507770999175942621721382;
R4[281]<=640'd4562440617091057225824404507010703118340759879918979007461541336673485425703588408203598667906445963120261386616621013453573374831230176443725963559318290503598989074562702609447135972117188113;
R4[282]<=640'd4562440617091057225824404507010703118340759879918966812945195951409151021543028410620670930317368765665570251143328240895799628143512577881550518265451924280913895844063551027254000568794009155;
R4[283]<=640'd4562440617091057225824404507010703118340759879918966812945195951409140506621524840728893851414501437394735941036380690432240754526083775026727390640798956496988885379772079823376848564330888488;
R4[284]<=640'd4561848870147247907970016510123611114105528514668870016215864345160158338660899346082208518921965358087464531591991733394890292347474916465041843572066159165252599284462835576595646074469866086;
R4[285]<=640'd4561552996539446613172648386396365618210017220269575243604733337156184223244604445038571990202761352958386357120683914836647588330053756494044414193296061291274554445793385140651701264393163246;
R4[286]<=640'd4544622934776476679094686656662154808936145271911321624706452584891744690259054918831896234830827907179021394211596886928151641371552933589409037103422213681892397514054665217625582296953978672;
R4[287]<=640'd285156753446929198620384876583481304920618955714194707018587956510993538179434900107608886310861441587571717683263493200054960524771458571492047682983497061132203348865732923736393607081874089;
R4[288]<=640'd2039437107918181467193346316109841411788805173792417344772328679818767643813620461167148172437380483833031656144594949623902499817343604009770302692257744464206942094291927653849913696427;
R4[289]<=640'd2175275649581069652683208499935635263228348613651105756657366319754706820663610916983414840552513159879584161813996682575772803897966650553415689693558422035878077977202440882338544242950;
R4[290]<=640'd531137992816767098689588206552468627329593117773549435161350648312669802442485598330549677085822597722248618625588230755145444631423942549967225106936376190517738670153024367314725465;
R4[291]<=640'd195109330912251078518046330051984774099427920822876301995010855919183686442837736371413630570670194214415456674738689644734384569801774246705013;
R4[292]<=640'd292663972744087502079385999966015600402560541613200366235104078352862794424878852362800563743225183068718154074901196374674770581368128728830502;
R4[293]<=640'd142948280278171516249216548939075277375397900337265334995762009639345050880159818553881160888066146095572251921014069235313261534247322343377;
R4[294]<=640'd714557421054119036835082680877735237476649969300338216161904215786951663239577899220139237910336789945042150822194037122329025408452050445199;
R4[295]<=640'd39536350988354473992366896159518577825438010849746028233019251388880367432136417080614643090458541259858872456970597816800879496179136709499024;
R4[296]<=640'd18196227250887499068726270821291102098207537313368064232597446977371424870064575707496783155334887802645964895371861774437606010981127143536095;
R4[297]<=640'd2953314384832596782348650797056355634027377887386535494194280970584516118951513670179854888225685494173312909395027718680554054143042209542086;
R4[298]<=640'd1429023081902320562151050013231312387548344409620137567732477745561325031496643759613729800956865754938118309521278710437622897613914157415710;
R4[299]<=640'd285804615812621359075059954791049214901222826533381252495993492103708729710220765859556375870130319450240213140874413005343915832761151282632;
R4[300]<=640'd149844025683372897980103025111061862439360096773273112425929167627544560530862196857892793535378321312837503233224378269122142525451431952812787035;
R4[301]<=640'd174817918817695564957369444988209859478822693184966930463866766542528754373614560653039255341550233584197636274664163836544722031585268500071242827;
R4[302]<=640'd174817918817695564957369444946607920161409846415395540118855087022379203031393730042431846181572107289949668307258317072045437020365625042799296294;
R4[303]<=640'd74921965207583813553158334153368090589235276234026481799920123738910910149096055725272990759773257677240624796641422674615399075419129599870760639;
R4[304]<=640'd6392560593909573091811665744766952403604452088570196792067251191632861825564775054451946887628445395976299176438394473855863204396235258334775746861;
R4[305]<=640'd1597945039192998523438456092605969711773027970481682858486978387795275902979669383604688835637224830469054021521326344678282671080168711974633231915;
R4[306]<=640'd798777410312104512204771306835669589470951238842667743935900371325986074985245430980152224792393542883720113102513815205565295725861628381813917940;
R4[307]<=640'd2926639265921242716987968172533163730062380419492979368560972804497613259044587893331207887642177907655560535581692021093527508097935379416132725;
R4[308]<=640'd6345390961119968174523645197810794483232678913471280594377567592797506809005935982746806272140959236836491291833582403405908057759998965519979349207517;
R4[309]<=640'd6354980972666538902658449429656058703640379955409354513765501891703895427556330907839267421542553652653830129645672127421906529385917777383286684602301;
R4[310]<=640'd82377578366055063680981841505599323409270018019221346188858206595772667419316123011571266447939620992791315218739357156731589140231187492151856647282671697579;
R4[311]<=640'd82377578468348483594745450927977584015854675588103161996329835521687256185789803328506841634040512157820247392587779226966469954838423946211108279057905140684;
R4[312]<=640'd53987745104694852810148161769446358284988695407777599883778793095125356377592232959140402594851391195307317650651805690812152558866681587751175398292518494788865987;
R4[313]<=640'd17404329748620063947796289795478575851775777972504030965716135261119977794345337311505470170221848929698648258348454872825136701960440647198781136255830827262810527774494858666356302767764;
R4[314]<=640'd3380343056367347061038978389947770728608055301782835230648937398875557868069957123521827685785507352574063456729245310223605975737106004255199738428033547179522003;
R4[315]<=640'd2281220308812134988212806051089775521800738037348107964774169959515669323741865657657649901020922851873561469059852816483257002014742519961311335349080074158659130594420362844350107546189310798;
R4[316]<=640'd1013065324433836171510912179456672368586522247120003675225639594185675289948354057787138165600231513997380576551786874791388864167975929619374092546669199637196442210404756289879599;
R4[317]<=640'd4562440601156982277502155311838005559928355440941078541181994580582479233955344645252032814223711292535777643658009716406450610834543548029932960123773305752537699877255677968448746910939143541;
R4[318]<=640'd4553529332100448582591135861043645015498747637106109413609074472383231506708951218830386014957090955416652163593568031474353692500633288363933383098466925020663814993582106829377080590269478030;
R4[319]<=640'd3566094935506657882960618945219405356789841286210962540300353838751575451150453664099227166595582603845768785953157989382526077585920513307394954882197413438743036716840389391504618076817612317;
R4[320]<=640'd4562423213292446598816881745273939013601248452646514650216890579475508175033302005320656377923587662604952263269483912382152023476427449889799397921443445356167928093764940350764579351044823621;
R4[321]<=640'd21852239852211945619713485921077371642548809935428174493400248414062465995022739298576288293500674700970704108424781532594565929616389552314366002;
R4[322]<=640'd10576325594451655342829781613007222773908256947816611186596643921634208961129326867108880210339355988167903661890157625569501;
R4[323]<=640'd174518161094061982475082059367653376911666271228188244223464737932782561773118543851222565485257115304509688235053125196961928;
R4[324]<=640'd3992135540419420816311025154987754909281574943842490082159101359472546621503750916403159278666137816972147314202569350495411981970915722445672254173584031741975322027718257271247493424967827377;
R4[325]<=640'd4277288079020808017476098380344023117087401725545525077913336248572749188430979119078768312471039800289863361869285825957200731540311339139642215263524784921753399979804519690071036281398629886;
R4[326]<=640'd2281220308811097609320585802850145662446614253624280012906254765035928420249618448661745928607008968709513681839406336158164841486328469141073904225194877484171344142379997088330390858980366779;
R4[327]<=640'd4562440481650869057548794341165710447461259910873020601179389627185959986359745121562738096180133135430884994088880345745288542350171681459887066890293685953990434071403768825865522959991183124;
R4[328]<=640'd534661009877597011263327915142897775226991270911208870881042817515808727721071970945842809683904376115355096247847267536459792318540698575162441079968449950860293374070233814622261952607153227;
R4[329]<=640'd891101683129270167466909614228116594248317211386612441103438918855521309341705238747988127521866044918256761031407267859018266440739105951680427279842101670970298846278503156686013996738528643;
R4[330]<=640'd1140610154405548804656432137403791625277744106519588255694270562980322227359812049923028380294623901131935168177554745322112505876625736198073420438140626998938693531867544423005111999104905869;
R4[331]<=640'd1363120159161290924351105486864489196092911474341766609708993416385626435789541240676282021404129400721007803169028542921066280912902649791030286254736801470184613152791442058473706929441053015;
R4[332]<=640'd3513116172744022059727340788431384374509873617290798718615902436671422273324952889845734026412896460408742486297777431996271020962176186333668914155324250580793285808243398599448953272635484089;
R4[333]<=640'd6196085860042703607841155349365795333483037151785003790353650870794801119871530191193924933333508693643851707824480615633635563947271807936178688913934742710075433175343610713998178626938075;
R4[334]<=640'd3651410976930690516188427595659692216102680802380314799897828303442821895804992607980769879659862011268501552907349655388824897679343319315114884491895462321197070364583876399784714371833640955;
R4[335]<=640'd872865208864609294002134451256480273753328548310117830947713641181237391360259409222696429008497069420527495517586819394797346308290036582587884844812023046596512215024140358333086542851392118;
R4[336]<=640'd4423232647009580190172818921628138093605639446841564832262346521341468183286983043354964011714506272657604714123077225153611860353760308399710557032507878844383159576423666441606207595645062732;
R4[337]<=640'd4259531464562520572973292702959481008555428483014294811813290200441095625443009099244864970639262774805266821791238095355346909133996706105541379022496109649425976054823707513495015408385129823;
R4[338]<=640'd2265556530484241017853288329926949811765383608266795149714896857714364088556098878718452140557682253315947374051716058974915296955213819045685616799855135827431772388335088201153789960948125117;
R4[339]<=640'd3704477036998434862213789090066210466483639260198362857962310383969884923702220550629112327483721094296378210113633916071650890266476329191174854305648338284644911116633275236810684927069949805;
R4[340]<=640'd2896063617692964678629500623080393282251270705009227519847528243737790060647128511869875953277397817772675244002315766417519940135338564572305444357604700830800442772550941204169658196807250621;
R4[341]<=640'd1372070845625305969072144046578999531876900300418390473047781308842582574792398516781388718662196383092825007308959615070589533011797746847660197772468924580634479996732321027512029868586712468;
R4[342]<=640'd3599772993426750532845750867907330920357724648666468850250589734594958028224338041024757106285082062438156465176085546840289362463690851199615955866032608055872075983107406700441992134421294446;
R4[343]<=640'd784121593802176636244835067313692512710938051864020878701428642284996205792008216556981094438190157542939813684684596341454121542448667116126721599043595410382823797682764632497013104456064673;
R4[344]<=640'd40068582710277441101434270253404931277630310036212712604898485583614291390933958161995552977817204592153124426311521422365150206724329990618273480991410403017033551214804076290444689860222084;
R4[345]<=640'd571386066005670756876867604457900621220472672315219501996928387768283862416468158111856312844612999517857236100051281484965138384248186397959752259523043596279363011457944981628429614713366012;
R4[346]<=640'd2372527246815989733602800188686727565399507441766246370626956828097493232335121304912579426752885995641317006562046311982319717902418307268607232833578914358280487559047701109325083283691166627;
R4[347]<=640'd895490837570956088873839165056644781268744860076421818731338479162341368138826508179232117338714204397414115226641672005139570784512508907474182764978082949989477479254534721943566755594822277;
R4[348]<=640'd1290359182298943053708971056048505672667712820893508417951190880443307857171774454616311224062657275051946322043126900001578571186552635806665121085153125675536474128258735665561390451069566913;
R4[349]<=640'd1407807951861138860600093761313963251845335513182870713844658662890993194672207185178289946889173267559122996859426443356631068990285293482173411296586351867732773726745166426507515757503805231;
R4[350]<=640'd89110166453935313816188998902547243544183793063408726438307758823797549913132514083144507812095650493320334027940672813274044875530877188682371185557059100080198742695590679300015214380703342;
R4[351]<=640'd507927958323392070173490371821391157208556897777049770133247923932223411955963117910519749349473452458070287180761947640951921037593892056331671715621326448638866958894283212220851281056889359;
R4[352]<=640'd93565676664207899415056654994852232330885496234327447267187364320276875680489478687127407357756374556369596709545944213047228633338696049591011457112459867182931420830964803423481460205887236;
R4[353]<=640'd147031777700778606976782890117992835190777884660985062937979318529336761914706273145304596264117005801511744824928844423107108027890664003150456139035455898436755861430321575320041605772246751;
R4[354]<=640'd158697029722115447327527331826551439286530944124884805696090166372748367348235044075339213588800570621847960878936348845498813556332264922969936752377764741699845654618001311572598874685073534;
R4[355]<=640'd152010502731741722824895988965772175705071194611978360278607558570340684191762148629890777761138326808087111502665516440544407375323882733944462423369730105795636944543549559216262827829636418;
R4[356]<=640'd71288270621616355491149216263720617296511042905959957641291494494943859118905399346484461720295277791312232041217226348848678420839249159634194162760037797452268750165364427473753183245362197;
R4[357]<=640'd534661026873899513472600539554597913982083365263144360950652406923902200016320448575577818846749593851046805821084021734562584628654514113749845846875279053157393397539399883208656462853401539;
R4[358]<=640'd285152542850491131070376943931148137849077709034490914542369796586593910431115213777139235934721188254489664779207987843961253161014212928079455240607129497788567165259425984236179352400664792;
R4[359]<=640'd2459440697488487905768851246773866927504454361903214174460088627677841381706052452394806425344051742042323721692390812492262794784162275735209945305398433239075830800190073557962789123058236988;
R4[360]<=640'd1211952799746489895289792137230886519186486205488611428441046591447212762261228123541038841765967692421074374280324064932440908575476069594585109983619539316328184576106377984270927439825711613;
R4[361]<=640'd1316540352595209180513225113684071460555106434152599600985358022578458615928316342839871033888151672823944242622535710372793700080861603655576391047060345343142027865815126472818718244195939624;
R4[362]<=640'd2470030653935093844034228163072019689103309338716152124524636564168657084774077402766226625535704109320252060110114335478412186321609619970251972684385295282177668819861663026735344303592054071;
R4[363]<=640'd4075262031864582460416900890187013045948127192206194478579124046016291338019331117168728123013629574658245738801163018775953009758272548701639151175247205974975038640326019761721398667566051222;
R4[364]<=640'd3974601728259572899871996938820109565082045142002000096954102209945696895838616719225264583188445462362112797721085052256831520910974133446174016581236017621941225343581567713879537737305755463;
R4[365]<=640'd571662662726364136302973327566507061987649180787163973464570798531671252430436614469522847917910136790029760687516102104933729085042475481017400266211395398556407531067296887624796581493376607;
R4[366]<=640'd1427035417571171799141317496168811727732155523663988573978562334742953850459573349632346519071619454935763971371057428949674295696988918470091331076556672581237379754395182779968692671373710240;
R4[367]<=640'd2424118967316997710114869096903409969632439250312631610711531950308488777849249346126587211657091929557291517841884294808307278187200723391946749104530884839344336480396841560700713358495778128;
R4[368]<=640'd21274578225205333566065868132499435539441464692742919797214608528876373192358538692328825006581517177392168977437887795672612895085274049291898990722883470910456771705575069273293753747;
R4[369]<=640'd16199785886712625793802537287528654769623613226539562825648676126251294824003041693145306395039962144534836078003370013540818203434964869357023311494406100113962997992151935869264740201;
R4[370]<=640'd1759399360562903889528145377902852185022036668532391012057144461537210874510675963134009001132625661320927335165834968251157425528303730129160690588797926304519813118665314205276222338;
R4[371]<=640'd497941980170711034917540706805749401326766948014324774977791729340307757395156874326982164238326257297401368221388433964433675554984709202055082942233835568650109325612880548365574279;
R4[372]<=640'd47719436953602983055558889702748766931306039279341302150160739642672728325565371232403244852436228974968808489536367764961949698008040291719230932391623667372413734574463481159288966;
R4[373]<=640'd32807265851554715629686072013761733963906357421012462563628032874812994501863052518003991478025225586415657136113441626197776579332004258572099413974119255840482658365349355098899925;
R4[374]<=640'd1261775149442123280036604250421333677925214647980879692328702628129657296324219124597269547479530872813825691939377328242768371638340728303564101493177258110924978110658656552486249;
R4[375]<=640'd714116078862638090589739520766068715630699217099891752229954714342736617788068174025798961247748793947377681158101647846280212768072103047214534728209657856000574226274264823693626;
R4[376]<=640'd8618351505957782716384536285272658457702877594430729325774411374525052505419923013159513353288109185457519125621941627822360807883365276012383055268886309610352610114115091825212;
R4[377]<=640'd32177214241377978418011276272463218150011583387913317909386604438681102894259669670293660080101536041018709781494467277768323456092969394948105966185486818156457186107965562618770;
R4[378]<=640'd14420568835998464844262472187453866012732927876272002650248685874289540902736991455556549489610473238269713088828242625347253963976660441522889814227517777252321263585523181289559;
R4[379]<=640'd5132356830026461297656214735473030387690490504459229001822754819240286159201743735386097701506127189009611947052399594563974192655926373343422744516216651318524971160918141435939;
R4[380]<=640'd2817645924771374141972927644073694008509342038845846291661483496400698219250335267684009239115958191066246286464596238662778118657199693429061212622114208015714400610795915313186;
R4[381]<=640'd8456906657641975642491392067802515370609462004811644075224472025234688091680046623879308743030365284634049581061692332633415089548623296199064143278441650822420656350350607908898;
R4[382]<=640'd56946376700404010783858762331582253187204693458237558595392242731254392624166925942402590109365550875655712808128173716152026426720148588707485591671177457585941246136962514952;
R4[383]<=640'd389021165509955244048744262977727540746735217734005492121721892739493055638097429065663510828581481454918876833353523610285570689380853955782152080769507098244396603024538880442368;
R4[384]<=640'd2227754207823348159765657568788595921524715490574281271133104402067066107479017034174669821268181896405344006991423264047457383990041477360093784232296538040875161011384451363154764622725120;
R4[385]<=640'd5433554794704402150393650180326387356856495715529536818657225492406173285634325482661969911991699451776245895253750412916352508502922390832428987509537752866520457784818925568;
R4[386]<=640'd69617318994480795513216875863198185266881588722106918489616947435175594376458364211033605538914719158864821982900326741397604288489418405185396725495115232111272184711365530371943850573824;
R4[387]<=640'd1670815655867504067040907998262342429516031725805109890896589653842154240270119192082653091671713884920328965604568116594372871145434857908201446858825854202174937146769122169407881143648256;
R4[388]<=640'd1113877103911668831958808796894426174789277042457504131270686105104329173936513614084436356455346201932904299370750158370477830440928307498688684849541381177679576835557686862783923210944512;
R4[389]<=640'd261064946229297403966963902254457934443963607239680813627906982933461585819225658639303799314246235098659755858479309850344635850653586018628480755855084464504639525445231748949420768493568;
R4[390]<=640'd17404329748619828999772903543537694189706892675444919625065816965633323049014427147086417009493830554521515842113125560602085779945938413834931155639124039535445291870758284757348544151552;
R4[391]<=640'd78319483868789215342240135867061354392432440950778708122645256458234584196797452827198300507782881114632274107953769580764094687144515257174853293902067709484046528102316595067331991830528;
R4[392]<=640'd635258035824623587259204229382227590640776266226443732927342875428556955739749431785595827907754498687317575230361066257822113137350924828017174052882000670214978303839145722352563046580224;
R4[393]<=640'd844109992808061478482801393293371304240239646213255830560954231439094430402647373696102159048819402011578889768714550613473222091527285855746986903676854865378395095223271770643575276044288;
R4[394]<=640'd261064946229297364423503580106875463529129530495097778004306109296586645542148363213505581314188959744092266643518457270579943131463657407698719356077796388920974106773900767354185595224064;
R4[395]<=640'd50712807227139654715598192200693773714861872005183148339708702860075353369265835682816495546836945653145608033992093442693326305450814008938726585545375582559028205584384;
R4[396]<=640'd11318201764286721790598179220961970290982355484528045684747815526260514170440658384243368958790249528934025483244786477522103200239811706242326660681470133008361624436736;
R4[397]<=640'd1903598566255293282705482212608676262773458182126970597455039759678229550131261024819200281336488381952141921803422917386473361821032274759961169621966309991091162698781253745994505388032;
R4[398]<=640'd1903598566255293342339311583757690760974560622774960126553680957827201165877387739131648751597934808763247615777601990846621565665804676118608474234723943660502696994852272869497926320128;
R4[399]<=640'd483168721188783988058984079136795079282191888032909629967583450004268220029193649688022324175661850912480194486718190533709082040980981423722109882802520561228180784939008;
R4[400]<=640'd30315483513987715510339020878484947248264284245253000596293072732686753740088935103881183434183245906135061778818458001013635531956173302356701059869162130482046959616;
R4[401]<=640'd26575533675746121899333260656790674627623847669059908562723836935428141766010339521207091942311716117740307342327811467645864057608610525839995639583802174034373771264;
R4[402]<=640'd454560046287189941071409706211829259797883566139370716976722272383841934460888350036900674087546352566351099590000187127811848860940929095748051242743966167547772928;
R4[403]<=640'd3136867643258638440244703688021872167367296739300533356576688933933981070906557879449644109138420571912141361739902005613271777338340447991315314172478832364039962624;
R4[404]<=640'd2831328860914861958616570136424809044061574700897880791753618094119286297427612415023740530145387719089810347569707192718030796514634766137080575004949553554899842629632;
R4[405]<=640'd139466382454999093651203143013763616276372215875929737750808130015116301368970609964223552373752610960497682383581923585739409940275348922961724801237702824805007360;
R4[406]<=640'd44227007889530738621131778244270482877430404819313664533930087432800985430512100923035908313534436464429680250700184640428482364441251814290214377777631755721181757440;
R4[407]<=640'd1415314233021334543813749418404380450292981863126233708393448521724922004096779684189460159970033166795201602572128400303447081257467864058452707626155355333637370281984;
R4[408]<=640'd809155535931793626914953353958330497147865130811924057774329929938150702449012208803200683919594292684191364688979560613424410220605905108016829788250087445661493421711741296828219392;
R4[409]<=640'd813305051500674619871158529097328344684848758472629968325486217225643988166432863858127639390817304784382254301389668638751968176092506145149254075345469486849144240032252254677368832;
R4[410]<=640'd248970934132859577511017332035638778480134974194525077141425584367551118378497544013141677575858133379148976177146462803921732559936174941466698856601318652683833527430366718570004480;
R4[411]<=640'd232372871857335605676778728194167468950120038865058034870413387280351145416205385872545223864412664770381960952500081840231446019065622424814273875053395894676913040912798459260567552;
R4[412]<=640'd28118204104481053419960921934583127599628174674883437850268513011609410442000921379241825592532195341629565289282257260406765173464973311215232084354188317818880;
R4[413]<=640'd2428420863119553378222277009198503284306908095958139655837029150168205642914170434108036097753693434441263608358450069739592705835315112880555432670290266554368;
R4[414]<=640'd132784498204191774672399301575916976373064406965899269396607903643092626690355702248307859956892546221617085551278470028664491957286810153365728521393454659422538810417064424442429440;
R4[415]<=640'd199176747306287662008596403148286718490060504437444675578409884790493585179353508955496037071812719344009858925169247242919098195215088554318715603667138813599278764275594804376633344;
R4[416]<=640'd63316582777114760869656094196561586869004388796254485305790279032283226954618077198885858440255900085724811481059153997007801273961007116118139700324268260864575251864098963712;
R4[417]<=640'd3462625620623463524900615335018174066576809567344468220643348009037248355586495822334408664890234577456717753321999277560842801246996997183192636001355701422436164019029016832;
R4[418]<=640'd494660802946209074798093368574222221249807624484279467755539491065761455191454089131662538131362303935825199155261676173932337039652825506255138681015524894385335170049769472;
R4[419]<=640'd494660802946209071526588278720914530287610845695056265055260297526879257713753244831999701885980527844229833183697454747643942098662449843845151298824917587840637278779080704;
R4[420]<=640'd63316582777114760720608195860723935941681789197390963678934639244438733253476089751675391958567597061792192988331120452904418099208438685662753886046076629714061789539084533760;
R4[421]<=640'd63316582777114760719842282861963156494997552327578071533105007462343874521330864039584633473228123380181189921753393978065861209623748673333753176100818583636705162097644797952;
R4[422]<=640'd109969158118604284576902255896759354759252202647509376195408635607754686351374076199305177799027913751523671763248928781638627262070957205782442853792701480960;
R4[423]<=640'd881537184268667480877638353478771476306595083461422347125957452462591295628914127971979441382155372547382772527705813472759698246248778254779127502689271808;
R4[424]<=640'd9040644586860307109103066916626024413881146914127272889571492516922347022474973705669643456153488059781654114893486844498777613968853234329217874570248192;
R4[425]<=640'd5287344354222221341421370079156434470917695836543991018247911734315486140325169710248690910861237413886730373695892782174526233452238774856922958594572288;
R4[426]<=640'd943490606205385899446927079359932023941350293157844647567443168556599031469678876247465520769215794415441469468567832666463952303630914507231186520392658752456286535680;
R4[427]<=640'd2830471818616156243523045453202008505469035959010415996307490857657255207857816618907066218674301876836348005062871101987455910152416832279191402035353822184924109602816;
R4[428]<=640'd4052261301288176500039427513437821044754149289690841877404369350929288068448087733441271456811014017475924340857770324495352675780471980706366209416624780402320364422722853273600;
R4[429]<=640'd4052261301494565070146855517598076294413946988806611188816713815503039596147657661098111047878605358547828798313239968219528329588376516831295276132496447286348995224372024180736;
R4[430]<=640'd7091457274796073584682310491465327871499916875177418542316811663850723241294075380165179219815069216730969661754022725213024278575822621293190792640228408607560768192420648058880;
R4[431]<=640'd1872239171688811531006258708902494590671826933837671013205006277210147557882508600534461127137801475709521636323348263603274567138966329809240084986383836818012775645184;
R4[432]<=640'd2902173419177584810087374655667761293351404316292792227097304772877568546566293778927036001005618815643265353624044627851705117252671576394051347916694925202095809266450432;
R4[433]<=640'd3770276914641051565835082938016883551574082470068117969263253823175276600366548393204933766850865429678811536546577594994394900544910176176012409056207164280393902850048;
R4[434]<=640'd1885138457320525782899160419018644259971420543164466704511941419046010466742874757795453384704681061945890483519990417424253143689325307758335465696263901834543512944640;
R4[435]<=640'd13820663176836699290400854597813621474089188988507208449463733466484922088780156460943072134917365847721420297150376674638819408853639712244876477198645833775632613376;
R4[436]<=640'd13820663176836699288584373465898598048921615888264454722455470332380927974557148701134561089432341929734400046252853861840198475261837266739149167466760187896083251200;
R4[437]<=640'd2898417477601858690962468235227069902285086339769230196183485753744091066527379645530506730021673252390149862984550889876383553170872683668013465488404669308230452583071744;
R4[438]<=640'd14565683301213052609068564934792438335934889162472226406464945593728352407593428441589430685928932706012152039738077995615633353501383633346215755073550786415644639232;
R4[439]<=640'd7194662940233479757696166454046911874207525152955748096509839565227037753179991504107214121007491828185032696917629089293651443479345898177306431654420409417212100608;
R4[440]<=640'd483067277656084907224954389291648335426908052986296548651740784449803658036384293359130442978701467792180046040123543082222612563085332549407530460850296044089428047560704;
R4[441]<=640'd43189572427614685275252350037164311192940643596673558150107547665025301756099169671385756237558354994257197129900875405203018185999738458594660273111507037897940992;
R4[442]<=640'd25193917249441899743745040984883454337306724522601850936838956234254762326116973524142322904576375816035862216583501626356190838649412996844137295128362448681172992;
R4[443]<=640'd25418862939169060362096067855675084707150964603404306838861919329244959395550736448434338700057964824011527488286566626570335614783724000445780541818896954844774400;
R4[444]<=640'd25418862939169062010330406016163706905786016876307315686166757880769631452307334406270617718141508663357081509869932929664729696008146893005787820845531307278598144;
R4[445]<=640'd54211911224245516562710919433507708016225344483013908007964285590783762699259533668459969152141175422016419704350012338736366482355354478064896909341216389134811136;
R4[446]<=640'd56686313811244274424979756637685385198026312315606393283444120181204705778220222219467809118228884912364747852164851687689430594258764356957686380030279212242829312;
R4[447]<=640'd483067236715969376881842129484187352508503516501488141193986830941045971626099944734956605061775815732628388014536826632721720159910022411551574942870332206856602786988032;
R4[448]<=640'd74921965209854830353893114976975521651528110328674110446295645636295531078073058605018046148937565313708139268949537526897698693287908987189067776;
R4[449]<=640'd247330401473104534060502521057108172662176461592532326946807338744752493470925840003355931071837583690394979521980495544148853132096389540867078991978657216677450370271674368;
R4[450]<=640'd741991204419313602181507563058941570291454824163059014983526886564806459620400549202768847260599238884420531126705388107059875298848651478469988721492180005668439716211458048;
R4[451]<=640'd740650080353392514210327766613105336941552877688410087520855129046969808957545513240677429638263007706100223294799558158469436084687208448;
R4[452]<=640'd2791083497488295799976000275279077200176930848682339923977481261852836336185204142898137339594699892006276598257105046725773982190111031296;
R4[453]<=640'd2233570255760549968489300648395040819232114963418312129943281285767218421270557897454750353992402389840136450811184294112892553122075901952;
R4[454]<=640'd1571181819613545437311146000935290375595447422438189577540746050491815210670997825309991662785972014709889007007626602017448257226337446528000;
R4[455]<=640'd6245067543222875479289493122088883645844833463043344425242596689469094668000272245192282645754613237625895270228267607158008507519555786946645504;
R4[456]<=640'd51920445716931418627941055506425579560166797585488155556993696992157875508862259296461967089991829991717049723331819362644875030443311826534400;
R4[457]<=640'd84777009757886095844778833338952854877368829864727369248330697748909607935332927069258965360010164643680862533669739284285752978952301838336;
R4[458]<=640'd321787390318625379271801228040112000489524307835454329024497500821447657955492270863522153832685991807191694495152205347357170250184167350410383342934430464;
R4[459]<=640'd536312317200609564338206008910304974811771605910012576778739007226506243688965707019503691419900440306583443581099998691829419103216941462068165912453722880;
R4[460]<=640'd1501674488156690194271767992113256497504673032948576655257371864068033340902489119814366245260362954143707812125274030276923325347124705350352840071598575616;
R4[461]<=640'd858099707528810908739973765739691376685074470234581960069039409435578345349301538770113679811527987871195139966833906441990692101150623755857982390448686848;
R4[462]<=640'd4290498537606602712798093310782130492002325198791009890357605088747341440357238837772805441414798642442877310214307853618593916022940082825521298188087592032;
R4[463]<=640'd23187711625447378152385878811276641251750559684128060883314819484372569753004615980254065088388061916311718477715304884524009727637885306248657608429199320850875207298581472;
R4[464]<=640'd2227754207826376728279879934086970110530891801225216363136272812290896005848167044162338021685050462976889752523623869332752300852602939853674750510971696265611554168598669146695385408614752;
R4[465]<=640'd53674952944743664743095463100482098000120840438710242058761054900550229692075329704871876026916598601660876380097788013448077616138772442588059702449319882822244632131828005869877106124009728;
R4[466]<=640'd470120864359596985928445002916096020990314239991543428592704359952153159898537390503580370598680698112889757808377927875120104819905830701383182103344500781254486157780480744122844132151296;
R4[467]<=640'd530764071669824125085649339642764672811809057113453592337230523566602747641375130297336303839373587488330645215876187536890263119926698922515202964229726986388345800019788461615905706606592;
R4[468]<=640'd16316559141357061340560387563030983867592480381156719368408518661575014406278397368770494013017370058697924099970493187263592180360085260423730164070214017880065331213898817071503762522624;
R4[469]<=640'd2364813304596757790445386406764097888714938266854536457091169394853189100498113258748627178937673877212685491794225083203009545461261545748650877599060265600474578306257289980765765214666752;
R4[470]<=640'd17804629332869548528335610486107759507786125980306599698634556070191243773151219763854939953482451439420097925179549876311076045051758421752308127879122155210451701937409406789484359318504448;
R4[471]<=640'd285117729942326845937656398829517704632976591601273358772530245867457498383720993311279466044138444215143884612072923302307146919125497495019919867528282543457967984878444588054129446039852800;
R4[472]<=640'd1155960773273384504695170505830081040668028771333613581914299927837312415144509846221855764652938450005338535496414031291748972327791298083694214179244687173593715527078842410263323107151582976;
R4[473]<=640'd1751815407646183192811976948934752665563299521959185716057995881985366276981243400976101156301976386550289131298751733480155224789241704282224223191333993457835712023976255179217384094795628544;
R4[474]<=640'd1434745283105819162979099952413491935703925505924937604503800573307380877235202418218051963439109706255852910166716879262697817939677914865343738069406434720321712357867138328195915821252345984;
R4[475]<=640'd1140681944900537987173327972652769300603595575052243546457464673655100257734050248651976188085351992583126994490122979542809497746621874365939231060642457641880670693412764743323206657666711552;
R4[476]<=640'd1149503953876014664651149481978249745789859699365667725566678330677427670323931710860395709914305479581166274184940505298187755603341603884355204399344624613242503619628697157569241614674561024;
R4[477]<=640'd552428918611849294055718277325147603185172029935371738691954795392155422071543936517515870618394799379679054041453215691456435034894796865560698365200205870963422576726794161849521286483542018;
R4[478]<=640'd138345934588064155642400151671399778565597450066829308193754372581588358259931872165919564355584639097265209658281397423937033881484182956466962298670020582363868098871062388399783784260044315;
R4[479]<=640'd1996006460156567337288751693756555171013120456927870592141741571724426103545411691868126659200259207235753695523481301867512978982058941416814287246351271245959691947570799806039509704624636428;
G1[0]<=640'd0;
G1[1]<=640'd0;
G1[2]<=640'd0;
G1[3]<=640'd0;
G1[4]<=640'd0;
G1[5]<=640'd0;
G1[6]<=640'd0;
G1[7]<=640'd0;
G1[8]<=640'd0;
G1[9]<=640'd0;
G1[10]<=640'd0;
G1[11]<=640'd0;
G1[12]<=640'd0;
G1[13]<=640'd0;
G1[14]<=640'd0;
G1[15]<=640'd0;
G1[16]<=640'd0;
G1[17]<=640'd0;
G1[18]<=640'd0;
G1[19]<=640'd0;
G1[20]<=640'd0;
G1[21]<=640'd0;
G1[22]<=640'd0;
G1[23]<=640'd0;
G1[24]<=640'd0;
G1[25]<=640'd0;
G1[26]<=640'd0;
G1[27]<=640'd0;
G1[28]<=640'd0;
G1[29]<=640'd0;
G1[30]<=640'd0;
G1[31]<=640'd0;
G1[32]<=640'd0;
G1[33]<=640'd0;
G1[34]<=640'd0;
G1[35]<=640'd0;
G1[36]<=640'd0;
G1[37]<=640'd0;
G1[38]<=640'd0;
G1[39]<=640'd0;
G1[40]<=640'd0;
G1[41]<=640'd0;
G1[42]<=640'd0;
G1[43]<=640'd0;
G1[44]<=640'd0;
G1[45]<=640'd0;
G1[46]<=640'd0;
G1[47]<=640'd0;
G1[48]<=640'd0;
G1[49]<=640'd0;
G1[50]<=640'd0;
G1[51]<=640'd0;
G1[52]<=640'd0;
G1[53]<=640'd0;
G1[54]<=640'd0;
G1[55]<=640'd0;
G1[56]<=640'd0;
G1[57]<=640'd0;
G1[58]<=640'd0;
G1[59]<=640'd0;
G1[60]<=640'd0;
G1[61]<=640'd0;
G1[62]<=640'd0;
G1[63]<=640'd0;
G1[64]<=640'd0;
G1[65]<=640'd0;
G1[66]<=640'd0;
G1[67]<=640'd0;
G1[68]<=640'd0;
G1[69]<=640'd0;
G1[70]<=640'd0;
G1[71]<=640'd0;
G1[72]<=640'd0;
G1[73]<=640'd0;
G1[74]<=640'd0;
G1[75]<=640'd0;
G1[76]<=640'd0;
G1[77]<=640'd0;
G1[78]<=640'd0;
G1[79]<=640'd0;
G1[80]<=640'd0;
G1[81]<=640'd0;
G1[82]<=640'd0;
G1[83]<=640'd0;
G1[84]<=640'd0;
G1[85]<=640'd0;
G1[86]<=640'd0;
G1[87]<=640'd0;
G1[88]<=640'd0;
G1[89]<=640'd0;
G1[90]<=640'd0;
G1[91]<=640'd0;
G1[92]<=640'd0;
G1[93]<=640'd0;
G1[94]<=640'd0;
G1[95]<=640'd0;
G1[96]<=640'd0;
G1[97]<=640'd0;
G1[98]<=640'd0;
G1[99]<=640'd0;
G1[100]<=640'd0;
G1[101]<=640'd0;
G1[102]<=640'd0;
G1[103]<=640'd0;
G1[104]<=640'd0;
G1[105]<=640'd0;
G1[106]<=640'd0;
G1[107]<=640'd0;
G1[108]<=640'd0;
G1[109]<=640'd0;
G1[110]<=640'd0;
G1[111]<=640'd0;
G1[112]<=640'd0;
G1[113]<=640'd0;
G1[114]<=640'd0;
G1[115]<=640'd0;
G1[116]<=640'd0;
G1[117]<=640'd0;
G1[118]<=640'd0;
G1[119]<=640'd0;
G1[120]<=640'd4171849679533027504677776769862406473833407270227837441302815640277772901915313574263597826048;
G1[121]<=640'd0;
G1[122]<=640'd782221814912442657127083144349201213843763863167719520244277932552082419109121295174424592384;
G1[123]<=640'd0;
G1[124]<=640'd0;
G1[125]<=640'd7856604604333170949743877766454759612755986011919476912003707458509542094434921138512834176236971360256;
G1[126]<=640'd644889003695414346689444777971923024932903075611476636687358065354032681250220038412775185761064401764352;
G1[127]<=640'd645028987745581198224681424290572787897973484321965327621933292354023594916170530164222243531070262738944;
G1[128]<=640'd11037427093440622621436285598605659520641623359661458616588163477219863781927845948822192710631647497682944;
G1[129]<=640'd573365904994618745855007733816613264713679834614346708084651506764305079210124404513811744224823329423360;
G1[130]<=640'd5160363136974761769076649524420787146306809812950908955559829185538150831387094020653848850445074702532608;
G1[131]<=640'd5160367511476211335100498269425241381549540519289770741984702037079363651293092419405695297471428748640256;
G1[132]<=640'd1185308749101867383528343525208305352855182012758193426475207759204112866078574056471934617032200477336403968;
G1[133]<=640'd5873219911436570654128813737715762151372875389205482319821989601207900799163625007369548846695244672561840128;
G1[134]<=640'd4698231897357655693270671209046307281280792457485868434830751246077946660387637135736425620257987052722716672;
G1[135]<=640'd537521240116874746438391167318609685778272093980868742676505978066458769459245031884024810279769523355648;
G1[136]<=640'd286617334975565882569772691841493103715879322224246557669232980263960241015086220979209166717100973096960;
G1[137]<=640'd267019568481510095727395071886519216282314924123443374238858075630527062142259812707126488650974410833920;
G1[138]<=640'd123605912958937569870138845858871018598838310878637221207293148509439263890755132173207176659926817701888;
G1[139]<=640'd50114288606228369211222771027718940722971818000625283343387256134064843117656101152897133911952209215488;
G1[140]<=640'd49834320513456143684903090742647885188206612313470952151524757496444369133758581034724524225293258326016;
G1[141]<=640'd19597766494055786842377619954973887433564398100803183430374904633433178872826408272082678066126562263040;
G1[142]<=640'd19037830308511335789738259384831776364033986726494521046649907358192230905031368035737458692808660484096;
G1[143]<=640'd0;
G1[144]<=640'd0;
G1[145]<=640'd0;
G1[146]<=640'd0;
G1[147]<=640'd0;
G1[148]<=640'd0;
G1[149]<=640'd0;
G1[150]<=640'd0;
G1[151]<=640'd0;
G1[152]<=640'd0;
G1[153]<=640'd0;
G1[154]<=640'd0;
G1[155]<=640'd0;
G1[156]<=640'd0;
G1[157]<=640'd0;
G1[158]<=640'd0;
G1[159]<=640'd0;
G1[160]<=640'd0;
G1[161]<=640'd0;
G1[162]<=640'd0;
G1[163]<=640'd0;
G1[164]<=640'd0;
G1[165]<=640'd0;
G1[166]<=640'd0;
G1[167]<=640'd0;
G1[168]<=640'd0;
G1[169]<=640'd0;
G1[170]<=640'd0;
G1[171]<=640'd0;
G1[172]<=640'd0;
G1[173]<=640'd0;
G1[174]<=640'd0;
G1[175]<=640'd0;
G1[176]<=640'd0;
G1[177]<=640'd0;
G1[178]<=640'd0;
G1[179]<=640'd0;
G1[180]<=640'd0;
G1[181]<=640'd0;
G1[182]<=640'd0;
G1[183]<=640'd0;
G1[184]<=640'd0;
G1[185]<=640'd0;
G1[186]<=640'd0;
G1[187]<=640'd0;
G1[188]<=640'd0;
G1[189]<=640'd0;
G1[190]<=640'd0;
G1[191]<=640'd0;
G1[192]<=640'd0;
G1[193]<=640'd0;
G1[194]<=640'd0;
G1[195]<=640'd0;
G1[196]<=640'd0;
G1[197]<=640'd0;
G1[198]<=640'd0;
G1[199]<=640'd0;
G1[200]<=640'd0;
G1[201]<=640'd0;
G1[202]<=640'd0;
G1[203]<=640'd0;
G1[204]<=640'd0;
G1[205]<=640'd0;
G1[206]<=640'd313311928306697110311803807986822613638199025029763407112273703794759655119198407764919090136231572864649788791982975990940762992329280168040802921234664679863442740690548435188188041969664;
G1[207]<=640'd267988861103656740246423867145287360730910185107880319041818736593842818549152164187500875492935027459952124528262589566299208684288699353887509762406554247947371730687622661021772617351168;
G1[208]<=640'd459311119024592205994633021641925871462751826168338780949152408524999937200485415184519346760362554173795116240172981133535284808687500956950815233563650040595944645111872306228081851367424;
G1[209]<=640'd455231999469027732468200345527908179771557340293764519713080026408558320956845215735973425389511062869019112661787327259139131133575933354677249915933747616932825503281037685890297509183488;
G1[210]<=640'd8702164631364184029140876295477713663157168990651150485354136344208865690277860045195168207992511065580124317367840887061049600634020064546028569235343724814188716477854459548133060771840;
G1[211]<=640'd8928421161030303780321715324073127003000968316841945920997478811977506108574178650495612941367778629541695961514758865444443592731252990709418564307146995669129238524099904265055635958136832;
G1[212]<=640'd8989336315162131331140063071623692371762926782277319709476611382585623268259494876113503496518513279800569773603677691511220387363917993092166919658463383915499773903646914806751677749657600;
G1[213]<=640'd106601519710292466488971541735361695339222342745245653012235616923935171069415002171119166344765869784759587183840588051400306734297725437701382184760856647128412208072618636373867213357056;
G1[214]<=640'd88109419352385881824206623572303431630283385935981590624916579503069233233748313665713336920838003579676477462191133815517593520684107863773194596183487924038169644986275704493504316047360;
G1[215]<=640'd32633118278662046878287562858316642211869691329553823795699297245112837686322715345281590873244188078135788707546053033639081168038122481491230909101780657524947994759919597041465472057344;
G1[216]<=640'd17404329748619453294258216695510201226554577810894329362375733702790952754936266944239217076442965156914705349414929384545626893576552249518431506860001275696403347280703382441572066918400;
G1[217]<=640'd784178183318689112868765898469809193051511296717339887724197064605486354861853129915951577777110562238387831159168796599620444531552087373990407885855659995846100315216932581943140425370959872;
G1[218]<=640'd2272413717958295978214458277023807115325782775776022248590344460557413126741852426664371429640105052489747052595520628442611715819368495296518012665770827493485030400650277525883008154836402176;
G1[219]<=640'd4559795159500405005341383745848705491822826715159880689817565956640738571986235814246918087861646807566901220944412668512398915194583249909476069398539854117890083405337585890456380955414233088;
G1[220]<=640'd4562440617622195218639239336938782695720880831303093936907043054234421949709348768880187051868712660154222880455163570740294269367377909089059654072692454514430764407749007580507734093410074624;
G1[221]<=640'd4562440617622195218640930072105102746246685047755376681370173834941168515021261309302697091510962348638221560623023179685093818127359248480349219667747104368301496251959706394228331511665393664;
G1[222]<=640'd4562440617622195218641111222301494180231592642375264118276937847159748504161823367205108881610741218169234457865671849841463575991963568722070004587058659568584851149563834249943270012116533248;
G1[223]<=640'd4562440617622195218641167831737866505068075680726631371055776800748403055085607835349530173818435964565738429196699549917870703476196900078646174067622205952622818418666118700631846561098235904;
G1[224]<=640'd4562440617622195218641171546732128478245430839257927892528895891810740401818414940152162012874814034754177120555145486710945536394411893246608775919031836092140761626594823920070377955175432192;
G1[225]<=640'd4562440617622195218641171590958250650987666220969255353467072756324804170843011452186266281330920354533674384883722098966129344785321085666934206298743762570432107738485294221246316422709116928;
G1[226]<=640'd4562440617622195218641171602187539921514534640823381227492934617272734083368454577579059816740758679300879023137085305911107797140787547732683978819641804298519992094021474204285045086722457600;
G1[227]<=640'd4562440617622195218641171604311702457469172610346825939213314509214747357246659884568837982482925282052336609976440267613773728213545914458988709479667344986197224461372343433778251642540392448;
G1[228]<=640'd4562440617622195218641171605700073405323906491108462711257349328013878355597212965432505169578059804260843873110092262239683911729224869951919578537858742390718308247009226318879978497735917568;
G1[229]<=640'd4562440617622195218641171605700263203249613782205863364634962841387446631914608493840550698321534191742967122006729679159317530542905158955606377567394297630641221104798857600892485597162110976;
G1[230]<=640'd4562440617622195218641171605700291324035128799732235240497696796876326615030739031502418711239400153922494081086525186072560477505555284043273579300441515573737906047184228562104684800311820288;
G1[231]<=640'd4562440617622195218641171605700291324464178653490399871975392009007896097373139941175314621992373945250252883911169622304166366304038141860833527790222966387988516158423110887231178178692120576;
G1[232]<=640'd4562440617622195218641171605700291324785966043809031348112874634813116786819823218381340226177164434486448952119481262336423589186062640995424053430772582311455753364487607069491660392375517184;
G1[233]<=640'd4562440617622195218641171605700291324785966043820823265488482663538540062713996833519607899287882700738129875193428458290447083693591886714226177578367357258791228036712318107804330684951035904;
G1[234]<=640'd4562440617622195218641171605700291324866412891401161730581308436828389863872891320087722417132584161494635409351948800312364018605522052086104435992850778829983942819016902685197244968256667648;
G1[235]<=640'd4562440617622195218641171605700291324886524603308562620431933443251225021983283034041605399769829388263654683235560607732845892533253631639893451664769815630750200134816616739458189325080985600;
G1[236]<=640'd4562440617622195218641171605700291324889876556065241910185193022883412596503858119322405837495173124037656050230171185704348234897631296164968910023698240585855699275609712348022177326935572480;
G1[237]<=640'd4562440617622195218641171605700291324889876556065241910185193022883412596503858119322405837495173124037656050230171185704348234897630492695946780529252141155107705052682643749729227425250803712;
G1[238]<=640'd4562440617622195218641171605700291324891552537650658136988897854644010563059147059951467758323016871557730542382596535041468460440489867205778705293916892503573506279734575995541940229267030016;
G1[239]<=640'd4562440617622195218641171605700291324892390525546383595697509479802187317088733198531299642343845517320470129926464236085286077740275503371977589207939090169255257016017550175513277101158432768;
G1[240]<=640'd4562440617622195218641171605700291324893130318317005108417396301947392592466920075590789511729408734956706332185224909279802186631377899161820005028224593108916582151396207434985445370145800192;
G1[241]<=640'd4562440617622195218641171605700291324893199264106683920905533454755382023774063638613884293781537226781146857003311682737614415507699073353391310669467416351801695336856945659279567790928822272;
G1[242]<=640'd4562440617622195218641171605700291324893228353808375185447542361031008128414967126350816903048709392749359430067322700841568944568089860219962800792544644117615293496160606310908054866029974016;
G1[243]<=640'd4562440617622195218641171605700291324893228404955103433824759079987097141346203879735848872471596728425787056569413269664608864619185052813651992767235414410897598307243446078318130596721721344;
G1[244]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998243518165479071942623648792974195658272695869732028416;
G1[245]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214183018159440957466004834783788439699968;
G1[246]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214183683097957403738169213916956753657856;
G1[247]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214183682784847707441707772724389513003040;
G1[248]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214130187848388438345803321351235325394944;
G1[249]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214159767055455326655389368590118009702400;
G1[250]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213949904800324066540885820982294660515840;
G1[251]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213768471754361423735895291916425218752512;
G1[252]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213811843008030157571299707572587627347968;
G1[253]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213699854251232106408629362375355407532032;
G1[254]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213766076813129948727513099929569531527168;
G1[255]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214066151240457114539795810395382907930688;
G1[256]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722212274704014911117209043633822896776022016;
G1[257]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722212614820385620127775702348391542247456768;
G1[258]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213231292294930482802909124182595979968512;
G1[259]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213709816643780217196839984627690157118208;
G1[260]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722213622007724642592104428891580632953782272;
G1[261]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722211256155813746072058724012506170882819072;
G1[262]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722212523045847105468319980954112594920095752;
G1[263]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722202553720590021307157363260780387797836032;
G1[264]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722114980099592035899225944848989123067772928;
G1[265]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722125584971261729564299382171262038225076224;
G1[266]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722114782293983637351823933446960578619768880;
G1[267]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722127048246513689366887393187776226622703104;
G1[268]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722080764922636767181393983866297732349625344;
G1[269]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722124342404553064474057487540397929299261456;
G1[270]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722082110431962186686835370983502372551016456;
G1[271]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722153612129732168348040553018048486662357504;
G1[272]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722207704208238708732488350566188081206673968;
G1[273]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722167566519606896863652761621469815663497992;
G1[274]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721797667607160274639288046445468090703124742;
G1[275]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722144576776659895024958976554344328442448128;
G1[276]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721450423881841699669615362278230429663398176;
G1[277]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722191557879911145882030391286446044173447432;
G1[278]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719250749240255375983464134326451300871780364;
G1[279]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722104693473622308971315664290119992714797056;
G1[280]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720817212061827106536182670219579659791835136;
G1[281]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721481932235710473170963404572086893099290113;
G1[282]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721157749605064336189493735271094106414270472;
G1[283]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721941809349342677350830750588098061763888128;
G1[284]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722118503953295317751347567552914258502112800;
G1[285]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319699282718403930853294125643366146151626723716;
G1[286]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319699776521786076725051430616728638931305785600;
G1[287]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319688694200172779477766554959799357320653180976;
G1[288]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722202828522998241280802289084114997576990832;
G1[289]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319532637392478827933647679540906175624889000960;
G1[290]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319627434530312708105248109275830760979857213192;
G1[291]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319652501770000723648316016112457681174933864556;
G1[292]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319687784694190267611790803287721481441082618404;
G1[293]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319709005836818768659581600625084285651684192856;
G1[294]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319597735992417730640147524422105734715972567618;
G1[295]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319704425318823092208692737258775695102791129280;
G1[296]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319612189226417260766016753715309521609399220328;
G1[297]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319713347992946084712452087202222552866472098604;
G1[298]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319697632297860641221165298606686137948392978708;
G1[299]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319715318043977135892269762072238106602411432192;
G1[300]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319695646134703842472440153818376074643682904480;
G1[301]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720922800764237520156858877321594117184610704;
G1[302]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375425444049190546340543400134240147430031395457970103997970212;
G1[303]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167191025287729928084630270389813777970588918684117520184614134514673726282552469309072705067719202583108049059387268444780;
G1[304]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167169589442003439202944282419761796910784019610258900542209387818122565223944208463112359953017334543485705278995595540568;
G1[305]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166564356157136415442331545608023544060419023683936768250711576003827899691057367009044971047505777841175771352668691781698;
G1[306]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275162049201463079179280438065844867887067267326201455591786138045564644151014980328933680885515862567273760736840968768387146;
G1[307]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275156899812337803157707737652906999018296705664839284185377959971661727930427743957172327347255213879205795348904982919305348;
G1[308]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275125932396597839862688035125525892647180810319955750924550986029677223929081561100447406079634971354490342258811961404344323;
G1[309]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275002580160764118474072157422553191623604818998629456042048076802429711979375279119933972163466601376466607558961332328620129;
G1[310]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275156224501324744261471393539734416719326353029795535290926532571364367509948170164034356597605233739940104879000834117738545;
G1[311]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166080834365950132447865906606669787770241554182498271541406155234811498601592500926517755643252789114521039253883502499888;
G1[312]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275164695775044134473714595873789069539457765391187662855493923449918656153074838476785160848277662081210204184944525860194320;
G1[313]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167207416522833775118479628795831052913881293016566527069834926222255363029669212179763079750011087471857140669827224756422;
G1[314]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275162074438371542140335755986067477795315974635437782380826164998151958896196702179338351723342489683919490903875839105728710;
G1[315]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275162364446832682772231238638314383038137283675279691450682625193579854620600621681013698712964369665599841276448717192086084;
G1[316]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208366498087649813788587882957434643481671737020355154001811087733773624886972124909777245627828535938937688557776429600;
G1[317]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208669998028560728666359368819883062302996480584021686606677333439452763175153451423680328451632044615906965945721831488;
G1[318]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386205312978440073940369550141924008404023980590268689722731364265093397033541242068149390970064834200110040367168;
G1[319]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386430763892330380474939960351168671723766720280875357595074132306744133313239191879581041281319056648837221582336;
G1[320]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386496519501048257069401691674887379167673002900263163333733932077534579801448565434258761562404890058127949959730;
G1[321]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386503635367191693258767613261747795844765119871069379424886064923069276550589739977944093899805174729234891681945;
G1[322]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505837340878538976487963366969842819125157653212785634563280061570343940750626786702581418776300687245108338761;
G1[323]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912739645539650088907571978275040648687722901927070582310167942847236229700674794166845690739756415371712224;
G1[324]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912810197499028689740204355581669908517795187019562008551292859805469865807055682353994412101516390416533552;
G1[325]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912810757435214234191256941822387528831467224193747421799431602269826934630406348521708919016604540669816870;
G1[326]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811274173197964177824068186057120144857430489393594228461302908130123867639196911911127073621172352726630;
G1[327]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317367127804570467753444438654695398060060704800514667469252294113081144409755801103274755917191464684;
G1[328]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811247379376585585927995571473632984372424597519073508683500867096281294670393729888056990588238325897224;
G1[329]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317370463198389254409027062208615233436168291065858317502430770870334209078690085583275711375278090432;
G1[330]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399257415727664530573536290932835601204314370578580485240137821837689841947240321583538867036889;
G1[331]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310682125445970789773677252681040654406515731857799178672312129654966474395;
G1[332]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310676732719290655270284643651673458914522018346975786830738944505320859173;
G1[333]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817792082077443838416964060770643043543706307101491112984522880008706077915921215686387644052673512854361901152625675;
G1[334]<=640'd552483043540187702257329374127769652623789389549630304093574093964365352279175777272200379495462942941944967174927447760268787085521499251715314460028262170293462993270246366730858897500171826;
G1[335]<=640'd2352508443461444409611854109189212714398070949050038714204896142041813758091974277417111293335519628010862440873884616269565395557594364053286754204806724397934295253686703518793062741057497141;
G1[336]<=640'd1220809305887188954987969746056523264668695909166118575174510497953516988100759378811152451465781019081394524241371941018653844411354947854928813111347689986337899096241027914677060549565905014;
G1[337]<=640'd1211967906374890084248720649469549128342685166667025449088335610109077169585203012415793398013673686199133056142680435743276946591876701373908921769012924445404818056406325459032397327459813978;
G1[338]<=640'd17787292988752540970425987999352579119887799829795397524792341530852631625865517417545638778260317913268290808508816742416698434471421547225673351712949099098974021148698609235762643005217369;
G1[339]<=640'd1358895530055390963088476897804922810104619777090639068674129900788965983129476931072970675037099460547809432175343289266257784031464452332234360453815214741473113898864678065582084149991715427;
G1[340]<=640'd17827472515633143767907657968001860266608028889965212035718533081019215754361871168004370943231677978270570948505792317715775796702564707288582076588780219909900646723395937071618930036843068;
G1[341]<=640'd3635701393791342547288792320952301766258784092753926824448566312470555105428358362524258050347358169336067889753538770322707712475809406745267219803158565157956730346117737397604215186361034812;
G1[342]<=640'd2156579201316356737668750359528068344929437221326533070671207559544212858605998303606570851923908801392637092210460166195075063263543020602307870168767245832012818948735338483615555366474095628;
G1[343]<=640'd249551982100585350580163723252615460060049274258359819658698089286417987766348345590267299061104316008476496718677457461127030053149052549694298991463428630292037490649372274242623168482253390;
G1[344]<=640'd35652769490047710057779083382709681621718515766520214148679641238848362655742552285222482241858065980858851336357973138019627689488466993095905596147265631450570583626502424759950559111295600;
G1[345]<=640'd17826384745023855028889541691354840810859257883260107074339820619424181327871276142611241103431027192164834877461761065410470343887933485202384473354062150970900198707931140915108598265677865;
G1[346]<=640'd17826384745023855028889541691354840810859257883260107074339820619424181327871276142611241085933021393646606337334485750453877350856865075079459398866583258341938622286306917980665900465389602;
G1[347]<=640'd19814829418803669954006095402106405919612658140191976474626200415147112952678982561252524303796180024070309343201397479428773083188900569770923080229680040270948913982912375393580001777420548;
G1[348]<=640'd22068690121249937199543020614730718231066184033169456451318420840058444641191874912780709703336226334472046753321625318645805318890609620586705033833308557046102626559033395045827144940132641;
G1[349]<=640'd17943974447529544730402627003579904945201011162779930125880791956068346520327593275471075026868540818710615558051699178666257164866324664181024731522361485561066134118411313555817575155236905;
G1[350]<=640'd106932205425842395961448104511667716586385540205487165482536106984652009257604449665878261228951562570763930626695899624367248088467086999358041877336493011152557481474130544691199774375022889;
G1[351]<=640'd213864442178452579189952549312758600109192189979437161279349590486521507974063517159366394819244034873929252833373623650788331949903861574000544120755080960938949184925751757658894305249726763;
G1[352]<=640'd89110171765330453673071524406157157530366946924553701369832354661607111247746686501598990761777225762586392262502995651726990922353005330956623799462035742198600814847482681816359946011281664;
G1[353]<=640'd213864404216609397282188468361995259130604399942072805609415610876250592497543594208378322287961787634875931497518949978299195024990886634828377282200711453384447770603964930722950326868510976;
G1[354]<=640'd213864420951605686579233070042536173397057321975268460243163628558736603204938036918916078981109468789055488462749049527899779295724413847259235597623528742774363010546305458414046268163620864;
G1[355]<=640'd213864403951053063386536537181755317886813098899552677856796746743793643770492086188557130891168892319832992179075148074761487192893458308378002939113801443910847549752779363480467585777008896;
G1[356]<=640'd213864403951043693332244791461741309206387084879571227599538263758038181686141622277018234868857785133374243447542253425471256111980176083948196897361704335306143415229603581624861440366084132;
G1[357]<=640'd213864403951043566702943774755236936366370592017946549092831933627972386549698618547506297271048925983415327038963207890289352171859101475299172603701027647729679999918391870426937856508297728;
G1[358]<=640'd213864403951043441058616759227754034170208857603021270333298999319558124773983079928088309475514766698219188496441723587839319851920941124028744683154554378235726311332192664331854963407849472;
G1[359]<=640'd213864403951040401125000237620511548719903057088161373186381516685831279052620557643828245811823449381702910600223873600033882053537430605162746006178028454993144025975896235007115632578658304;
G1[360]<=640'd214412640338121925339041193445694274201962037358388047315545048274278322806556624459874713672177814107053367483710110953592399697793294318987507440932167413096222001569981318942547532685770752;
G1[361]<=640'd235949487115300634773081896752335710222757643093273017084350995345694745624487002373123505318932719171320110437701682830546161757000089696924451782627693077014127843730468608097270875883046912;
G1[362]<=640'd158174373878496731298704542431671560981136220758180333395070426223417094505265505576407389431666979497967716935414234502746044452180586386490672703304813280390563870287540544315232251480637440;
G1[363]<=640'd262876054550035517074112469285017208950057125267387170538412639015930609138877851707782002813139236208494630259450344373758745664339644252707642293543468247119423587537649838317984278464430080;
G1[364]<=640'd169309823844528833803738883974492267108581811167652608179099078993059989855644130642740796093482106717921143098383080893314415021460212278343549461659154331983977822663429582768324338316738560;
G1[365]<=640'd249508477649869714820644256461793160890866785692538449232208597931959641298372379043208043152359920271122640179809362037389510159652212212090880977266680762518238157409865218875964190206459904;
G1[366]<=640'd213864408183546281132417736699857177250080290059389529833793190526786436959754839133047052751538005996224824265869846838462387097673797687489249188639542368961341361168485842418126502085263360;
G1[367]<=640'd33066452189520412638145750594933764169347068896536611239870907618162729113884237510647641944163920246255535807597967088743110318713581428969454304558398678526102983078643423023990784;
G1[368]<=640'd6457278377941271757216330441264760700712897713549705477192735743892107259615990940904054358504426825775401558236344542459320459278526644853649558299057113293275859406343820416124928;
G1[369]<=640'd26086432104171281416431683347155889567299536128265546458581483119986644646857687426044790057824687740116781460792216595022926493846412879058664837204917758526987189896822729474048;
G1[370]<=640'd498681975005706119718415443603550458209022701280760120740941217579021625809595699272531790780375824423490652465807201670177033402564091709809379360080753009095633633265252827136;
G1[371]<=640'd134424073200632314264243522963138317429612392961260708681273656747331527582005749120878897595083736055198279923117109681201996137013021675765006098282618757199668704584589639680;
G1[372]<=640'd3214419659867800372223267764855257974434770652469545324097688974161472277422284446470995378367437480965628434352797182487544723703303849021129214820106142038254443948815810560;
G1[373]<=640'd31814503241245648517869241101093238211037236662470666513675487398586385230280889551289867013389016058135324265727212478907860184024756462034110767510790921051448693588230144;
G1[374]<=640'd14240811337467453353817160855420349959722467716915775484722400665777604250043735808994121540395556679360352406957162114264537806967286271322355081070308966152410369097728;
G1[375]<=640'd4625315276569600435850153138487010407025838809032380927394481921881458025966916954634854090431212573210998788213197731811480684056193088069219541597457881968781400473600;
G1[376]<=640'd6219298484494922147767102511535678781180038836403045141666350261149854808328520389349823421304840125968271441850929663885675359301369023635791167926954556406825484288;
G1[377]<=640'd222246396368841369480581681761195929635717682305948900112495288670472019629516030720749335167407759770305585095129655050594856680599024767590507470455303687553155072;
G1[378]<=640'd8042288943634546926681745854549143942737816105528798614696593507125235632285197568440065774513732688971824444017473398730140011953639833621979316523469019759509504;
G1[379]<=640'd54506493473811290887492686403752511150351043915146240052750576885099601396671665391990330702801691968195348330450476794143304873079872898023696644934905435783168;
G1[380]<=640'd24150358220713734752040845208999901391118450915055709085187385447491648812305550271622825000733043201471689252403692293611533253841309212091388601284239720185856;
G1[381]<=640'd82377624295820163189945864115897164684202963061206335262583018399775145389067764591731230514108314900953979434172378784312256296908477983493883314754906226688;
G1[382]<=640'd80146925515664259041624429909697491993041433969265642683377937561860051458731381772988533293119192159132189149183479565815941974483172098710552258281472;
G1[383]<=640'd94903155409552653219896978654888664062512640287280996341893416924487618845549636410547013626296083537039394892881200885219567546335912978332661860794368;
G1[384]<=640'd50833454537855917897491505520556480922396135233496363376469383791601698252359607247831096929680257277997136291987576893763248991810373547247522755379200;
G1[385]<=640'd11388138711552743048282475217503546880153216693526359950477921944356574431825851899402933128484325360138392795913318700501498089961463929954891726848;
G1[386]<=640'd2403746383743314034799848031665627212899254217293303840008078705985847618747429646165201141908358715606687464156825015176633829799177474784417021952;
G1[387]<=640'd699271675270784832866953923589858941256048873218119811162685942861755759984363543074034377582063078309844035423782777902099144774478256289557250048;
G1[388]<=640'd156087427515889046846056386464406610689191669784131867802376860757207525103272814506226887280659783852528250784833344481153690598190598415726936064;
G1[389]<=640'd37460982604473318080606298218668852224751276303483189059570178737492045377006354207145494486563605452218253351452467535635346966304956720502276096;
G1[390]<=640'd9365245836836980432746253947369064100373936087978757373440584703858683969238042111729668876131391367126631781794857119458154272973682555414904832;
G1[391]<=640'd5463060521265126663943887134366456813987168841791878890026903649916504694909687191218902837067966501023622511180714802129622241375467007671009280;
G1[392]<=640'd673737305887759676150440562763779920458615381183438664442178194697370582331723468400725865273546992727373186386154546405289889893170448288448512;
G1[393]<=640'd229304429753450354476889534457514368756873237972151519432364351696609024582924643193817241835337661382674512915652871234525089564904858220232704;
G1[394]<=640'd381072821083495145432323880705459263017025753860902593171800056510026570651121441827778136084913325607556128876129234248999296809337299664896;
G1[395]<=640'd0;
G1[396]<=640'd0;
G1[397]<=640'd0;
G1[398]<=640'd0;
G1[399]<=640'd0;
G1[400]<=640'd0;
G1[401]<=640'd0;
G1[402]<=640'd0;
G1[403]<=640'd0;
G1[404]<=640'd0;
G1[405]<=640'd0;
G1[406]<=640'd0;
G1[407]<=640'd0;
G1[408]<=640'd0;
G1[409]<=640'd0;
G1[410]<=640'd0;
G1[411]<=640'd0;
G1[412]<=640'd0;
G1[413]<=640'd0;
G1[414]<=640'd10086913586276986678343434265636765134100413253239154346994763111486904773503285916522052161250538404046496765518544896;
G1[415]<=640'd3782592594853870004378787849613786925287654969964682880123036166807589290063732218695769560468951901517436287069454336;
G1[416]<=640'd315216049571155833698232320801148910440637914163723573343586347233965774171977684891314130039079325126453023922454528;
G1[417]<=640'd118206018589183437636837120300430841415239217811396340003844880212737165314491631834242798764654746922419883970920448;
G1[418]<=640'd19701003098197239606139520050071806902539869635232723333974146702122860885748605305707133127442457820403313995153408;
G1[419]<=640'd2462625387274654950767440006258975862817483704404090416746768337765357610718575663213391640930307227550414249394176;
G1[420]<=640'd615656346818663737691860001564743965704370926101022604186692084441339402679643915803347910232576806887603562348544;
G1[421]<=640'd0;
G1[422]<=640'd0;
G1[423]<=640'd0;
G1[424]<=640'd0;
G1[425]<=640'd0;
G1[426]<=640'd18788340662190665823115844774314696219005460391266558965658327772257672200916867547709591987078149624255479808;
G1[427]<=640'd0;
G1[428]<=640'd0;
G1[429]<=640'd1221462192088228855580650243104452027957471917384428846706397095531617374916413528953842253901432384865005467699511296;
G1[430]<=640'd0;
G1[431]<=640'd0;
G1[432]<=640'd0;
G1[433]<=640'd0;
G1[434]<=640'd0;
G1[435]<=640'd0;
G1[436]<=640'd0;
G1[437]<=640'd0;
G1[438]<=640'd0;
G1[439]<=640'd0;
G1[440]<=640'd0;
G1[441]<=640'd0;
G1[442]<=640'd0;
G1[443]<=640'd0;
G1[444]<=640'd0;
G1[445]<=640'd0;
G1[446]<=640'd0;
G1[447]<=640'd0;
G1[448]<=640'd0;
G1[449]<=640'd0;
G1[450]<=640'd0;
G1[451]<=640'd0;
G1[452]<=640'd0;
G1[453]<=640'd0;
G1[454]<=640'd0;
G1[455]<=640'd0;
G1[456]<=640'd0;
G1[457]<=640'd0;
G1[458]<=640'd0;
G1[459]<=640'd631873750011343120187508166102022593913370572403294667525865865216;
G1[460]<=640'd0;
G1[461]<=640'd0;
G1[462]<=640'd0;
G1[463]<=640'd0;
G1[464]<=640'd0;
G1[465]<=640'd100433627766186892221372630771322662657637687111424552206336;
G1[466]<=640'd27590906046292506828803208781780371200385814899000868864;
G1[467]<=640'd0;
G1[468]<=640'd0;
G1[469]<=640'd208419393557760884736735195692442048972148520616969895936;
G1[470]<=640'd0;
G1[471]<=640'd0;
G1[472]<=640'd0;
G1[473]<=640'd0;
G1[474]<=640'd0;
G1[475]<=640'd0;
G1[476]<=640'd0;
G1[477]<=640'd0;
G1[478]<=640'd0;
G1[479]<=640'd0;
G2[0]<=640'd0;
G2[1]<=640'd0;
G2[2]<=640'd0;
G2[3]<=640'd0;
G2[4]<=640'd0;
G2[5]<=640'd0;
G2[6]<=640'd0;
G2[7]<=640'd0;
G2[8]<=640'd0;
G2[9]<=640'd0;
G2[10]<=640'd0;
G2[11]<=640'd0;
G2[12]<=640'd0;
G2[13]<=640'd0;
G2[14]<=640'd0;
G2[15]<=640'd0;
G2[16]<=640'd0;
G2[17]<=640'd0;
G2[18]<=640'd0;
G2[19]<=640'd0;
G2[20]<=640'd0;
G2[21]<=640'd0;
G2[22]<=640'd0;
G2[23]<=640'd0;
G2[24]<=640'd0;
G2[25]<=640'd0;
G2[26]<=640'd0;
G2[27]<=640'd0;
G2[28]<=640'd0;
G2[29]<=640'd0;
G2[30]<=640'd0;
G2[31]<=640'd0;
G2[32]<=640'd0;
G2[33]<=640'd0;
G2[34]<=640'd0;
G2[35]<=640'd0;
G2[36]<=640'd0;
G2[37]<=640'd0;
G2[38]<=640'd0;
G2[39]<=640'd1901723253132729822027970863076119870813604833725471934611447705983146550580418757496524795109054613331443048355345843719025021161173040037501660228261006990745203113984;
G2[40]<=640'd3773962424821541352241554580988268890916921220416440428376206300245624162392148852086126725177658767541468375030763844899770584629924792632561434251432696043649395326976;
G2[41]<=640'd0;
G2[42]<=640'd0;
G2[43]<=640'd943548417247645218133907760666890987596116780712080286722786919770514102710948841640665280967231126882881470241392601968444979383700011259891362322278248128267887312896;
G2[44]<=640'd57586096570152913699974892898380567793532123114264532903689671329431521032595044740083720782129802971518987656109067457577065805510327036019308994315074097345724416;
G2[45]<=640'd5398696553451835659372646209223178230643636541962299959720906687134205096805785444382848823324669028579905092760225074147849919266593159626810218217038196626161664;
G2[46]<=640'd1886981212410770676120777290494134445458460610208220214188103150122812081196074426043063362588829383770734187515381922449885292314962396316280717125716348021824697663488;
G2[47]<=640'd30191728191620615894389286635352600317619266529393080559276102246800658014897707114211383843281661205233232759739938813731893465572301096224009483665958725886243835478016;
G2[48]<=640'd45287549097858496226898654971859226691003054644997285140514475602947489948705786225033520702131905210497620500369166138797247015559097511590737211017192352523792743923712;
G2[49]<=640'd241533595188578646543459493183249209018682958106652187416077203215719946393097526533512110411370161122653976001968886073585317416315186728483931792091692546793561300926464;
G2[50]<=640'd241533595188578646543459493183249209018682958106652187416077203215737864351034948967196569949614708676878949165946763269864517329122897063453373079654739566739734157852672;
G2[51]<=640'd112472844863579909570263462692149546471742427957547915827518889315295939516787196757976017152597271428748022765838022378080206651387357492225212879521629096378368;
G2[52]<=640'd30191699511045175681512346218169613819484916235073951384557566229483882614433130333476210559397287292929018428994133525036187055119604992447848966236674447870824258994176;
G2[53]<=640'd241533595188578646543459493183249209018682958106652187416077203215724425882581882141933225295931298011210219292963355372655117394517114312226292113982454301780104515158016;
G2[54]<=640'd245779303141450286491306093879816682380463357771409856171921302784886400822245369411479245907160092181242836145013285254851451950398774703467278319235933232392997842190336;
G2[55]<=640'd94821727527122285711321918037529694547938926092008865952620148137298094023727970131157764059182272196801491841575976919889949212676951459207298717594428311944968695447552;
G2[56]<=640'd123680307819365779785565640862950558313379770095669165401472765132349665169959150914799158551154061555665397435141489928820669630604205684395321133994701439408079761049649152;
G2[57]<=640'd123691618502340158195604159540227241239197554476574956937122118248265532146088809917907696665879844329496343487814368376144062930595296443713989629368504786842492096265322496;
G2[58]<=640'd966135302153061689825002280206393209077879404715499738738791153244321140807611855702133368941742300413947419961871663311445506305724911647050358109389512191357583974465536;
G2[59]<=640'd1328672491643376705304319143961487379043069749784219261379043574229532437673683005150430278216367289990533912541327073260788722805942240330468971769176048043171576576737280;
G2[60]<=640'd977456273427966180654057808412012811721331920771366734191627017573908791917472804984877164516867171833727044851533429418893081003997279723326149740691424788053548469321728;
G2[61]<=640'd7547953643173190766710376318793279134453264493331536479147672915071404686308418024236892969198647892719555484316302762711266649155587938409748243481202378323107711549440;
G2[62]<=640'd845368965901221244783768921571801663400118244268809909695626809425406120017502834082212835398902437578684305683605201200564897091521208026463698652450207311520738071019520;
G2[63]<=640'd191317262220548974119403460150175902760825312855507354451765230402747119376628716831892112821663507779380910340699826662652200083097172097194952896696677114400179068094906368;
G2[64]<=640'd56503017277167885077315901968766902060679328715087424350659120829588736971817048328622331919642531072166440554948368625243657459943866251726356282389949853851196713861120;
G2[65]<=640'd55674180589016146071674003524552998090997690109902789869352329026196712685050118334089431411851086209316394529760618676923854208387795526562026937770501178622619414429696;
G2[66]<=640'd498274469296377815030202032336310598585961457728355836734915844251117791473317089247594943020006923285529366041475136457890413440169440908382717014620154392785264916299776;
G2[67]<=640'd30675663620200135418787855348310084069531412335989422901791898263804303033191538392454996384515311468001488135391369024693661825521070868407595929305127178973600163355951104;
G2[68]<=640'd909302962773888334745256282156393699299937425977425469173863103769644318123025383077724687166709490180637752362785314251809272973192465833837525412789209028990449699782656;
G2[69]<=640'd429340812938289701802719999055420129579121594624795500325761599830829425687320946904721048970803343997522156783453757604151132310873260427853122493358479195531141827264512;
G2[70]<=640'd195350118199295176109552792838509945939054026642618882130022493347218987683378895500580465910769069460627316148500877207070547188610384084316043689141653203394851197943808;
G2[71]<=640'd193363628016719766687403835018815621998757129951234270881729669415065439947127165415193987183635688650306818466607058348359998354568769177405972271239325783594252153913344;
G2[72]<=640'd124395091091218982335383262241573647462503329047571521855510652895787853962072238785764231288102314124227404534643184394661167971296796162241234790452337447830457455761948672;
G2[73]<=640'd14520305658612579595436662078690854212238330567706714560784052053581005200776079772393522225463343811912241792161218043748926884547775129944231342100897989763878696964325376;
G2[74]<=640'd11621902516376937136895136244720472989306233873157651510684066040457597654089813957590202217905898720537549142172442231636802614899386348937566817089074018417177711123365888;
G2[75]<=640'd185863875460008890872681288327051028846549831269385311696469901702825563366236329932985980831895654094805269835642797049957930503462884540955888688922950244358698467032301568;
G2[76]<=640'd7139865162446049003352700960437419652583717236157389876447154626967343559576757745483387588466314499683273163935530656604588435526477451109657260300948126417171627982716928;
G2[77]<=640'd27441424281483622907426142720200249588853133786942257467082857766525740208542499887540958447681340037569019817122946399435585480344852666279756846801984768383112060646457344;
G2[78]<=640'd58360554937439985127920356064627883498726986992607514564436952872689207182397723088912400757799078038454798478321276999587441828896583995007458262775161778527479501890256896;
G2[79]<=640'd2410647982928843633051246243335853256645000890478680921337320899924576994866471481884946450391422302227808312938987866763687301722197917391670710506117384136687235425632256;
G2[80]<=640'd3290895227245222698135055935625255195410760850584187292220882071759478754419113467105137846260805169525450500392333219441789714390240889761878413971634933152826550608986112;
G2[81]<=640'd54477147602298510072556590823779940359734384220430331048337215376739184598598627969250702502342704426306462908068247930906233869056028624606031076088756145140550686400839680;
G2[82]<=640'd31929235472922592617302321926813526629433726857026349022798414046981171885451887876662389430841445017294641017808191491409180262497152073675780988981784897757962419122986811392;
G2[83]<=640'd3807928057851881784033122648545732773271710819804381613511476657797217370687599516737874054577936848370052515365277537618409879182383079366934489682078607474513985641906176;
G2[84]<=640'd4144490055690520277056032164647398662812935769829116603034424637819355775532873146915185339165810631295358156016800942362543558978168121177348607757178305659079473663114739712;
G2[85]<=640'd59716350938557454201856178447487324658287511604739588262512757192442475608829846362676597819907063184361427908232054907473842841147793775818788555443975351882077572807262208;
G2[86]<=640'd30792702914725161278276904177462638077587703261494587226031040781495488045397684260605920670061056923969377785733626545279073188208206896938191293778630909478199434785325056;
G2[87]<=640'd125586147610786429862342796337404499774913793817060690221574225633299447259210721909813335710453231040364234422075980087516798761636383051646999726527283051585930315209637888;
G2[88]<=640'd247266244111882512939133133545312789977917330322113560677137309284642155413988829832915807932938527798670058144295473352012307418936220301871333700052374979208489984524812288;
G2[89]<=640'd30855916785340922095926950252488879686749421078608065844332878334195839686865723527292584333312130470989747239344340617047124717003862206779134184417015997489677362714902528;
G2[90]<=640'd251164747296723220074379940472358178991889668802039087130070820258637775167532603859516153873362101672088998913547666083119443633161906571086335766385377763530243829779136512;
G2[91]<=640'd251149651447023933908970974255607294614794025787339738920000413233193975205701892596322074179460013082571589766528768653529997884199112870293446171187186246368448993554333696;
G2[92]<=640'd63366776477364887219473458056956824574724621728699908355986211608555007098755050018163017365086161695831306123311664128587163073440182810115735079478332616568602705197967343616;
G2[93]<=640'd49755920608847201187952655595749265606694736214630585264709727264681793320031856423935185190479292233418090550241112738038880961963002464432975173308155853068617759980519424;
G2[94]<=640'd49997454204035779834496115088932538632764736891183827872024964271329438779096482752984119117636807777786217516217630029501530684676326437142954723390523660855472555124850688;
G2[95]<=640'd3760195009895792369388577389876822495150290405882031777934166332371732531090779749302410945044291714016589080734049560831216806894570119362137954798777160266964039853431324672;
G2[96]<=640'd17822033662586700953931631832701665578404404988930348572694676946112503370956413240471977634543041667202039169121082236217164349539116844093060716613848257572809475435769461648773031581974528;
G2[97]<=640'd15458150092069033378781407563719375238721330678053515211094072698571338300219469211334730506054324381815267648395167981754784951490535947789932385529998384457249697703133184;
G2[98]<=640'd2983422967769323442104811659799485655846368233312270958160160029610064861591740290556516934534700359856712409323113940163642032971396578632067333513132683118838421462276112384;
G2[99]<=640'd2982456833388569127518637821826752658824222788060168983563809975263313504319276608368017246395795267836132472762334198327039345558161146422172192859503419019650430128168632320;
G2[100]<=640'd1716820794600417019630910077546532948365564058940531619600691004388970405032810160801242218664461371307896556264049603526627403280343632646372356394028892989086228215612047360;
G2[101]<=640'd1949659180362206834898805028975186555340025199366023223816694629877813906339552064579718013268824945105811201780927479688958494860846109714387131506322030137121548019051790336;
G2[102]<=640'd1708125585173628188355345535791938061577164626491470177608270010504829207289446931114766564023465200522564464905885127461828935535225738697653989388515836945575594621990338560;
G2[103]<=640'd66972435273889087113570448269851340320188923711714521147534983355250524005062649835943873727673649290719359426750521572825430521703088107747431087981390628162831004153298288640;
G2[104]<=640'd6113883859214407529708592068345168713906710024883376950649697701138899716336432840951039256040713979189466115269660055393762789883605403731086073064591233322029547537647483748352;
G2[105]<=640'd55278344729238863362522313447891146353608522263441234911342536224643442814698183734533805575595119089441683749874707160442893903067593076143372876827438458778189439973954945024;
G2[106]<=640'd1115784248728444521156527692438460746877888193428984589286963242486274495038087242962755277389105216514341250803245998841864195539454724728564864823091873243970886438786294611968;
G2[107]<=640'd1107993824149232105490914949945328227413988651574598779257595633350360888638002163145938984626592021438088403485608740883788280164693284258567202898824253225638073948139004362752;
G2[108]<=640'd8231107454305881177804215207635221834457544526285975521589463048074718508685201069625780697747842835070129946368404150990151884071079420901191118054355636395032424291595897012224;
G2[109]<=640'd94926567446634425349924276172907871125168411783761013577702658288670840656535575269547307199381236508063270883637561369842858770966882853645954326738161406603226585831886028800;
G2[110]<=640'd531141253618847851338256631045358074412680547139368362996015603474483712826656612551131036318294591530710057685557622279214344594250714992020405142807405470819411546088111148026036224;
G2[111]<=640'd199180261374699523116306879904646706450407420731960347404752637390544866324009978914739175018229136602291253337925379642329153004941773021251533366130837840949244732601856854608314368;
G2[112]<=640'd142344982581410786515635656078591973765004672793227407312812743299699497222187378841611519340111576221076101172495101909872516311376639457645914002035331760421889046706175578901877620736;
G2[113]<=640'd1062276492166196414297262169014100302896631427394344740989189302979346309842715187222172281202960085141327656348319595772418436280962487103840606100097792419825319918964632310614327296;
G2[114]<=640'd52068122371380159539726848127070320867488133718713179970069423264655597773849773560021777367704848395619694990729002508051915909906261213891564544762769096091146340822704519405100859392;
G2[115]<=640'd52051527348298676600639804401898186836363289091806805353241633288088211905616767773287175526842132628274857756726427096830947312121622245180812267977922081876236159988294735723279417344;
G2[116]<=640'd3186832009158035789959198028243420797986188254608644318354226316786409932059068943765091803345931679597895926593468027659040013400976723800067123469183780347130042996358926392520343552;
G2[117]<=640'd143606438860094702043542097393897009500138300741036826237401242233719752644337651069731340144624972604038364424621436993323987989450146311345431268085819366240478854479858312601726353408;
G2[118]<=640'd17822270483743299510144940149594406843117770338332589359756563345159902327273760402285869357759310217693599897107084208482001560234786414214577122813358155020350628663563955304828695440523264;
G2[119]<=640'd1086442768358958398104897362550347881588582283846235507425989657313292392625226840946156296078830778300941618738928203539148906070494464255221817964922625926271639623222463360245044346880;
G2[120]<=640'd441842496584493868454225131577039989326280342567882099176608758698359373924967145629159512816185591837571046851222975644376030255345439094215883666042863135036348216457153214613624455168;
G2[121]<=640'd2299077694989447625140676598344756009637433705871696482255329380967590185055028836863736967477734325543583613412512158106335822594727414124978989726378502421412166295472631779728657334575038464;
G2[122]<=640'd8911560687557958464906582378165453056880906845411684087060005496337922493140898760799473633873840849305492037700051009018823164914749978636326762991017506399377977250765018425330564427939840;
G2[123]<=640'd8914552052585518409764943212759026362195075291034935367055688841660776584602873570169065886929512651598469000411451903365519345350009807939567192400245336677924786701720429868049359867740160;
G2[124]<=640'd1015923496483355915375329977482294045889407100684799993946723517125727767807466564272044667078294152950378126134044068435286878667347576677050340116727722840951034117861228754115297897502212096;
G2[125]<=640'd3439774565124849740289073638868362480303650015175339184029693714358711626480457398146825433904779196544700436519199804510474076790080802105624179060302953045092475227187363384552686902140993536;
G2[126]<=640'd2281466110963518803489591654035532640133423061542417578711507442477316392723844198869264114118028192063941071489689669498779930729720555340989868882568343160915094079488676882878838000903520256;
G2[127]<=640'd250620410755596373965470670993364959670507322742309486815510394339361376966901393043042232124673340811689544928020446366170736289403697312397303868798914831859254630560259258330529844504297472;
G2[128]<=640'd3557304575163923343649820784800922232969898657221184806266521646271310849818935404004244267580709430320554896403769051439079590381411339480943794095433535063969344845793001278532722114684780544;
G2[129]<=640'd516837106340795495212065920679429701448915921507100304939381277702539206644062961682799431773349079865932353751734443054927689734897993749885293434415955041437146505404991592466777534808195072;
G2[130]<=640'd1140583911884045743855509953722579615335550063454305128348219521505852624126230046680435212251336561651546448573675562579757713745712983566405616663624301643761795298009843742711265916977414144;
G2[131]<=640'd4562440617599763356378312611157830168118991930958553819756926959569392855088652890242360887377814756738470535661279343672711350891404602345083294534376430038680369364801498608180205224856649728;
G2[132]<=640'd4562440617620137113118001490403104346475118137479064392416582675173571182076291072033304545850093687363023355982784204653557078878221603183591291592185165780578572721387690765414161651746209792;
G2[133]<=640'd4562440617620145280957179738207237160510372290307868112230109192742934935205888061248598936726543522351508285875794357947171403052829062000719190605844830466114796768872578851491300220237512704;
G2[134]<=640'd4562440617619642800556260555466167298620628438762237698247878347831567918647017849794763444036843413239098744224090844945539438923323761508752719368646581647448608130306665967962747375643000832;
G2[135]<=640'd4562440617619936082967684151037819970026033368243003742745432591669741760776697462884194140842271136730816179681232557027039394755256255239969811436753622349736294950198666986502637218684731392;
G2[136]<=640'd4562440617621603588491702245376128422990788165912575733943946283134529589280371849352080009905762890799550435472488965367340592204308390176425981362628552907828159101064850994412626361505021952;
G2[137]<=640'd4562440617622089859847430486738454095787314473859960005185100596871621263711407241231700332298166672362113687320637311525115388201941838865316371064670061401999524054734656067666402672451256320;
G2[138]<=640'd4562440617622097932711734568870445830589600555144242751873800304891392543136470446860893679199884946798666797874715171093905111415285907848627332697267725829962466880458408980380702724388290560;
G2[139]<=640'd4562440617622195218641171605700291324893228507248559930579098168758396217485541951230997165430565814565938221255456200984640248482401275934089963532128885595602522525346474699658648326747717632;
G2[140]<=640'd4562440617622162800550789722942802946706793420052067645843000295694551253247492744184693358630758377569255749361674694742077732224337045914604987235099642814196625065352281483773752958187995136;
G2[141]<=640'd4562440617622195218641171605700291324893228507248559930579191985525031752970936691111334123518607971722800001983135488329983136777339235141926919134196641526774577035523109835158099203631087616;
G2[142]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912792279541091267306519835335022478912340687388711503731613162641292498527455245442245473957317363405684736;
G2[143]<=640'd4562440617622179009595980664321547135800010963650313788211097816719776175366928563895093430879447855678758174094962258344879797673013749498303372753445890314778473435487558968802655600321232896;
G2[144]<=640'd4562440617622179009595980664321547135800010963650313788211097818107464865051418422814954045501840822486545284573581393867214548713046386461568149587125102318281866268384449142968339696501915648;
G2[145]<=640'd4562440617622179009595980664321547135800010963650313788211097798698777006205714405766054756500254898431485756942865367673857484410697231822188787941928850256579090035718570279049323941764005888;
G2[146]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252660640352312460215091290616145620974733132092669952;
G2[147]<=640'd4562440617622191166379873870355605277619924121348998394987168843644490015199566360477776665899259681314727322167545297742440060872948502065487939049513694642789085185248870134131804587436277760;
G2[148]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998156880339854697090654770459060304079552043282434359296;
G2[149]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998156880341594157938399094431607799297643073341969399808;
G2[150]<=640'd4562440617622179009595980664321547135800010963650313788211097820880134559172233282393368229644924525922982359949397969037694129327667694052644397264281494710437770383916433589981256474939097088;
G2[151]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437409582810952780251663771748546042003355591569319997210624;
G2[152]<=640'd4132344820874302116831888191731547817920948449816611003729138585463607160864655899966314548511390689698537577114925406900301440700684261955608711766370139245744544424569687991237813745706074112;
G2[153]<=640'd2256715012525040892763175898976418818370260678257320354787860338517312584999205063710172561315264162372478920714472185735640215134304914463068562730812808485698535149224830150111282931081150464;
G2[154]<=640'd2227719399163840265496268428673468205931020723526042504276900962240074912465904066830904484442801925006637176910495713710418934532552398747640824793779033044263232510775323932438166147344367616;
G2[155]<=640'd4125765984229323827208573508520801009106595575551224234708861935188654996824210392687883970543015135967736335959086794397842408023914081875754495149514922923843583886915928114293827445704359936;
G2[156]<=640'd4050022341163330351899100933035542266408172836661355563986355809403217811431097584513469402386379087338598719491556418495223552574438122455861628701854460954612993907197229465050710144966459392;
G2[157]<=640'd4107769907269250928395298621584039121319401484664474383080956076860701938886687253959561390285283478945988085334406356078165130939922941720379857102148536418153070330486144206745607524598153216;
G2[158]<=640'd1797275515820974774174987300057509734768439890628414401782092091507364496909289260612986696307241557863971645048345268887514502082474146253929254238278358882243223632104092849390913234290081792;
G2[159]<=640'd4117951423175777754980331375554194034438660059337169933649561593523284335274985796645024408909551805729693340703509938567078534560220194002403557889184502119272888210944603051408521003823792128;
G2[160]<=640'd4331293680237943790985225032236964230815381616886725170843994321879267389085153800961848732405466241986251610220224812750318004269633392256351975562305901766450843047360907516454186371004760064;
G2[161]<=640'd2139200978058210326557127785907992208093398735308046483715465815178930468666951865052377650228709521202753545061005137481083324102235888724113683813783055424344366002841947872380159035824930816;
G2[162]<=640'd1003046332068308197409790531673515852730516491309254521401518632709086362168666883573159473072129937678772167211939852731416830453129514436701011661067183081226298551987022550369339749768888320;
G2[163]<=640'd2600116579483230783319532534421139522372993923472426097440376894787477539350412076502372652305620589708255386766669475677160121800182377682518527780992701548238533939677526851417977842678366208;
G2[164]<=640'd2307724927477027023988893600997744425788419971369627089669400472043208524884745657751324127811329874512397212372084208880059701738621120111548188875238355549252829841988744458868622078517444608;
G2[165]<=640'd2717788204708766818592046779824677351964779751966543737738803045730677671974451787475014987003586071070934590977236421346808561366798254897869344131632644927790297793418952297065775333025775616;
G2[166]<=640'd506811770763115029119615895985002344318058111033622006498432640314010550893746972181371206553940847785431876425686303390285146842178532393246090827649771989756979408835350930886731916868845568;
G2[167]<=640'd2802524553533918109063291971340872170011717609926898275299252233768418054933803222206971266178836669495155044060366318563007509629269054393529360093768254955292075097094321325585875484117303296;
G2[168]<=640'd1774414112867683939757274877820534058212512499074646202116272573697350931601963530291064560101713722025884235116198695241923728601346686792653882013829901941882457712960383042388704637625565184;
G2[169]<=640'd2210071544768509860346770863811648355771041341976688867611755335599183897977110482864151408829147261296198385022438866752406348706900762726926106728169473977930920315833456075942156134296584192;
G2[170]<=640'd1643160231083168434596302070214703117873423174534268184130611951115023082882215793765869624140609173162760723701366680151881963367356346736368726049409470643427603318481204106013248174048673792;
G2[171]<=640'd2440557824981017110404230533516664884112906080112186595587976864405950561172284267892832796815783902777528300478921003709436152137188433925212094010996722252001118884534052024532668514731819008;
G2[172]<=640'd2453879860100673889026786223040587624957835197565259457910744916736764394069104949264597756769783382921057283883876300639279101153621388288885722830045077596883114056284221479141192142868709376;
G2[173]<=640'd231834271368466517577388719432872494519393042115438361258333384732135170932863420110082951191260741578710259403267618467397088635688788199670858414053229940202025851818203722303534021708611584;
G2[174]<=640'd2237090780907894066654402906061723348626092600342299609789023711486007141625145285862253096529916247321333473948808090481013593993146876855096090617823306987491371193959158093106215203509370880;
G2[175]<=640'd1811025195516055399233454108266049354215666228797010951501120028216247943232208957642915457002248215795637319161717230969747316978165932051358659806756919055322312354793357527892471270837583872;
G2[176]<=640'd709417032937634566720371634642017541483115753986156364456989631754122549555777193729439996013155114059744229266812716569011304188675783563892106649499247262171125163035075849121662018896527360;
G2[177]<=640'd4131365793316512653125217826084738458692718788552773547239455012240745797373291708114563577297232650172902446845193435517810108487969810030276248919524367145933907018685161463920151656388362240;
G2[178]<=640'd4134711741717853281986422016692735603400859509418567262191427374437033740018017277126854284838551353804750311987809390830786702931717181933889159238800954112027834621856834285223576733568991232;
G2[179]<=640'd4562440481646719541979913351718937674773124266234045441863763031428793958694193985198948043036856232363644718917923044500517749823268247225844768966375505025438981592797801434058724732061089792;
G2[180]<=640'd2281220308806948095235687220145506265864364220713775810323459659910847936748851801856597032405846002802005754165579499537450546515538530346698944673776967773504279628771862570294141177414287360;
G2[181]<=640'd2263398274876717640475385293376011086213828207205583442028634725437045815687026077729644902905757637416453950561730340755597583526292312188638213898189973160375001919569155968812634205218410496;
G2[182]<=640'd2281220308806948157068287587066011611402069799319535944744236710936550914994038142356557356052133042381489736152253185697685527818337743539317384403862669509134710260300344459401698539556831232;
G2[183]<=640'd855457326860943995605036997390587002191466059201238443864791806920651360049085189189161207921159286508860704550791641454767232816724332712225196397343012029456356251940944135562094948565123072;
G2[184]<=640'd1140610154403474046999517605687866004614420274826703981285321394659233294260780702653290347024694019049228200268422103217498553139840791206381475303158655814716271861729984721375480098953691136;
G2[185]<=640'd4562440617621157839872616558197222509213164461019063983032264643949446830830880647879289302672924423819468758258957175651067291574370373165637888682225961031759968971257739871373153516805685248;
G2[186]<=640'd4562440617621676529195061481580479007271676295083636407730113981338563070574879341089102069901094880747177729507461543521171559140002770371686861196725382702199700357351943943578245947210072064;
G2[187]<=640'd4562440617621676529195061481580492431383500680490934054837126585002999440955608771322830140774389318076872863623871469186548872614385028474623787237543274294247233803248920169945150389475082240;
G2[188]<=640'd4562440617621935873933574693732475519806566759370948423570255705974729393435090724874088744033279747461796631877139545367383970707299233631698325664542819187463049270516494187197333202429542400;
G2[189]<=640'd4562440617621944041803669241720724570542824511988314400057778764201751278638458563012460940886177453359591623953866912724927548967051965986325914330854563009031379525896884107431616273423794176;
G2[190]<=640'd4562440617622130596323914363960391720930610303823460173668293708009272858764935392834685107443957675837211090398518829034548228725511806888808753469856583254988653618611381504702553473975058432;
G2[191]<=640'd4562440617622174981310273721775935754789341833213717434236125404057492264323711551249222030657299420735387769477376622323474632262454154240476801138677007017426708909828708751629777000242085888;
G2[192]<=640'd4562440617622182805615253398483905112276146870273243828932117172149132426940395788752283764117992523563880387998537839368622664008553551871316874640095906110768760730480811646283302871385511936;
G2[193]<=640'd4562440617622194789948024177395823351904679939889531683015844306257418826397518732405121566089038679423916320360307820859126596447109093155429367048541287530825231924483792072586969791728713728;
G2[194]<=640'd4562440617622195202498998372057203634099214706408914219457794806182845515558736620168677181273551312567001205397329825133091457419785737790264802340661900775604045940658501644746965530607353856;
G2[195]<=640'd4562440617622195218637790135367651333678382636433749881363343741788073512895817107953779282379283381375864074390332059015925799640620753229963449139587530168005027624737282255575898473541664768;
G2[196]<=640'd4562440617622195216658663856397837424230446600622744306701574651059995198082678821960540075656991556322253634842674062307380668683614203111322950282151704488712843645962021254249067339057201152;
G2[197]<=640'd4562440617622195218640205471319649525198803917485381701469952329986853756662261838986623082962202993123477046639350221934028485140205459712664065345255289125361622802948566744753990729237266432;
G2[198]<=640'd4562440617622195218640628155140247538669856248398190075942210407234643161672722636519055875706200725375784972993783984263922866288280450114175360815759392055316395916295475942166233576359591936;
G2[199]<=640'd4562440617622195218640206887016473440411796000961706555542776546328286749969490281118469453046576123297158649006928255904468402778885135681862188795876439605011665917435134579941537009834655744;
G2[200]<=640'd4562440617622195218640386636259403237070004483236292316048774454520700236583045508244564080205921927902030883745497487981643054270148270600929710490443901044293498447544020123989542361827901440;
G2[201]<=640'd4562440617622195218641057443396079198286262004248221672302103085233322564355405200911726321802613200574108755343690193535427881104885347598041700421478625741616052639616167504751935054485127168;
G2[202]<=640'd4562440617622195218641077256915004286558674276554906178090648887846713959395021728792603978876533948845034072177194073402099546154483886212364555966463808821105473780463046917739773791744032768;
G2[203]<=640'd4562440617622195218641168053386667407889743163606142251738436784914176905507608786492740672262485602258716100181554702212851350342920816034170098191705395141912351251261959721699380234779885568;
G2[204]<=640'd4562440617622195218641145660413965565800107106092747743521901170051942801650748874896505956952810740999742609191015886761660610430681467668584998195133551576447676194304224628420108517935939584;
G2[205]<=640'd4562440617622195218641144953904628064717245082818540827229138302639417854197484766015141973473817417754118360616235044732731736703824894396033681603645838217979328843839097527591617410612854784;
G2[206]<=640'd4562127305693888521530859801892304502279590308223530167172080244195480407553558188098147892227235168205777659784802424334697763958383108718084620516800979523572131231619574401647395733134901376;
G2[207]<=640'd4562172628761091561900925181833146037532497596226823438775464781152413266805559664401101008207666196320928292269466518717425219320449113677882925539126190093467072366649519845370270891047387136;
G2[208]<=640'd4561981306503170626435176972678649399021765736120620305194463398858334495460329632647145975873094411462301033093680773206944340232714115255724852823278735244413065906691087721049561264413474816;
G2[209]<=640'd4561985385622726190908703405354763416713456847613248795029888003844997784410350451367238599974874731787488458976938796467939842677991323828861327119017487988822139499369992865631752476405268480;
G2[210]<=640'd4562431915457563854457142464823995847179565348381338068056807389891342065335504638318630226539419101200195343413074813551849146326328283911648482980207128314481977630520088326083734766618673152;
G2[211]<=640'd4553512196461164914860849890376218197890227537333382726896407016619919879446002059312134949331538391909212250283889318169524263627047460239035353521583678458422674513366801498022075196518694912;
G2[212]<=640'd4553451281307033087310031542628667632521465580466282610869715906516689543940417891629799307820852886498841739799990729619177484334011520005160494400063750804336494900456618035275840489814753280;
G2[213]<=640'd4562334016102484926174682634158555963197889284905814684926180282282351232037607971503741692151026633908857549986410566722637304414641140272814959937537453331604866262152192331446489862501302272;
G2[214]<=640'd4562352508202842832759347399076719021461598223862623948988567601319772097975443638192247097980450561775062633096132216176873187127854753890388888125126030700327956504715278674378376824615862272;
G2[215]<=640'd4562407984503916556594293318137433008251016637557230376755396818602030054370991063790567529726498155590564173784886861257655065640207399875771170088813112407594469726365505030485830993767825408;
G2[216]<=640'd4562423213292446599187877347483595814692001952670749036249830142165572376255922450238968572100294956813485394868244992381304159094481861446003142888215354186976298271012984246700432287392333984;
G2[217]<=640'd3778262434303506105772405707230482131841717210531220042854995453293788812346824256589961233540260837540254478414425610711068260189823350624262253433866554192405894359143332368139733020693495808;
G2[218]<=640'd2290026899663899240426713328676484209567445731472537681988848057341862040466824959841541381677266347288895256978073778868076988902006942701734648653951386694766964273709987424199865428667007040;
G2[219]<=640'd2645458121790213299787859851585833070401792088679240761626561258536595222441572258994723455724592211741088629181738798289789526792188088776591921182360070361911269022679059626490635224416320;
G2[220]<=640'd1932268761508629172347675945465993672149463664853217499328617625725759448658739624419429118430836570394435353997528909193007247029759673821230266611257295788163391758041104;
G2[221]<=640'd241533595188578646543459493183249209018682958106652187416077203215719806409051140420748950571227625594886594016189517903441651975109819950498422400558334493613662923915280;
G2[222]<=640'd60383398797144661635864873295812302254670739526663046854019300803929706630181609407851707922557469225128729411869276182656732663554619667143524796430626352627271918289024;
G2[223]<=640'd3112136676664518681309125722921197385187894197597544825868855120337540764942318608735215499614208222611005807776476837065334282913046083580923391754761728459442126580206681376292937;
G2[224]<=640'd14977157756429892927793568780807952770067586169796671774456591064614646344944263783468807654258641775957884846730832112918752250056699777192282284965613135448426182404043575555830401;
G2[225]<=640'd32612598924174068775349129459260005950543021718650164085374365691203408759344854949561242832786568573106113609645052076034739221801769442538875024719251369227967045037153115244368385;
G2[226]<=640'd33163706460666064423362288101788068436785988208008001788225126404859823193067096402916629158020217542421807946482163106631564012054200048048912022195272774493969598573191338709004448;
G2[227]<=640'd66367935534309476656671109603288159920563917529614953555747415182401790750864486668171119725969435869470648473203926044186230359882207754110114549743362495474916032984433401833208976;
G2[228]<=640'd66376040056904945957672256295163050958050216669627483266186720850070761943469590409260034445292147547916872983791030225361146732480782859542365361774689088673359623036327500087307408;
G2[229]<=640'd132768289159000833293680984188514338276848703007892960292548961807725678518030592008180959746322559359890622249938224038599180146000572234933000119197599649876704556581551783079602896;
G2[230]<=640'd3186811747855411650758785051079693927895637254075592563200472773343915610056062974840499385591863992876208759882612657914191886249836437128490522054008791981168368581483668513969465920;
G2[231]<=640'd1062271933372236462034490366260682722517784758465840681035482194227233539024166529385210740594933009594154334410766696599603518879959825926506463649520448030407153211715602701450061376;
G2[232]<=640'd1593412965388841399755610366291037600844349539093706661450500941986444326451546796145456102896438661375850778618904921235277303209772914165386278773682694977023200506517807825693509208;
G2[233]<=640'd2124550958213337573491233089532896931944014714133728410583934674289988741677034404058479459759059411503956757307052854975157641182978227414523109780425293474089253477972397279055726156;
G2[234]<=640'd2024947388568733622375310848414884713943225818964098591249625472188380534275144987955397404314533602210089737391644895843154475905890283349872933844210845376958562348883386569542618148;
G2[235]<=640'd3992135544668395086483634413474507048962287517633263052275550337252344157844662711643442409983967013597854335572472035680710833792435999459580839607007124337516422633794307657168718759326745894;
G2[236]<=640'd4419864349902211662365661817828022559608855082899204751839031172712319727976156027064316411314914948297250328268223019682305363159974679878721239013872384460124184911867538522485102877199246338;
G2[237]<=640'd2219817867703910556813876456109094180437867810106676781185739828034114554436340693261750714043676104164492276528703784832000153757969175382807735237753561313442002814067863866109741529458346240;
G2[238]<=640'd4500898907632108846614063951197598717902617221014090903927879307561737300538873075604975262441263830182991102059902169686135019226682472034486714848082332967152469682417163356943459499120870152;
G2[239]<=640'd4545175522511821734885535334445261311350609771306604376299471469286716250637847726020716732892232666725768631091501567130164337684122601937906560344821766259636478977382258992544145085009676616;
G2[240]<=640'd17822033662586700072817076584766762987962362787994509390621186724926618363666206956162021507171146852321298910141351184443895842815411641113330749777785978508271877159792436345946212504230190;
G2[241]<=640'd29243141876009673659063143893143434613747892028517535834172997495452570282724573074289213676364644861350650254797836450299337500538855585857211839830020;
G2[242]<=640'd153440184745131650156868267038793710260155095908268662007029282879506271706469119760153285577778289860527177570070636701178195671122700697043199213572;
G2[243]<=640'd102293456496754433437912178025862473506770063938845774671352855253004181137646079840102190385184600668552486799777354396367116647761224185238603203846;
G2[244]<=640'd9143154243142245628345881385804288506464786863760416;
G2[245]<=640'd5233830162798486416158582881910927378;
G2[246]<=640'd4568889111050977898048726205009899835;
G2[247]<=640'd4569204756048210344620200811022457225;
G2[248]<=640'd58064141215313010447381988748107583537;
G2[249]<=640'd27155685870231588408346304098211647504;
G2[250]<=640'd445245460324152851054990970187215466226873065374425001088622824982584004690;
G2[251]<=640'd448779154453709619714157565188701303437302628170085557501025652974469259393;
G2[252]<=640'd901092003036976008087481725378888443436462377247879497875909491497079320808;
G2[253]<=640'd1807484547268287169163713343260005642178584519766258678798998711559010300140;
G2[254]<=640'd22895419815311617052303699948472142832139702861650518898866955748197841366923067249254426805540895855436888338686265029755480615542692196;
G2[255]<=640'd23077129496385518774943339611744713954744457676828216203808734162978760124828242412722614365933436042498820616905102546776192371962037392;
G2[256]<=640'd23167984336922469636269316006849186293407800070545475455776777048633330476392252023363898450173131911401889117763882325377943328340362368;
G2[257]<=640'd23236125467325182782258526748120701839120657617426447955831049512785276051673226840313810606753414898839185187056658680952940708371637250;
G2[258]<=640'd46142902137767380065496887304791685659238411560833261716464382462467165084689821804880979356768740550606615240064768316684958416622555200;
G2[259]<=640'd54103525322466562515462086292188350117699351701388316223469790892453627240558929462272852536800804546454182997865883184891364295224856176416851512747294400590194077686202512;
G2[260]<=640'd61723155457956415220274357196513720302547219967566568820946051829750034916239124804755634887100015776451813403195176406728154362843305830304618357867694595921356180360512288;
G2[261]<=640'd30915474629859394004543151965315236122947302709170648555409007509240472031640038089804319714829075554768790768909058465411852030444337935942458883039250692381052805485838936;
G2[262]<=640'd1932239277434214780044219442783777340708970002428699831946073019757539473149251473846039118997674317614417051827442587957953365337466385257218790070928364111244171068646404;
G2[263]<=640'd120737615846881945639764057123609930939379089975253816547659748353278469829351837204874270236688448951626019779145394620154553507127382418661828367469083620796340118962876;
G2[264]<=640'd235685721683183012331141657098874671513008558759175149554300194468636144523282287392041576183926271613791237993184632790004303101354479062879156012977992487213420668821;
G2[265]<=640'd106707036944493345812662868644650354626067981909427276715744110776408924732529400070970502959688509662155339720769019779856461491251474172200566219564303218940405623809;
G2[266]<=640'd1669996800534434497298491456961972307442321941469815657399664230060734886256507439336635236990616144582227146568690898451978514024478049314698731128557996867503226240;
G2[267]<=640'd4019843207353463771313985362844050763459800246888445458315586782705744594914299078377691788761823152493760708895431509560709958753199653971049440710363992567926099113255210969346489;
G2[268]<=640'd796690780179959721397678842694631304588936441122906005790475440643208793129243325213130718004974811755611612309372981906684020703101804385999608563465742386052653614809254790738158209;
G2[269]<=640'd1062275981676247891745829643810064175892716773949708457431636957808693167426344228115820824086167800529670042784117999004181953542464993376761773077695923267208328566022651349481572392;
G2[270]<=640'd1062275985409391492789478531805275875178868265165153010987501901804263228776124995191778910648955229162943529228212512053361885512637065244737960784157972880926190456649348369007294806;
G2[271]<=640'd12448546705193777304405751711812726493937843442615046591165411615683920510093356175818329801415716171401862464323141634256903799247341022960790371867795635491817582810962263054746852;
G2[272]<=640'd365157370061527380349091892004822181289095268437334097843236385790105140524148714854627587316273636544472942541367312005765989785807733190315067401662529129864782320383382542260245568;
G2[273]<=640'd33196124551047943668099262909529289208099569857939323294444223147003928629623848300008043332478157053677922523156408206938077259814665724040480324363504201509160619969014017858055220;
G2[274]<=640'd66392249102095887336198525819058578416199139715878912765179081892234376787009374336051616562915550185747061412352555417521703859689143285639832182534841944512831600964715461654939160;
G2[275]<=640'd1062275985633534197379176413104937254659186235454063763565381164541463189816580734203699364366900944485258475754415531168881587982239926159579300266505695475124746554901041021169780390;
G2[276]<=640'd2124551971267068394758352826209874509318372470908127648781645158633678343636083797685196217007478571084469187113622661804273055936304063198037408850985564419387030451292486389681886912;
G2[277]<=640'd407913978483277131793603742632295905789127514414360514133943199964027581869031072687887635628731087637279743940034858888156840476942334401173118993944052089505054843649872231319237626066;
G2[278]<=640'd4351082437154956072465106588077822995084026820419845493512766749030975210494415218446118578761656794644944932926905723697900903715858995601119728256331634659569315533120121753557052590573;
G2[279]<=640'd17404329748619824289860426352311291980336107281679382014638748990547478526184095995641377872118045112139367920206701196875290525718152202374784317357446434578281929307805274507856884946988;
G2[280]<=640'd570305077202774402330146450712536415611653563406069991322396536616369990967646252236793886220439962575263817352719551708297507238830282744067315434536344710593242505688184457320248839397197202;
G2[281]<=640'd4562440617622195218641171605700291324893228507248559930579189989871650903336926575444560652131866878561807360788663165764702414427850622163724022990549856226375286183202653099243416961331261552;
G2[282]<=640'd4562440617622195218641171605700291324893228507248559930579181316660294630881746547159910646277094979502412425696607790469492969228119566746438782703062316733443820157961365366129247453112776468;
G2[283]<=640'd4562440617622195218641171605700291324893228507248559930579181316487002774999195618436259759768152248037635108485619254521337995439705735008587181263044332767383251502983791130247814405796625182;
G2[284]<=640'd4562440617622195218641171605700291324893228507248559930579189845089012998713790485095552019011916969919495976589163076955411735673538171309614951143603113278232392845405196161265880544319777101;
G2[285]<=640'd4562440617622195218641171605700291324893228507248559930579191264695896388570998589243614300270773129375278569007249564240957010359647767789933947611239184070997406050943697126455439014402104840;
G2[286]<=640'd4562440617622195218641171605700291324893228507248559930579192507458440850284983930905946899153571829025808947611535116434351533969442075792693674559405889754030333517397855321971241471347560583;
G2[287]<=640'd4562440617622195218641171605700291324893228507248559930579192508194931237785825377981463166816578437751112545758236394214010172570200860678562980679451463393720745764268046169144176311826180929;
G2[288]<=640'd4562440617622195218641171605700291324893228507248559930579191048384337283176801809946395215483008578466992360390809566956510978972082301016672450133093122320026239236252904507743510506451007631;
G2[289]<=640'd4562440617622195218641171605700291324893228507248559930579192440264523731825861318310315655311027703558404199050730302537260447511978819440735216197487341901763970063933046356308035561496628042;
G2[290]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661315405642889965560387311358996625454767730294924;
G2[291]<=640'd4562440617622195218641171605700291324893228507248559930579123312063709911669782309287876599948133626309240929191878152140356563773532609582701583556352758671418035478931323393905006752902149986;
G2[292]<=640'd4562440617622195218641171605700291324893228507248559930579169804189140929493347720136916311175672848486120830884210610741964309743621894313148717846882635111531841556350311148723822139758167322;
G2[293]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661318353399434544605999182138683236876501783708594;
G2[294]<=640'd4562440617622195218641171605700291324893228507248559930579191098292391777351469282357850530058515240322859717155507920025143430035265841517933664851916735207646892488407497630615469247189514033;
G2[295]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661317603384752938111135459315721846269534434001824;
G2[296]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167198590472919635824639027965513005544439493994057449550374380674886765756545990292397830065086183228098042605254211585668;
G2[297]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167127982077815696917890623925653548188500791101284775469945417333106357423130185685614820034584876731274572720981105741652;
G2[298]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375387781438778223050394822354451649030004477163395365008842418;
G2[299]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375246546649732021976070331643319091348739946221361461535532664;
G2[300]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721351142475985660097644746049366434768030806222937528836963538716;
G2[301]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167127982077815696917890623925653548188500791101284775469945366119802573509672226839203115383675026344365243315903388730880;
G2[302]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167201112201316205071308613824079414735723019097370759338960718209909272165888138777038076586990640704014701903526425913366;
G2[303]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167187242396926531224335643657469475925740772641092888171550776382159873446981654552245315173412202707255481438071501968647;
G2[304]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166925594829748474565171666033775491581198215832250215072633589279214035103223232981773032643333774443040061598516880368901;
G2[305]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166562464708127355605043624403813150841326528988375403849056718604729413445209230024181131482196228145487178938184962454811;
G2[306]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275162039744830082865505521589677637680339880396753970647483764204347767223250517040531257977290895533305963363058380935564292;
G2[307]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275136201544405057391318485624943380701382064480218331207266849140896187101329886438487786128122780382224643562530205844155451;
G2[308]<=640'd4562440617622195218641171605700291324893228507248559930579192517899269589509223461666233250460106833149041093565485336529135180534088454698961329756742589652554400039279335434450813064336955636;
G2[309]<=640'd4562440617622195218641171605700291324893228507248559930579192517899233024255191434185472430277808761698526061984619639671512383355709900820722129198386680617230531508692717692098804872178572456;
G2[310]<=640'd4562440617622195218641171605700291324893228507248559930579192517899190563028848297649058540639130753973395137475332913578632849571796223775499973433501560118351621741587726811498164783929898113;
G2[311]<=640'd4562440617622195218641171605700291324893228507248559930579192517899248726097768797249400266703272906569643343683374971270010396949459340143896717475916399735193191510310692175189323644922011777;
G2[312]<=640'd4562440617622195218641171605700291324893228507248559930579192517899264592826079085496335187261593326540851615463606348740136074421144675755211088435167268454038165686021905106900155381506378340;
G2[313]<=640'd4562440617622195218641171605700291324893228507248559930579192517899269889091187440536893677491691429156152619745625453363772339772875251689394216560408525355479887240235589887826896275313009176;
G2[314]<=640'd4562440617622195218641171605700291324893228507248559930579192517877613690357597535379234017004937860795362735587483541862782707340654226691641688376111937238702498161780888538371495423750443147;
G2[315]<=640'd4562440617622195218641171605700291324893228507248559927602061103184469348362877623219786818963556496577699272724106162266612221857731238850788449995403349848914603954119990567791934844523384898;
G2[316]<=640'd4562440617622195218641171605700291324892390519252938518260469319134162206995263381384866652186411226513487030368100786767571520783595199193895486466428263261671960759802334049372386167765655878;
G2[317]<=640'd4562440617622194205583576246908354764246475836801576934847604072446548246397102066373909325495920838174841493980085912696938579461180449107948663417191604282325954686545284524645705742314547361;
G2[318]<=640'd3773962424821541352241554580988268890916596298186660645385150054666297192237362287380562766261918990316254320244100708867464887852704836484976346192698161081866230351571;
G2[319]<=640'd33992831540273094316133645219357992149093959534530043084755624867769292041820444557712858821731192346761349485417725188525391788685701057757540726920171459953935709113634592034324925194;
G2[320]<=640'd4562440617622195218641171605700291324893228507248559930579192517888444426216017953470077941179676809439044393016825139063279951283578586102122873931934053397270789285631196794664642839953332728;
G2[321]<=640'd4562440617622195218641171605700291324893228507248559930579192517898936706552656779225526874805336762017279216144384150097712412456753670165607504584670682269115900608993210604446574289264075060;
G2[322]<=640'd4562440617622195218641171605700291324893228507248559930579192517898936706552656779223324901118491044296929109222501895040161489903585629982482525331395364035881381633346454342854093324100581064;
G2[323]<=640'd4562440617622195218641171605700291324893228507248559930579192517898598245896636171940586121713777591923592760803912551445167268815012352546438145230437941133677607290067172768972436824394332304;
G2[324]<=640'd4562440617622195218641171605700291324893228507248559930579192517897921324584594957375259289886392655777975842004690571955890105936034594517289073844031131780053196130182370037447868498198171844;
G2[325]<=640'd4562440617622195218641171605700291324893228507248559930579192517898936706552656779223249431239594806550701219007748000657957879668514582365690294178565167385166551258591756934234358860102502611;
G2[326]<=640'd4562440617622195218641171605700291324893228507248559930579192517899105936880667082864581121041713212206910723480164364677448331074401832975360891949936844125071968857030907033666271943801311361;
G2[327]<=640'd4562440617622195218641171605700291324893228507248559930579192517899272522984802225511517003656143540668554837775012982010147186591672057773838103746050015832816099163067980709210312890616653831;
G2[328]<=640'd288935169755614940720218082440619488819047955675266017010293758646984841736111227741875097862950090563316595211736250078167773064885583799718476683985115898885281793963840602681836833926;
G2[329]<=640'd1062275985633534197379176413104937254659186235454063846398888276400807119721704485478325941110711626502346119866641347696680371736603254706879576438834967345243091739208897067624173718;
G2[330]<=640'd2281220308811097609320582028887720840905262012069698977020705353097435121103913505714137619173598830843504194369645495118362053289182148774635215221154313144127723212191396690106597142663804551;
G2[331]<=640'd17822033662586700072818963565979173758540294633730181363270351598902816459307015948591688724965205767896542253011906878872394874418010565758606190651187244941503488259740291189444451961944116;
G2[332]<=640'd4438104085898055193914408719839379454985707356828242425146843307740460727190173125696751016634280167111914889089523814460052740223501270795421897836167123003989297071811827278816188622727530;
G2[333]<=640'd4526935784935010777089856335941576289253342848393933991178017771437351486555655757674155982493948222780654999846165934962622943015314215726748119303507924117126434254058333099664153540778146389;
G2[334]<=640'd4009974978411748031685536621309501889014810682007088234683630474810860061735129077583730217862559213567302729487897308316998117519727438684676388051341394183390810930862970573924101015800131613;
G2[335]<=640'd2209950122375804073223116415075754431515012279809155448237045131473779477153797927007788159761128084772219137958391528326890032447824413047840312687068734183371065838309634800551793966894708474;
G2[336]<=640'd3341631312000566918101804524118837370871737961086812409358055495872543626689363886387578088114355469463399667972438313296556018390052652117538629251711162095493829452673153345229427341860292616;
G2[337]<=640'd3350472711249379401473374930070602824445387218177015674906381509435905436787216412187731256017673092917724913412614078260779646834045689785703352191530065594025268433443958879676096929935556012;
G2[338]<=640'd4544653324634429655821084078171720532596032635021779475581272289745895602059726977787585415618350908721718935667192704814884611212046659616869326516013841002975534382700706421076666414740808446;
G2[339]<=640'd3203545087601033959042590967209172640860890678921801742317406549154216397373612411865744244870778801039750128895640911053691231882516447366742357538932847296417035807939828163975759216198944924;
G2[340]<=640'd4544613145109933556041107503130045295334148433337873090449235325017116323115255055660090279705715858305469634463032421097296089937460140226036523752553395257559100156045459329947974191794107181;
G2[341]<=640'd926739223837133612807684965469532095396485360547549409427162435993675687985518422220996344949066107588561724437315909718194840309963785044759409079592944307534723295753511866472587926569237075;
G2[342]<=640'd2405861416318319445524047975093652676853145011497375286977919777656971874249904811091498381589674362891325592855219150559773865834212420237122138538738826858186629577538180251244575084749334622;
G2[343]<=640'd320753095102448388994191548100678769471405239793519941498717012942862805566427473152132688874359238482880910019197301638600202582562286443841748971992313977496209023158968330239758376376547617;
G2[344]<=640'd106923499810654556982991281259052216875705241495269111520467363240801183838678419974717905651521787666693028476815047324714230482288524280536113929115739018574674751116263546944167721464109323;
G2[345]<=640'd53461749905322945263344899028466525726771275515231638677034794305178601909428616834406526226646622185629019232651125930509607525713883955568675836560526985161267982513166826986291763328857920;
G2[346]<=640'd17817682580149545117710745858932999751042927802352264219384852759090514665610771844361777536815576591570380045464599131709716478546484130859365039824026613679309931437026414166827157434929013;
G2[347]<=640'd51473305231543130338228345317714960618017875258299769276748414509455670284620180375963776758758554663406964586713466501827109635781907437906826658534094529841560749004716329281889028419235943;
G2[348]<=640'd13575377203923462946574199745179965037749082666076416424368886622242616459559364138118305976487476417935216391747044824799446445070388199326676746781875343909228037734968984773374621179325442;
G2[349]<=640'd53344160202817255560880775185186433171664650481302771864982758820312572417132964749256304363377326204685008194187477356581440255648391514724773378523851503451155827277711944710926722066946850;
G2[350]<=640'd178220333175544805203626064335206696604779301886193077245886154613680871491003766476989589136553014885820361567257136612762450381210705162414148579125865749271866859595244622409792291633891872;
G2[351]<=640'd285152500373975022848926538551316968936342738389519328194972320388339896237450832663178069012765566951020075173385449095012226029560253765547963692610331297170215497478253003612797530339154448;
G2[352]<=640'd196042366836056747492003405153052947380787871835461728965890459496579799919368017327923639608005185096286127671497467974237285272177999427371748920959390530222789271833445204840869736664685743;
G2[353]<=640'd71288134384777803882884757886632499822813010041706164781378212164024672117742286905144537362854707623313413991741698896117846914006325432412173629885455540224271994514302168710547561324484656;
G2[354]<=640'd71288117649781514585844106187617517800263796921509565673990930715451802680457794502143825086043997740855051916391300149467932464297051320834668788235513733713914707055315782742484797132115225;
G2[355]<=640'd71288134650334137778536688176094484384826071969695738895461540436121204616103961196726576178642287949327424524154222594556293133806472684864632838234885072210446835129080811732920530380259503;
G2[356]<=640'd71288134650343507832828433894639371444722270730844737672085686849602481135051550148893066540382098550929974608691887526464835667717477165933027518949186326771215121222542020194028570189766912;
G2[357]<=640'd71288134650343634462129450601031271439482172226160370743868272259962969085719694643079567558844749003700681984848727479605202899771965867700424332924060232070274537453905526979080122985087244;
G2[358]<=640'd71288134650343760106456466128514173635617924100208834612232110057297074357660637015096899929068054374522967195873354282898841578637568589582242111457068418300468349024886723639203746862596480;
G2[359]<=640'd71288134650346800040072987735756659085923724614884292513263224503723818798664438656735801723744026785591941012984728605500171701218494718398243074260848355946191650337518854061572579783621632;
G2[360]<=640'd70739898263265275826032031910573933603864744344658617537903634680552690614727617691070025808177173645497643149515504681574648638792570886038282226981940663202637115107435842477716904644581376;
G2[361]<=640'd49203051486086566391991328603932497583069138609761980239855538211358517902918033485878028787337356323879380335200768593308704264641463947016622785626522255977664906627707448448701791343895552;
G2[362]<=640'd125868638701415956067890080744636801960944134105647601659842395318352488424868673570228915903690130618081554163308655402763063174143251153833995623899254017859422895083391377555540334887436288;
G2[363]<=640'd17822063406314297811774603201706327353379409081647104144739182819041399805490075297726696431606795475304606557356084961064959671882985917889278574824266386131840374426290141333709053678064128;
G2[364]<=640'd124755091301413328321515525019968096085165119446306154386761035646124908391493626972737795753681367518081169609690536540833173726412602162397337023493474828404060715757857071672990238261903360;
G2[365]<=640'd17822048534450498942295839893236545600143013562104110369967597948430926498925566479245571278804332461082574105231588228703712780067056592018727766448896953900124812217982222681333702592561152;
G2[366]<=640'd178220343016120976804899921956775739324483058460035688697597242996874672077145801069610655123136610504775688011137277024872173766899427318319328374461349802282834292525182843866481302884581888;
G2[367]<=640'd427728809794389573518870158146013809658684159540870221312356021438980527723954654403496621553269497260497470625684273923405174240588867793009692979144179134782301149195596422694350259541643264;
G2[368]<=640'd9622094451472575957019249822717465845350076392992350037428194648230466255805677384018541328234006477691016878346920334524878140641488876557711777053702953415420652097992184029253696;
G2[369]<=640'd103585929423359748537080854572169982291584365231923134476007534440003864401481494612333229033840599659658918377680629626589930979938238079998705623859047948803196196578630142408704;
G2[370]<=640'd514383349428130051793196737446001564744469354003454130230747794509707801921081947602326587541059845010849058330744922610603289840519660853673544418566274755382029982655137718272;
G2[371]<=640'd49794558935160931787920385817085068023438388167781593962046500426360586578309373423419158239886993218613989851091603627707611725119121857820316328594857797753444269934893373485088768;
G2[372]<=640'd742866763701872173174660413212881585632423109607096115110387839124566458859896173020005571364198597769229726668253838546404512184314299370525579680013117803380294963029082112;
G2[373]<=640'd7780341708144077593680843819253666659957864612359568380200657379997637573172993988193794353494049999491702697976235923928726881167966657331001623396089470742328581562360430623457280;
G2[374]<=640'd1004960801854316370200773738622911571901931037752646339075668241332055228042990724705409412784879109088981649364423923189609882741600849086684271479787756051394636573550510627356672;
G2[375]<=640'd129419095206893105333296437803033937280627450126556412427207501288122571917556394387150778297976162298231829709700744646200545104091586415870474959515833696448478558262419592839181;
G2[376]<=640'd24816143162442440902867493605441452153074577596816164970691482799486526957641795018460328787353314385216863738041662702145596765689966790270628617803758689691583827018286144421896;
G2[377]<=640'd8108448965594428521114630688168482203276826604479045123339318880932217497449099691414540588727458269570568002263352577412581272208775346064294267573699102909276682265232270163968;
G2[378]<=640'd8104553270237412444928433034496668500393175944223711634483579786591646211230523434120708748582111115239556725382200295768012302063193767417296643430990969150015389288635840856064;
G2[379]<=640'd1828266447512495986757484195403266031661505930683486301783475051955431264433057156326889065069656787100826872443999046240890432671535056636293044507094774410254123767706029129728;
G2[380]<=640'd204665911449959693118923406758316693415412374362975317243030406593927713197415582445408124478057247985182868599972642958910531421846496282865548453542554329006894890667514789888;
G2[381]<=640'd30674768316533263909759637598169020556877941719848415019746973417032971041173242028354012854823035325324676835249652459988189231409812144282038332905056206273629214216290304;
G2[382]<=640'd6183494022548340121575310402936616067116402363348485034370679335801656072762071365073878908928250203561675297770597540978667088435993076150199849698758535865548635152242966528;
G2[383]<=640'd3091631142494742114123005921833631362906024116459792079481279314894919022696614985975681139357795052513439092776113504403679607945388385815241705621797423311554863369772072960;
G2[384]<=640'd231872254627451694824174385091650733176312570627734139960098759434982749951057001501355989227369895117336676011467392697836368387608634395373149404884713013371426573276676096;
G2[385]<=640'd748723953385279641076885622835542364708511806301169172273381535615005804154678710788131531030736379762939894297101869794386683380515662238496565436078429019628866444631998464;
G2[386]<=640'd231932516843507693445908940443394842208721369150576046146872050833085479886291730403808650095168271707888535850029210967617858864842352159490790705660907097608980519538655232;
G2[387]<=640'd54107298392081953563722179072962664087109728586411085689811852203760569032368640105819879413033143613076974728569453044918203648313940296128845380783153966922804609729691648;
G2[388]<=640'd15216618166876376907380126244519951600059365702900759575493214712874440389278311530450212280264381031626381116312168815469869947341863145824817129260072114531827152261742592;
G2[389]<=640'd6747844815584403456136364952116163081812777201340225073939750626732428651737144930641992209788981323021417437415706060407000769847268337833489537250962242466275105991294976;
G2[390]<=640'd2958771799019393062226847806142426237372475210075287451442049744518805608892556682735240377427617893850830596330065391283959277113430426551309984659912103908914689147404288;
G2[391]<=640'd1690970970475639772564631495264411331213454859746898982464529999590888045117794279959946352030246267860595417271094182033237941627768974060573401990780229351462755914219520;
G2[392]<=640'd467985909565985966780833791839081418728900149527493089239661387662908920413560492644433618293899001770717350049819988457452107855884161612223302808062895155123611347451904;
G2[393]<=640'd58496475170833786249945063306340430006380363563121197005947873304584803232075588339684916287927736013091535047824135227245998523887068180491048829989219116777910757752832;
G2[394]<=640'd7429988523867462749466079679148621218002143151264323466577944736894607273180961272256124358587684220816569210236477020903507629832120922680377021812268409061622071427072;
G2[395]<=640'd235671100213351217492844234147001107763484707529366194079596394471879813521616320956606198245569087136300619213260770119732197363648079418379103643289249717611057381376;
G2[396]<=640'd3685165787307366687730439367660571144462103950520914684017033789092750560402928583513070860464296661638077967550077036167738092432122355465397830737093285334495526912;
G2[397]<=640'd884939938991106671122094067516557306135352974678287926842806457126129509095392323331517799737175118920904069855038555812658664728243245767273999349626077502469006426112;
G2[398]<=640'd232187366316547949537474922875920170737807926435216821611283762579450440770312757452550393912888935543860865351780127760184173304196846464020171274701723435674307133440;
G2[399]<=640'd29023392671357127399446976974513894469593819282470986823233494850095033843668164683665114850771148470128175124579533764998714072028013440244894067935760104796440231936;
G2[400]<=640'd14741112824467509648154331502106848963300583324736293259105677887466135140869022462778926390525775756967434762893945802353974023893807088280957849855855029135723200512;
G2[401]<=640'd2994476143382822308087637626941345667970563784377173008533996661239113237678121844090783166370801346829784844802092568654256797036885847127747382933960656525251837952;
G2[402]<=640'd2767731766402974005531595327149197115112194429018990351835665817194042130567977676841628914365792000902931246800890255549844844624771699849762215956899030953411739648;
G2[403]<=640'd863794963221439775613576526085953721565844863489929851863112478449275316692504628020147036374945335548516592306109748132617207006539736834574450942106008846300348416;
G2[404]<=640'd226745255244977110479942984312888166397132288341501640866317498447525326591092500669649121318043608510614773781109630488465828116088264256219006550520509837200064512;
G2[405]<=640'd57585657223102665344068785441908082893420897918109050259951152995687711786911442458784988372955183903820977739351084491205806823849655179739210293429053141356118016;
G2[406]<=640'd7198258746132696440040734551760941211706415602133085812204446397677103675688928231898053329036515984657924978477410289570658013397472266502261137582774855336460288;
G2[407]<=640'd899782758882452129846707669018228556405029589560107058400892166282112726934714826257074659982432738213742952141018750701300185345346624771727219686464273720016896;
G2[408]<=640'd7029552793961771891108730088707715836096156447141512182818308472906340845745454867779112023009068065305302711440097562176969755658724351098615073804113607131136;
G2[409]<=640'd168715917594290265720708165979837368823044123204198251392377919465028782578614633022764138658690694672490338012614109664708389211756633647257769813648719722053632;
G2[410]<=640'd49206869654028908664329781822854624126934820155492604327043921569602924337350334755882492017444429399550381257978269416855074852218000704138221883538824648196096;
G2[411]<=640'd28113169487306397446307668823927839443198504430892712348047704258146554822059440782779642350914749972895870560310956585429101266755268058308097918041861985927168;
G2[412]<=640'd7029552751599494621755562429749616104056656477456158232196843505728043407132655829706813642372317988217425796050975683060108828365688299447364805606390682877952;
G2[413]<=640'd1675010629071469186641056161393892829098338385773778266784358086230228009216874515308786433254864878171951319731683484982623710027538053835720940690202939097088;
G2[414]<=640'd110641225104865913723027999334204914571533266922213934776772950265399498447708726754303441096755129965161301013311680843183630773367325451528428420317663199232;
G2[415]<=640'd205943929803918291449460477521087363193211748259389957819322793873395817887417514990042003236796942041065139380520583660367714905708057515753652874847868420096;
G2[416]<=640'd54703538528396460601482517353118444190508130918678396132421891733786226108768476948709980756772825338997715639732669544308216041865454519412227010997174403072;
G2[417]<=640'd13729595313867878398915921055528634010953059075298691804774264985116164887447608968568513604825329360274972134173964959332433228172276947794487945581616431104;
G2[418]<=640'd1716199415032646498299679425624612252421342753202071575924974310015487375508604408253579236277344842319182342279360775991453401965952159043108516953422036992;
G2[419]<=640'd837987795841699512360999239197981218694116332483521331274352637053688833159763208925406989699705656774959378930168351552602499843305128667846498815311872;
G2[420]<=640'd19182998509440646362117232734105906683543094102589506359705126826184147409432713662676398597969039568392116008194301107311529922030102581670204932096;
G2[421]<=640'd106581994680138257821170773257517066429705946177573397360309010833762727792369558744682023243928320136305679872403887534509250855068239779891517600206684160;
G2[422]<=640'd26815615857543882786409923837149905539310004875819395414992178312350212588720760098480680655504125058712995109382720330933973751800456080559023306074750976;
G2[423]<=640'd6703903964970512795129695598652567765452751433603417762726784606288464270699763720802750884832509036771456631121932577545642587580309912239538841820594176;
G2[424]<=640'd1623555589537188622827788441298826778107402528017773656792507973915958176115706977201833819396900823956482012460070509007039053527811710011127423899271168;
G2[425]<=640'd55546135161926768106176192132842808473534593830393054381844012604821280617783628726199986069466662424514491912493965969077977319682525309384715103371264;
G2[426]<=640'd1523213354315020689349269595303163907987190583618082477516237402076442361834950714270256939129658533315046434813280994714780179268175564122198443556864;
G2[427]<=640'd26187124863169129488940588990069797186297186603758457959401761217498990226001486020379619961983425408891524616204970593761990974565383317125259272912896;
G2[428]<=640'd13093562431578659734901684094504011389740014306331530158054089707964043949989953322405916960675956942941457223107777973380897110405966215593064935718912;
G2[429]<=640'd3273378309866472278500774320617438670364656627937194556035169290831780415052165553978591466427282685360656003511809472420716684470747703816547578413056;
G2[430]<=640'd204674322000551817293690941442712663594057980867200026935484535621515972815682438353165954258083692110652189734972670186890580489558866044855177445376;
G2[431]<=640'd24973988402516582057398198793178160987452213592773099050415056537560797603612309859652527462400430800521620970857071644957957115218334414809333760;
G2[432]<=640'd51146728248376489885777132752966319099343434898679994349140424469918149543697242236701674705629815558242380374061518850709990486299882123950618050560;
G2[433]<=640'd12786682062047789423777960664390531040470407595762304816430181088038189674369279288414702268656516976467591805808739994548545151031151921555436470272;
G2[434]<=640'd3196667632916776515483105737306152258304807108195610310142927389948504320793033792727593525332306203470067369015817876486505010959317505926399787008;
G2[435]<=640'd174427700260535484454409995558775480696895791352938179513922843375555858473900457447279767827098646243735356985659326256207974739627233888960512000;
G2[436]<=640'd1466097668673159735926663052971101491612314573097950892521809070832490626253472892056901295379564281244369399088376755362137792524253441032192;
G2[437]<=640'd12194330135550370081628357784673045778267093591158376863986609397782624917845470717960688586214980538287652756101781027052567016254991027404800;
G2[438]<=640'd5511837283788254421385329163578897354643366328466019007892039976697801876763329028968216501558382486222187642480852307746642243091976077929611264;
G2[439]<=640'd3121695520162667623902862751128142796956119689919215976226365389262856214903677386521166473154332605685179000896538108179666093419634467073425408;
G2[440]<=640'd758334913956155339410324522374072381401340783185913607482677477529680105839042855727424625255408767755238766414017823617651332055112696750669824;
G2[441]<=640'd182914954120077669807515462683193338227483799358681787021180417410415946652808101549891001520795282554357674747849081241624725354877557252554752;
G2[442]<=640'd36582990824015533961503092536638667645491384484355130674130745620609825064294128360784837145275296537029221849078983862056030964991659593433088;
G2[443]<=640'd0;
G2[444]<=640'd0;
G2[445]<=640'd21778071482940061661655974875633165533184;
G2[446]<=640'd65334214448820184984967924626899496599552;
G2[447]<=640'd0;
G2[448]<=640'd45498746942158376823531662710172809431928012800;
G2[449]<=640'd46624053413417497702067085763764453759452071046146138057418857844331388268056766578688;
G2[450]<=640'd15541351137805832567355695254588151253145047330982434499375513180732554693542846398464;
G2[451]<=640'd803469022129495137770981046170581301261101496891396417650688;
G2[452]<=640'd678469272874899582559986240285280710077753816400237679918696781296365993984;
G2[453]<=640'd355713524293459643974404252608769348018815418810786612808440337637902899709214720;
G2[454]<=640'd44464162267129419042726583464160796784821703584684468588144940524372210195890176;
G2[455]<=640'd27790101418251544025747717484995636021949039966835926073793760460882201379078144;
G2[456]<=640'd3242178891714136715403541298207443281236101686359635329639207548827559044055040;
G2[457]<=640'd497323349422809205664337237748171441127556494867906959341956074376860018740190118936576;
G2[458]<=640'd923491572736239776007688205621369224794710674242289550539758604836844045161523779305692134003450091895156778205184;
G2[459]<=640'd1047775657723002353703593392490229966418231880728904146622695342080;
G2[460]<=640'd421243369770776117191986708383149396995645111076943482481371250688;
G2[461]<=640'd3450971903502377970092160189047817747540850290210418873094766113849344;
G2[462]<=640'd1763396507541813330823728637376429109542650678141460553463892669248831488;
G2[463]<=640'd35835915874844867368919076489097841541703699533500557784095158608790385643135203998890281299829682339840;
G2[464]<=640'd363148590109069717659969773082973616634517417042783895340709839821654497096626732693737376886382991155882167555116236800;
G2[465]<=640'd3290832945073043683777322166267923332873347864995608589133414400;
G2[466]<=640'd411300375809017583180541975031926789551107591029097915754741760;
G2[467]<=640'd235872651551346334515097161311766805682307576276027526773512893765351510149509303255382920323603672971341773439422741802813338166214887780108358342188355630403011215360;
G2[468]<=640'd3685524239595394424287089428429192857479364847116424799335011575275877090990080384152110225167954195031789900001952798127511220825227390363830060533262061431825629184;
G2[469]<=640'd64727672327610783638048341725481295396301880319856995367090250523474968840748190949605691326442749096001130536057534520560222350999438035348399237923718940246398730240;
G2[470]<=640'd1509216418910567562248941993080757920732889882578644878339928850119671669595906523425723218305156916230068209569893770633571508394641141193636226780150066639840047267840;
G2[471]<=640'd1509216418910567562248941993080757920732889882578644878339901805183991914672641608625725816095951043135715937198649909230092955841715840580642066413281902592233943597056;
G2[472]<=640'd530713465990529252658968612951475312785192046621061935240407570481892914427381952318641079567040380454382179411005230370690291368236149029447291925655383631491542024192;
G2[473]<=640'd907706530694132445583897298189532084751843214137126917331706206030471382207708348859666200666191849326585428487490462099110647035855838978666367952005418993782289790407978906550272;
G2[474]<=640'd556035086230054471676571961812622684818635665721320638444875738343708117807866555018008558228676181030535126941639975075535746715900662983244637958480189876486130247043377467460943872;
G2[475]<=640'd271959250384645781579658618248238313503419445804477940079173309443976844109423184577296720259660181141517841323128617893859473142214695073486277634364198318073555656516922358135756161024;
G2[476]<=640'd3898569871989872523100269167449213443684835812701861268143662462894260168990179232120811683892341190911249850737180737908409357795690671724828267546195147746263316217966889276908026533511168;
G2[477]<=640'd8493540452511685536852990364146478672238465743387590345736054417185761964710948261354799665769726401757289645018299299388685715543492194453369294722246131174706735015236652245188608;
G2[478]<=640'd141310488498574733605086743626626603593474654669341019677177810418996454630422671211508560441853710721374603401379991058073102569353424332149189048816227094851185049626872523996266500;
G2[479]<=640'd3992135544809721752245443513906446076859999717053895201636773974939114519369321708078590136155603354459041768719984881871762562341048480722229274127541089838896907548317960850515081656550687744;
G3[0]<=640'd4562440617622195218641171605700291324893228507248559930579192507477944065794863582909201480150545800289163001737779692448792991718485177888830404147442394227449287774325651820312408310408839168;
G3[1]<=640'd4562440617622195218641171605700291324893228507248559930579186828400661196967218489981954455041920776684341453399828328004558266703071323798637124324302646184240693414766308486488091186959417600;
G3[2]<=640'd4562440617622195218641171605700291324893228507248559930579183998880399641716858341521460258749037542228567356856891066642009228429941380033419391128986961505543944099329365939081930894547026688;
G3[3]<=640'd4562440617622195218641171605700291324893228507248559930578295325666595773079297445722858579360900763031005653100386366683987074137944992491500750990800433805718215081822789099843664952296572672;
G3[4]<=640'd4562440617622195218641171605700291324893228507248559930578295326311062542335315578658667804555518701119575393537998774960028041554647642288563344610115058574417230211003200972034474285285047264;
G3[5]<=640'd4562440617622195218641171605700291324893228507248559930579184000238936408417503344985634090004215440867810829119512787979343905198523862020510133544185278736141529050959790730494061596781770976;
G3[6]<=640'd4562440617622195218641171605700291324893228507248559930579186839452618572957366361271048641544624927679469219791853347477477199194761189722857817290642152104839241317637037399932544034354984992;
G3[7]<=640'd4562440617622195218641171605700291324893228507248559930579192517880120407512438254133360521291582681261273917834009041164545663836435539495357801846089086469061348602954961176434101262208798467;
G3[8]<=640'd4562440617622195218641171605700291324893228507248559930579172642330495161922349596686067574157515542001069852312430609191466995807327033051078024818888422179475740510612771025737402016310150080;
G3[9]<=640'd4562440617622195218641171605700291324893228507248559930579189677645588321411931159706720738323668948701887539340453050240277296616691687978218794526879502406467881906626885603732573145890998208;
G3[10]<=640'd4562440617622195218641171605700291324893228507248559930579053396416410312314844380971907212325310521782740231442012955610057338233452824998180782998887138782896659939371343552884543737475039104;
G3[11]<=640'd4562440617622195218641171605700291324893228507248559930579056235630177112042958008639857968011189353000852037975168376264285006336656376537773709659886158541141376109195878958897491491503931036;
G3[12]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274826513084096414410763589535643631263140198036365905011480626256584416557030741986279073966737174332713517466611660152045084;
G3[13]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274583942986173625435122786628423598335195351298452009827744096193279379471038265717377217107822523227589365453904847906537436;
G3[14]<=640'd4562440617622195218641171605700291324893228507248559930578829098515381431878070827295952988723008339682363211600835695245449636842345181393017121672511029480659873913543204176043083802032996316;
G3[15]<=640'd4562440617622195218641171605700291324893228507248559930578829098515381566144977651185966016485429061055844107204432222158198912317462481731717116942175199261185667737948075048152582155730155468;
G3[16]<=640'd4562440617622195218641171605700291324893228507248559930574831474461468658831790539112218957984792807693151295863870966131416891017205318938708629282027478679828498874806524175796131748455708543;
G3[17]<=640'd4562440617622195218641171605700291324893228507248559930579192501241594859402152918351264447016569567893335803726236772000115947273321535345528617494517008660427287275840129138627465728042727423;
G3[18]<=640'd4562440617622195218641171605700291324893228507248559930579191985481708788677517724169557847782148886412016030766795085213178887790801458443066498041185867532471119738288077332989265294514977023;
G3[19]<=640'd4562440617622195218641171605700291324893228507248559930579191985524992750023215596922268832699220739286483999902034102504626897855151306868265503279676632135726688284236578193263823229609244913;
G3[20]<=640'd4562440617622195218641171605700291324893228507248559930579192505745811419316897545103288776456346944130190266283910131513168602286871303553316811473270398661845886152940875225214673089186495729;
G3[21]<=640'd4562440617622195218641171605700291324893228507248559930579192506460571907153556509162675028606303802121656881350617159711376603532929556310466472949496639795817206399278965758196424016730783487;
G3[22]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274506152708596257313859402063367007602481168911443029469420072580163592461425008376388999041554959075417358870849168888070143;
G3[23]<=640'd4562440617622195218641171605700291324893228507248559930579192512353919913603622874210155623707124337869538746841369287713988403227056710425037934220467025605878180990240424030093995705165102911;
G3[24]<=640'd4562440617622195218641171605700291324893228507248559930579192517877613685223358520415456450503753558345545144922220840317169332997823709031021211139722414140563404220474396114446908787332743164;
G3[25]<=640'd4562440617622195218641171605700291324893228507248559930579192517877613685223358520415456450503753558345545144922220840317169332997823709031021211139722414140563404220474396114446908787332743166;
G3[26]<=640'd4562440617622195218641171605700291324893228507248559930579192517899272192456817830387217527698485252308963081752521068045201923801796703172192097918666000836805015955578450789628761587134234591;
G3[27]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[28]<=640'd4562440617622195218641171605700291324893228507248559930579192517899254013417676098550746350027514351105367800623739550311671595959926657012933099356655808133517923785245142031298073444780867582;
G3[29]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603774;
G3[30]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603774;
G3[31]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603646;
G3[32]<=640'd4562440617622195218641171605700291324893228507248559930579192512353935778967047667349084443031203992905768158821961256969729543492132822387001415239773401979972838479577843027275730534281510911;
G3[33]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[34]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[35]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[36]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[37]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[38]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[39]<=640'd4562440617622195218641169703977038192163406479277696854459321704294441441736742775058206828170820819359884813048799298256075373278327082652408942294701053015211957172700036689075883447043489791;
G3[40]<=640'd4562440617622195218641167831737866503351876265693978942310301600978054750768249010299612565693209007629790223446869229651921163253000407234407761549137584263459362112926013517386830542851276543;
G3[41]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[42]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
G3[43]<=640'd4562440617622195218641170662151874077248010373340799263688204921782494455128390663718993040803268688829800668908313440079561821839905196605650692874742830488240734782997942671834745924359290879;
G3[44]<=640'd4562440617622195218641171605642705228323075593548585037680811950105743044094412853602223139987939878746047264833510686528558901749856450342143593862145148382741667638340955955767800094900879359;
G3[45]<=640'd4562440617622195218641171605694892628339776671589187284369969339668631530666715086546191904630237194681836524129211558487364035692795532905492436245574364268985401514733454731865835995620409343;
G3[46]<=640'd4562440617622195218641169718719078914122552386471269436444747059438664958988463198402762688505290203704216266510231818481304933987187922616330211434429899225855678393643139233734852367548940287;
G3[47]<=640'd4562440617622195218641141413972099704277334117961924577978874898632745774128118110403666010659356502071528098189751125649483471488615698059438929426256641887155770664876598991356987948411060223;
G3[48]<=640'd4562440617622195218641126318151193466397001608593588071352501514844630169923536872030309863827422693992417276052892275405478207100875068832113864072706655090740403937149247757730350399502680063;
G3[49]<=640'd4562440617622195218640930072105102746246685047755376681370173834941168515021261309302697091370978302252108797463183037149566050745373469112179076002305899001523510742568173257536080630945677310;
G3[50]<=640'd4562440617622195218640930072105102746246685047755376681370173834941168515021261309302697073453020364829675113003644792602011825772209491234982796802393091291188541301280610210516134458088751103;
G3[51]<=640'd4562440617622195218641171605700178852048364927338989667116500368352803424780719838590085292428056103839125522376836431293536107449946689975486823297344133981600607316868039737203352563150225279;
G3[52]<=640'd4562440617622195218641141414000780279717546994902341760965373032983040093257292828939683327434756966648308833363035010023395775702946443864727625132667094583259546825394028275635003367987609471;
G3[53]<=640'd4562440617622195218640930072105102746246685047755376681370173834941168515021261309302697086891488817896500376348298476012677494502082474642880006202327697073939768382246282495781094087731445759;
G3[54]<=640'd4562440617622195218640925826397149874606737201154680113896812054541503757352505465203127924916549154409230830327687247218507461885230424712997809867771815413548527396041029016850481194404413439;
G3[55]<=640'd4562440617622195218641076783972764202607517185330522400884644578973183158342724766357775513223347671808511151809535225038491903229533862021332771370509537236792787375642670521770929223551156223;
G3[56]<=640'd4562440617622195218517491297880925545107662866385609372265812747803606001807204621373563146147412248863843151022440345755023307286233948069431991689118008503856673540365563510674794431196954623;
G3[57]<=640'd4562440617622195218517479987197951166697624347708332689339994963422700210271555268257647279171282589860734612907714562981192361233561069622108598389126917744538005044991760163240382095981281279;
G3[58]<=640'd4562440617622195218640205470398138263203403504968353537370114638494559667469938595352668490176563787922940176204652665010274757301413566334941215813416489276604944316250875437891516608272138235;
G3[59]<=640'd4562440617622195218639842933208647948187924188104598443200149448149490947947298342931683278879697716773491879295378040020698170808834110924991872596916271947921525702591088902039702615669866491;
G3[60]<=640'd4562440617622195218640194149426863358712574449440147917767471185978503800474485759488338902525453926973657432409077540138854977676523904568833768238718216908528668524619573525294820643777282046;
G3[61]<=640'd4562440617622195218641164057746648151702461796872241137300058064634781835672198238832997739912685091360618072680625208662795985165891121695489950053073058600313584926116783747704551084535054334;
G3[62]<=640'd4562440617622195218640326236734390103648444738326988128915792399655006357298981759696487405197353896944560096738195504873110020415691832797052096422630692980225530975707814742771353454175584255;
G3[63]<=640'd4562440617622195218449854343479742350773825047098384027818365785436884422899704051955103410681886523490967604333844412245762519694566014855281464769729116771593055913363575597053918689382891519;
G3[64]<=640'd4562440617622195218641115102683014157008151191346591163677131838570560079784326727385083222580399582730313687241674764779616538280820489629627417662262270322000268318077875000229022995532742655;
G3[65]<=640'd4562440617622195218641115931519702308747156833245035377581101520209165264418808034176886614604686349660308220142182556224479388326845677379575737465513826392725432647422494448904251572832174079;
G3[66]<=640'd4562440617622195218640673331230994947078198305216223619980606556441546811371942470661661693525898082689394714630574400387403175355333962861794770906282044747343611957345644795690088927330303999;
G3[67]<=640'd4562440617622195218610495942080091189474440651900249846509661105563285744306885488242108508284179861386187313189079095842687216585984068973558999494201143319844398745055137771109274028890652671;
G3[68]<=640'd4562440617622195218640262302737517436558483250966403536879892580473297741739503523402143166999248374395564584886427697820508066969012652684000852046749021722418157148947475741053883742546821087;
G3[69]<=640'd4562440617622195218640742264887353035191425787249504510449613396304650371708351624906081981891684078831737588524623603966691182564591984240648510187411340927824141551866906470887343050419339263;
G3[70]<=640'd4562440617622195218640976255582092029717118954455721420633253463872632548326547364012565592329688020883141729107683638241228077405226937121045590772533603804167678630671123296879479341048659967;
G3[71]<=640'd4562440617622195218640978242072274605126541103413541114957193760769323932937795656836497745877424272613227115586410771622038397902908830939904301321367645419074588702089025624299279940092690299;
G3[72]<=640'd4562440617622195218516776514609072342557845245006986283116689188851703645353166733610124957355299160992878078285492093186461300186732253603591493348425418026010759883907927502252416736484655103;
G3[73]<=640'd4562440617622195218626651300041678745297791845169869076366954187331568452647893334452331806116595320006248787348131063498776462929214219954503734435174439058307763332259366960318995495282278399;
G3[74]<=640'd4562440617622195218629549703183914387756333371003839457589886284026117515697993320465455213663281585821052107355688508590151155579202995766615858704822827839314427857271190931665696481123237887;
G3[75]<=640'd4562440617622195218455307730240282434020547218921508901732642686629889855512207484803087247951135069845656328741698753215883434885732640948294730816259329647296105985437314705724175725214302207;
G3[76]<=640'd4562440617622195218634031740537845275889875806288122510926608800663117777332230231878945467757794642033158921985128092811005431557439907341648072884195736737142337414059316823665702564263886847;
G3[77]<=640'd4562440617622195218613730181418807701985802364528359680990339384112332909741594528739387071108828899891101351125913067273119684904252491598817075839377361521972237827558280181699762131600146431;
G3[78]<=640'd4562440617622195218582811050762851339765308151183932047080465530906667652644240433633223604134973676689729908815795329272233906243054160998665219490825630193244536411585103171555394690356346879;
G3[79]<=640'd4562440617622195218638760957717362481260177261005224077322547517008796486287340065605988234322504928296757363123202985008460896408436450131488974018000016270860323963854147565946186956820971519;
G3[80]<=640'd4562440617622195218637880710473046102195093451312934675383781757048690979916456504434153332562952286311537171727333602141163254220983104778810871605331973298490116260388630016930047641637617663;
G3[81]<=640'd4562440617622195218586694458097992814820671916424779990219458133678844836160340171129173626718772771809391607071251702884382241813307190067346427450666185563645963598271508804942323505845764095;
G3[82]<=640'd4562440617622195186711936132777698707590906580435033301145465660872926144410263339524740925865483523116252878732149390016047686913183946589072398822570140512471005692575367192120455069259792383;
G3[83]<=640'd4562440617622195218637363677642439443109195384600014197805920807079470785595165909848115593946683800261904435519016470462318652206010160460634251440539831108885060184678186342608360206604697599;
G3[84]<=640'd4562440617622195214496681550009771047837196342601161267766256748070158564174252748686557035784498252863456970407783776015330548704574495635709102341554093010903386917181959291003400529131864063;
G3[85]<=640'd4562440617622195218581455254761733870691372328801072605920905006294535578946164629313470335708541553415965711753687344126327276813143383090778818478574420412433206118916289598200796619439341567;
G3[86]<=640'd4562440617622195218610378902785566163614951603071097292501604814637780579982646345724417323271973715518036388903533350386719326935641811452973588131514007291313803380581634040604674757461278719;
G3[87]<=640'd4562440617622195218515585458089504895030885710911155430804278724082214476987103160872613364058160677868828973863141176270324470299299457910735862558085831136604994947832981898496943877036965887;
G3[88]<=640'd4562440617622195218393905361588408811954095373703247140601275187577161606531540077221270655903382569945726501640655879512018646577079964646240353900785993886380660974307889970874384207721791487;
G3[89]<=640'd4562440617622195218610315688914950402797301556996071050892443096820667101364344508171716971630505676251349725240282276839698957482031097381205536602718351981472860489943248952593196829531701247;
G3[90]<=640'd4562440617622195218390006858403568104818848566776201751587302849097236080078606566247275036149838795919126155700232305638599705807827771915133217686560307617165658907974887186552630362467467263;
G3[91]<=640'd4562440617622195218390021954253267390984257532992952635964398492111935428288676973272718836111669507182320235394134394228117114954846669344722663435523101317958548503173078703714425198692270079;
G3[92]<=640'd4562440617622195155274395128335404105419770450291735355854570789199366811222465777950905712562321381615624944487432711479382581409711309411089587879539404072516915196027648381480168994279260159;
G3[93]<=640'd4562440617622195218591415685091444123705275851652810664972497781684644581943967659241231017997339543354707124383115115077270614171134325260213780357759211723819019501052109097014256432266084351;
G3[94]<=640'd4562440617622195218591174151496255545058732392159627391946427781008091339336652422234583372538274917025658190455957599532902487205157807968751130635045887751109039950969741289227401637121753087;
G3[95]<=640'd4562440617622195214880976595804498955504651117371737435428902112017243389274511054134180280226591650476231364529302693294099623987325877167035854425152094826114039875583104683118834338815279103;
G3[96]<=640'd4544618583959608517687239973867589659314824102259629582006497840953162663837720973265440833682828358111440270404473325074471540371836321154159600603108365930679185198924495488434101160664629247;
G3[97]<=640'd4562440617622195218625713458374154492399604235836759629865812834054311440329601659837685999058909675164138321739686296745545536048751645873986522689980120211379957737632701698821527232680296447;
G3[98]<=640'd4562440617622195215657748644898773094932095105923760805676620996334281294636394890031023178475003657723026154997823142169188456921738167050927763332982048537134955769150295555205536822037839871;
G3[99]<=640'd4562440617622195215658714779682686321931898791984811134251707005312520278613511897701311674024935483472805299133753049980893760452465906753805726541126956331697438826666124751367887464689565695;
G3[100]<=640'd4562440617622195216924350825841788495271161389113639669109830825132572975984593721121563525705209304895232109664727673948301525645584116974028230068164656863697523412807834238908399483577434111;
G3[101]<=640'd4562440617622195216691512440079717498105882010823994037889412216526578658173722597928640304908954245334329901751621768171145225065344675789805808272365482548128794847586902939037530291722780671;
G3[102]<=640'd4562440617622195216933046050010730521679057314291012404944138192161562079523809937644719011823728709908440248776752299999446486061849449463787027115054784241953242132622659434554638276147281919;
G3[103]<=640'd4562440617622195151668736361295257537204129836076058853584013691950836083634583405175853395061027199330306407277307334002208108151103332469607850010106513210940724425357450956812611617279705087;
G3[104]<=640'd4562440617622189104757312420776836030838427358348512831357217247779387402623118580521793908112996434201094237883865022838073598088146696455699805024514677799814372848849837803660669137910235135;
G3[105]<=640'd4562440617622195163362826905945481288251453675513146551016119372476733282137068862716027416123898815303928742208133990457048490213885212163157025722534187200299249816729590933397522788166664191;
G3[106]<=640'd4562440617622194102856922928852884577031442151709012432405942080381446920760792016609039239361929114997807444814262806413065207127627694132771170174087837498452928806742389696618920535002185727;
G3[107]<=640'd4562440617622194110647347508065300242650885275415895298713400934076663045592988618790895793071081229269037424923804969287894791829841060854433969631806140909233778012079300313053623694869397503;
G3[108]<=640'd4562440617622186987533717351416241988442830998471649837132658729584720663000741438744207835420405083760372940449254270868978601305341498570762615488362857640603542672106929352329302245552160767;
G3[109]<=640'd4562440617622195123714604177493413362708521720363049013720453710046998407239481316497147929961438537456903464061079857919165321785643391164824884926790483987142319804040738477735236595580141567;
G3[110]<=640'd4562440617091053965022323772789582081694702284695283255188771364498709822968642541720994494534369121743014581373831939101861801498262388652578378659917725796949625829152598854036080398612561919;
G3[111]<=640'd4562440617423014957266472098216754305053347541816101562287096497911981551331907116094959583102691085843468829995290241106536604014444408346876636976366473984605192381320809716606597518917107711;
G3[112]<=640'd4562440475277212637230385091014750044336187882501771931999818046633139943520347668466863120071302019603915229290106184858852661149535110681681911215831012397478383488808983424587646740182597631;
G3[113]<=640'd4562440616559918726474975191417369471259542401407138322809568621671519971522590892980711948356304939180209254358548174741240661021856381105001251838990915961079046857241925760063024397044154367;
G3[114]<=640'd4562440565554072847261012065987728128029207711685669829885442688738492705643486491995743069948276054427814316417267192030490910305978211452122788367356049589024869247001816113955837209743458303;
G3[115]<=640'd4562440565570667870342495005117848073902283040619759096174174170736532849538367285702618893781421517667357911570960060585965801543924102297575871554799865220812837688021634574568037515601641471;
G3[116]<=640'd4562440614435363209483135815787657054450145407679672466646478177317179887780095584430199060576437408809762817153305426833013068224853983010643211636673979017745781806891606597556637127174782975;
G3[117]<=640'd4562440474015756358546469562187099452139566851788836425210285434090804451888303901251298154018409267625834310763721616145939912867078634835203967221091529739509659287435338370219825852441427967;
G3[118]<=640'd4544618347138451919131026665694662159486386865100145573719024620806913894144208939030497638333968183459737375741377263314825135484172135115172769505713292835635837852505355703661312176191176703;
G3[119]<=640'd4562439531179426859682773501021586529290190211482621661766785076804132025447627111301714565770329103415886076251223265449419619483614516700217032911586549172214310362499377695279629211610906623;
G3[120]<=640'd4562440175779698634147303151596635692474698403590177406171453304530236456144373863877630182691559670773805271008986983908461632057679747679683379252360272803272229821931841434677044651837358079;
G3[121]<=640'd2263362922632747593500495008277587779837564616761300196069501664385902710160559287234234853366919863765341282839579757505676347979404804382623016133627304475732152509133732409039633292801867775;
G3[122]<=640'd4553529056934637260176265024244189333812236319662631548069028620855781424018983366885759479383267388823700856636268109840630848501378058003650010204305898069944761263195839173105213363013550079;
G3[123]<=640'd4553526065569609700231406663536792127284776407040365592062880303130785036852527745144005701186194516405321799085182114519666795997802033299727883317838670666664004896883151079679179128762793983;
G3[124]<=640'd3546517121138839303265841628403746209554047894493046761442846443410395743557682948527896201795842621080012078124279078454858575147917920183111040348252125697116462652746242449685011057480826879;
G3[125]<=640'd1122666052497345478352097966980366199532583488122125162691801292840728380208564305842285958533532557322850326413752809075682966620378497807170921021550066112407718932631966667252032163471687679;
G3[126]<=640'd2280974506658676415151579951697573064569418068364182632807756146444755357447890005886855805271884131025288702905147284515562671839992713469941850828198046068916654088218427581115609766808256511;
G3[127]<=640'd4311820206866598844675700934710525516872977977022484998012798741515833037511817374806437411015766250430407803475549114487480087437351186660903514254644164332183039856440218789843743384530845695;
G3[128]<=640'd1005136042458271874991350820899369119572069254393499663588031616473877190398668856454878540968444307648831814327794318977339633938374488137908863456331042091899250010914717152207329176896667647;
G3[129]<=640'd4045603511281399723429105685020861624386557714119417719809085805465858705093551575969646751066841446797774534106360294892880636352736912001917152931290930085159201862575786392602373072097378303;
G3[130]<=640'd3421856705738149474785661651977711714338298125678274452224954093728508456992608842670445728966695071606988194725792580306918819519880488268321272874062515972463442538335182027691491260773695487;
G3[131]<=640'd22431862262858994542461163421826371149359607502469849526658355455041560854735299981209795408848702366115400717807841739717289018112002051108961507293229546691220232917783965176168447;
G3[132]<=640'd2058105523170115297186990431343527159512865524710689285194791996362379988230239001979855414152824866525101209951672359899207234013765533364069194259582252340311691291377006710620159;
G3[133]<=640'd2049937683991867493054183260709048440472390484490822571018229246115533765986568264295151054278305111932523557827401821058018058306178334800885258434935573888973842493385290656251903;
G3[134]<=640'd2552418084911050234124068533984276825881177450498858199431446266335785518455210701120900771606267051253027446056260645791862092891053820365708521819166991586624111749187018090872831;
G3[135]<=640'd2259135673487454662471400561004461156943244803606851551901978468401007333786826421704388634013958060403712447307367142791088797216528968131712699743913322830542885027155536026533887;
G3[136]<=640'd591630149469360324162925500182297235784414422067552412182412914241741580940937546174124978325282827362472563414322780109548955049895466973208077212179930696737652132207032528797695;
G3[137]<=640'd105358793741118961837255707004953608015265941809997923213074230820873934979372620609212083170738662918242386230567365426925468388493803523789166002373171808074124509761981198106623;
G3[138]<=640'd8702164971595841581967043021663679213440419157251500706085620721420872461401249751766454225020376553113057083368134389140731020114275002651222966855063804751858876923811151049966009450495;
G3[139]<=640'd69617318994479297159441705409258897516664690331309469162606253522316466477471774642246136511330227193867515007491905521947653628313631452414924249592335769238355302708015846118944030064639;
G3[140]<=640'd32418090381882757488467428804668891294215540638791074538029643285933250526815842327086053339610097218138874832019418090513605795757280446330289481559301443374793449213434546618367;
G3[141]<=640'd13729595320261213189896356888304023394604196511280053888778944642464354052241800096048511227458328965537572555593226504857992301205514690441189023169887862783;
G3[142]<=640'd9010046928921419052526139362568603675154143486566684770154400453104856051574639322311117466964356258832348387186486277229800342736643842834543112506902052863;
G3[143]<=640'd143857663094644780336818965425000835700678169285887477572279853629565219883245838067222021982801698440462174414961282210761324069708644813472835002096109163867310529553241532645360539795455;
G3[144]<=640'd28282666584082729572894295314314843318814090274364354596597124072431216253942951558159468373237550158690561262062355417829495886084723155647642346779321744795202299236636841010482890407935;
G3[145]<=640'd16209045190941385042751641249647617817592873864680725671430724610543172582156256630988868413466555262339799044205921221950306700427419832644572368170190438973493435483035023704063;
G3[146]<=640'd87021648743099121449302144358515942722337924604119081296506840152637726724387845364307475476293589132561970025935106099178596878275016732055245219301927398458089125258299534181757209280511;
G3[147]<=640'd52212989249911734167316623967928152937731174921616398581782151003789352147998516093558560180740707293526720446068591961487300058140683250334956373851139316734993260919493177753584674013183;
G3[148]<=640'd1313965177134374515711736771469254079538168780684457823563108907618391323722062977514478759845113136517573639308402260431452758075147199032782906421772550143;
G3[149]<=640'd2699348947116314326816178036795160670695283690140367516582291850354390000910162272729641235526109806111791184405063973404591965006753318158903891930320841463562239;
G3[150]<=640'd16209045190941381443537504021540727358436422292277123749850062597427795937298886801414396685886311925443235866628709673100347318956176978873632681231681278142693258378492172566527;
G3[151]<=640'd780282119339900436366747035411710174204332792458616195779106488573878851091536251373138126480983939031400210462320518697831959714460536608276421717035607763451903;
G3[152]<=640'd430095796747893101809283413968785684693014113787558513122048536933059791181170270173671321662757057859876644799047566709741716966225313431764311188730793912600591901000599786004290113422491647;
G3[153]<=640'd2305725605097154325877995706723926987381498491977752289993605626459458350706906058634566225683922306816343146541773227719842685942235116610171325828552582503321728081299043092584960780348162047;
G3[154]<=640'd2334721218458354953144903177026921532712357260086469766952292242645945858879145641736104363630948963121035433441216479825125657667504012186874635542273467114440846574914818180575579478440280063;
G3[155]<=640'd436674633392871391432598097179574670427822508590106080164111468757262013544499730079453969845159758178862888459813543400847258183575846957936391469521217700680800215995270606658183540382892031;
G3[156]<=640'd512418276458864866742070672664754330867535529757032556202180360299512079827715820647811747617389209629889838892761751823591345775310782285334690240509161278850798414675372936482868700238577663;
G3[157]<=640'd454670710352944290245872984116264505670004550657573163080916922739614887256183958365218424474791521747546481838761452094925980879218742005975722607341256090990681226035146288621151058021842943;
G3[158]<=640'd2765165101801220444466184305642792134621592176360950204694885449534546631750344574261988430785045849801517796733978204725991046364621667081032419220281725564954737999042181551781229796270276607;
G3[159]<=640'd444489194446417463660840230146107834958075911617165971162058697626230076845787949064812121710490431856713062017679494067116411495425374365302452694266809510191905725149984068920198417491165183;
G3[160]<=640'd231146937384251427655946573463333354826944161197665211611850299873774518518217645649631606014534146112213844042935471101741279662110379711604490752510035434424786417796891344419013411133718527;
G3[161]<=640'd2423239639563984892084043819792299995547561500378327352930038758211157911122495936744407693464755353458194313546867654141274361288788869801898907195734697688190177605056797688595173724477456383;
G3[162]<=640'd3559394285553887021231381074026775513455408488180018826575332050523361769720414257984593442982212803824617517085704856119963609101399780764589610887238539354104946776521551794885228357476155391;
G3[163]<=640'd1962324038138964435321639071279151802573865815495904221521121271170117660776097649512373632766864945910160938772799633805651820914659045827248631628980784444498629532895781347586457222890127359;
G3[164]<=640'd2254715690145168194652278004702546899118216343808875437994420449585944071764490623775777551468965065384322057984588067643850132705962147610272518312132070647292355326837867208658576311792435199;
G3[165]<=640'd1844652412913428400049124825875613972941856563211958789925017875898474924674784494051793267797525639051766827327554444777742092165231863067137442446116819719705717098172244788112482867014008831;
G3[166]<=640'd4055628846859080189521555709715288980578522348197423573340707784747845214126398661607306226358547818745974254998353418625113095608423727535546955803096435650469657725619253624039024834505605119;
G3[167]<=640'd1759916064088277109577879634359419154888162427036906591505802084935346188341231970246728854331592012017635117950920628464342184637060674097629899071445680739055980642742987742525779805539926015;
G3[168]<=640'd2788026504754511278883896727879757266684067960156399377702884111811098472399256641144396549307345000195220170021654235864839778697198313841702250852431321550899369351148301180890509578634002431;
G3[169]<=640'd2352369072853685358294400741888642969125539117251234963471054570701803884547667633529950290974587603390681041986314221687163652579988588266536800122873798430359982823841529877234091253213167615;
G3[170]<=640'd2919280386539026784044869535485588207021428729868895239295607796796165610667907509505517924217535834273002499897229008661173662439070770227439128654857591619467980226377901725869145183280431103;
G3[171]<=640'd2121882792641178108236941072183626440783667832337643191982365939247994787773490170542601568705479900462588260417188851487848166249620272886780295963646851645969893521729865933130994983475609599;
G3[172]<=640'd2108560757521521329614385382659703699942089746222825758849983354582037424366705040749370985505898816218760067937909488691873778876305278429601294002602021782419351532807011174006546314010034175;
G3[173]<=640'd4330606346253728701063782886267418830375916830092080721101113614892911580688361903905136223296757134423996379658055724207399677450769446455902288197659012984110393833952358157490537096664317951;
G3[174]<=640'd2325349836714301151986768699638567976267331587419916699206612987385591951869822486853249902598731158447385109102112641147960709348081731886207676846286784689633027455086658825757201638958825471;
G3[175]<=640'd2751415422106139819407717497434241970678392996319445584698099683197634822555724123835061688327905802440694430929862776281460556445343318959081690695613393820773001398485534074529219789660880895;
G3[176]<=640'd3853023584684560651920799971058273783410898365569865253595851768075109270891288498537291607176906665912752225211163432062226111447980078936297617148974656602316575107116455639081690081769029631;
G3[177]<=640'd431074824305682565515953779615552866200928712645994234834988308148841488296913323597350527940604607774516547974531490767678888002993491955991579782282981905865386149225455569002049662334533631;
G3[178]<=640'd427728875904341936654749589007555721492578494805497196934192117026376185700390112714874953466216973312898667387341447697504792402969699276758668064617971527000448981852790811106710488895979519;
G3[179]<=640'd135975475676661258253981353650120143521698699731363308027938133365954230867123687698549770316464956073846318432699080011546723448363593642641505063070104114278937046572970278203981561855;
G3[180]<=640'd2281220308815247123405484385554785059042323241186731598959938267867034885098145402451241460362958518486305513019840885409203259622325036802042780594855136631965105575350927655120914330333216767;
G3[181]<=640'd2299042342745477578165786312324280238679452674288800642621126006855420278447320518993507132344906132001622337761817905410311049441601378461507702393261675761916068538432270867071976570808692735;
G3[182]<=640'd2281220308815247061572884018634279713491237269298930871901455710187703348669853936529533396113873412988504640227176175876852576291019205874627392253714325666809291415162427163371395467576344575;
G3[183]<=640'd3706983290761251223036134608309704322701945757916681065847583623828251891069908831743354627977946589398611565509823075881946947341263104577513848684589878701118832714535883013559550008254005247;
G3[184]<=640'd3421830463218721171641654000012425320285552849171586836257265612774697358574610825986315230368619081752546026646938337459052042993848500136498478817531697274613849545415235098962645209027903487;
G3[185]<=640'd1037378768555047503068815680561601600335286838548720168673161430128189954729598776278240947909668156627788164313373801433290984365749381507660569899699618026146433275762822554320895;
G3[186]<=640'd518689446110124119812317621558758943017566628519660186391778791205845553576786400879852336848305086272500152766498789228097435976035224451284307154270174455017931636845171156451327;
G3[187]<=640'd518689446110124119798893509757696434435933835591729272056924952799245558774864998552481385648535518094882138171336793436064013692991565563721170483678543740091898596786937031294975;
G3[188]<=640'd259344707596911967815805086870017342551904834429432986797159242237939661637765827633815629311393121418210825390117652273590997482300548781276103012446067120061142574079186737037311;
G3[189]<=640'd251176837502363979566754350566232669762388856225847602126277038384476370498744077952892676059094832627981087359923204676290782566318772502267917034618881454130735530146360836751359;
G3[190]<=640'd64622317257241739899603962623318072950606230237253790896057429598104684489140894361742843443204652494608936260524733481837480735538571884438647864158208710068806535444567632642047;
G3[191]<=640'd20237330897883924355570103926005544203649190053887728892460289368243793324869503635040750833770522042343729163977507992031693803173776649091997378706729658526211567149585493131263;
G3[192]<=640'd12413025918207216386212617081661549720689734571165355591670572921026675070133584881654292394707537083886328792907172898397942994180704353715121921568279065050654740416310584272895;
G3[193]<=640'd428693147428304467972988548567359028247563348211642954354775318026875833716939657550985590740234964058101133591619368486801042132701842749212007957534931992624464941022326030335;
G3[194]<=640'd16142173233643087690794013800839645711121397711717601579924523738096987735014819366311615816007867551290090062680461181954651128791253318440596344613851372819683419474993610751;
G3[195]<=640'd3381470332639991214845870814810049215848776112347780737205338980071621913308925753655280692839274367016682552021164699521162282297633868853753663894087277468205242118045695;
G3[196]<=640'd1982507749302453900662781906625815623877617866839925128755691330244299821394684918107120844045517002425090467116803304675437774233753695291020089862347667302722364202930929663;
G3[197]<=640'd8481609822793715741580003473079157982432618327812781211509211879102880805121437790840860055575517978220015158117399191230940873220586089035235931507740551555912674627656100186012254207;
G3[198]<=640'd65283224674063340415599308662747519912271497631027120241526948021112378613709392480848900565392615547508056087713104998465617456788051668045739622107864794905637664532417583675621190402047;
G3[199]<=640'd35778967871402971923799200148961493649994099599011133664525056005088685832238658946956263636152411104488720506396405239702535560506899648385097848528719911594055439212928249465325158873956351;
G3[200]<=640'd138398856239667182162235364400695610501115042305427330051056983381010023133655567906800199959691012250598735289812131886058674228171782061441426776503519193433132992831995160908444002882158591;
G3[201]<=640'd1140610154405540700137811593039912863283664858013355169737840213631370446204351326431455150495050933490743583147488060488519576563930646649093554349147527001695582255278439060799850284517949439;
G3[202]<=640'd4562440617622192595207697529265785583477542282544468980429516231397850531812289185165198098323458148890763519758128473055809476180598535049098170605141599582005799678488877833049109788079685631;
G3[203]<=640'd4562440617622195155077261979426049988347565948841649770391191531872930575128654643934187026765716235166317389668477827293811231481732264819551914798803213494069483199588082839034386909203791871;
G3[204]<=640'd4562440617622195218270201948776960282895596126874901332583786842094790104958606412743614323047361978266823879174823316684524593569674433060493415129428413662949315112639075704357533497153290239;
G3[205]<=640'd4562440617622195218146537454549745516948206889639284653858984034956709132452948389894492929968704376671725082560110200938122688259082796805503651999309773222054018767420517424178006037788360703;
G3[206]<=640'd4562127305693888521283529400419199968219087787203882977136948895094268898328889845513080127170979944095173203019597815246852341226162573181247509400666820405931300704558817148906837624538267519;
G3[207]<=640'd4562172628761091561777259981096593770502246337390257090637721036412775536983582836009919151165662904127124088155489297980831650582795227870934795782648521518610014119447868821941244837180211199;
G3[208]<=640'd4561981306503170626377208909833390523851335496360183068334935811233181471820823431058729967766882935291087219619152644789162711870456042054105130273109724670755684177145340772984548035712253951;
G3[209]<=640'd4561985385622726190877787105170625349955894237075827638339858179173690431668569132190846159848148689427494753219758944435917146304845732348098665372207016235381697610392750984142653180182790143;
G3[210]<=640'd4562431915457563854441684314731926813800783944214072541615978062833761784369118726836060277114630499244380710802889351017371918118606479212021549969637230167804506332304734411697833770177527807;
G3[211]<=640'd4553512196461164914853120815330183708660027477270628127845015108827126670025432428514696543384656147686186833908802333235309487350602120571605409297441390119395283287825135589280839354695024639;
G3[212]<=640'd4553451281307033087306167005105650817170901356627937808446988839013028102596638888616792855405950459851416327964207011190640878695911687024862608769088925091242322440538699808269198745248202751;
G3[213]<=640'd4562334016102484926173716499777802335038007351023461837252975645457755406231179314915969878783465958345915600061750698443120597351388326331992348809183017949060331532309017997770721672288010239;
G3[214]<=640'd4562352508236038957309431095348826249786495495813786515762037635564810930123110877157233094565364892773488039665076926455089625329185826073933928883543527718305071726432604422789884243292979199;
G3[215]<=640'd4562407984752887490727151963278885735450827081928247197795429481795049576266741131182982955828485593508017380451865631936963780220470461988629019619218104416741071048629916452512828910504771583;
G3[216]<=640'd4562423214350585226036423757571206596116603280299846031646157886785056006337527249410418790125809773420298823341901525391825919029492531186803373187312065919298330177137899996567514739886522207;
G3[217]<=640'd3778262435365781078340615470773487033128302181590652868178401180538754700588616933496763470466864232013744956416043396760728264553278895940341633443522468507968262764581891696054326051038035967;
G3[218]<=640'd2290026908162106872228655799250852636452309870377588158197464225088638483195614171807782305733887949669228060763602581664194646889386391466890129822768881355634045092487488051703160777082666943;
G3[219]<=640'd2646002007094731036131363760387903820933041289227666731990718086756423316014965089809797264288893668567705176488586515716898677178559000905464011642177303375779781223879057918416841599549375;
G3[220]<=640'd543885304517738275772670310699922878925146071199492855061269742441193110893693346889096204757916313677523276254998133024876255597584575554869708563985673159113681420478340016757596454895;
G3[221]<=640'd1087770609225422676872757074878613643576129742895124352637536340746518164829590960036940822310548433554436405532382054433862348012017424530187803338675659479329024138952197796185670156267;
G3[222]<=640'd265416028666389003897977785909172375677516014003394377350847872526248837396134625060344970260320776402661954650402894027766776382424230149330179675143107674882844665372846327178012484304763;
G3[223]<=640'd2715075437672524254269867197120715731941824104550325331798116796819325988381377239280364193879956578744878927095636916044022920954130268486095818480352691568067131093026032129521703948255154;
G3[224]<=640'd4177039124691592904419622136072605180177198516699062263956194797009795361065460133064726867400504717814680066075842353678053344577908342586345014442166938240225606990655406560644324218850684;
G3[225]<=640'd8911016798680750988086231074186175522455201448655615423422802027262487747117583077182594994336093440533155581815187986523818751007114873022544750016486091336884931579213541082377823879654908;
G3[226]<=640'd35644067292009693684847328974079755308053015382592302722930476211706101442947925672191429728600673276262000500824191623248828291694876047493714045665360696488535020110259173936023743454334812;
G3[227]<=640'd2744593183971983875679459936775790980714249291435732885405385165867579386539878152661661121363327177072621961831749780774983420909785840526779718012712200618126272789450935450521569668454433132;
G3[228]<=640'd4428775365086418928038078201958507040666071093881887609489871096089584712907112072312396849508494805684564789222021287198811422134433319124535547156346274054972899949261647837887269312284611433;
G3[229]<=640'd2281220308678329320161566099744396813838544016404186218779416719800629506638861321299059243918664379813959760970930795510567539758141447027544165600239238957345069600142721629829435472589673737;
G3[230]<=640'd4562440614435383470785759011450900070144386113825103121173758627945303911313074742479124846032469545942534450106980441472714592244391861388869763967949815369397252992270066047948009873686927288;
G3[231]<=640'd4562440616559923285268934671920497856797969915271556873503601463652004905399160757833063043749981397434091145641472833098252875450116563772264730582482890137834705963516146987357304667391400316;
G3[232]<=640'd4562440616028782253252329970072029407470381318186106244651315940313514709972414622790617420100852786502697734585287391472941531038009696627911350831427275813221650912513605276075355991875631488;
G3[233]<=640'd4562440615497644260427834017467017513615710594966445964641458460892587184656329327456932370983536656926575251613810309208084382217634049171722584629620527350999656681391117978456485290307168616;
G3[234]<=640'd4562440615597247830072437975953960115552402071403344220618149411219308543066008773394870681564860592541152471891768198136527536568742296271259297907897293254717575973665982151955351392629140300;
G3[235]<=640'd570305072953800132157537190383029185699455559096094925849982160550003360158338326873015741887226548848917547975604031314289205452601446949066198791342196157319982710506581116150969749034674688;
G3[236]<=640'd142576267719983556275509787411579992729854017116192076341115792870423595728043630579092977011947647383799646391022985247484184981639067815972451420394266782828043221019143162824115858446569074;
G3[237]<=640'd2342622749918284661827295149130508371900841289908720046994407137548628769267858964381658674282913085175959821639995657319399691712977033071068562630852067465246508091393554861059001661639417403;
G3[238]<=640'd61541709990086372027107654445106510423810311730297720933521969054534951854600431106137983535521808175178386739259337876738144676499473737336973265915656932137101142074242072538640369012645541;
G3[239]<=640'd17265095110373483755636271251430882508660142240059793236938339319638859116076503127941811914169379489830269978681177359546231894568236676796609447382667243178180281336211123444149056455515532;
G3[240]<=640'd4544618583959608518568354529108769161660843754005111116284216530964816150734644445776063396510380106400466290748910833464140906086550757250038368443967897440613884709021785686006110179664579809;
G3[241]<=640'd4562440617622195218641171605700290446199157253672392422569549304038853153861206809538285607215560391796482284253815450110144115662383274259422309387126786625011119063618821958400221336186050239;
G3[242]<=640'd4562440617622195218641171605700291269974847379643866955855636293206398324268743145936456189924972256299861019407280096712702001277528226060199041572859995272753948561157501349833097419365977431;
G3[243]<=640'd4562440617622195218641171605700291311163633289280796997369824368738668776385162032202892808618385787297191977144778742592649436747579090686162200927121141287262819517514772243323172539998106256;
G3[244]<=640'd4562440617622195218641171605700291324035128799732233716206454929104697820593117571121937364374931168632298949076072147274899398937075746777524141915053891712306633234540354220044692022698662551;
G3[245]<=640'd4562440617622195218641171605700291324464178653490396823392823995223625772524311855804382496130203290613607810984814342428677476527627423800762023864485835568831468589389699571280539948925285538;
G3[246]<=640'd4562440617622195218641171605700291324464178653490396823393205592208319962718316465063629692890354917980039283434781548253708851188393610349402082140023029568875241615601917923883450078927416384;
G3[247]<=640'd4562440617622195218641171605700291324678703580369478377009266957105441049666585279807358100866884263583044020704119071290135312485000635382149983288505738846936933056119194509504840932507961374;
G3[248]<=640'd4562440617622195218641171605700291324035128799732233716950737771692802470972505476608886376023339480647904145610618397186189112455824252550335299413281339738843999424545773527162795350591106598;
G3[249]<=640'd4562440617622195218641171605700291324035128799732233912697128289191285378591998886365240200566249679912130975232201455263165992243605798276986572283845164474031712177283290378651190912730825310;
G3[250]<=640'd4562440617622195218641171590958250602075982892538662658512313896850459227093799910587929003608078740956774562824130133194320776827873332236332809530862438870582528785288594028087842366136960012;
G3[251]<=640'd4562440617622195218641171605700291324035128799732245910536729589858754849414176853543881465604525144527172954260428481977613338792985389198373005806303450215995301912891935492623772633271604353;
G3[252]<=640'd4562440617622195218641171605700291324035128799733453149233922102479484451467885929576182681292541971736253769836241060729753217547075498172074329026433767473571142649063975330586599866464045257;
G3[253]<=640'd4562440617622195218641171605700291324035128799830568795541408673302621327788482712619080476637010058632512855877086608760706819404194484770839003547746975345625820285619119455462667121466347816;
G3[254]<=640'd4562440617622195218641171605700291324464178664876974660647509962105752369747608080516495805768560003476670351945917365649925985201927771145801071678618159159559108133217202806949801800684324291;
G3[255]<=640'd4544618583959608518568354529115524561047264650050566025280497970185145062714710091828832894220667979752315194934691412465678515134883508953092247299801413013146078036681717376137068204773122181;
G3[256]<=640'd4562440617622195218641171605700291324839597381018575113188047104766155540036157783508631235525920502546216537365626215518434300292997140096386777213800330615731240539313396651443521388759093322;
G3[257]<=640'd4562440617622195218641171605700291324889876715099234227551624977580561657379297485954414001735499224482380445973071900375059768971225113780352513166190732643691304026861321637138692417843415219;
G3[258]<=640'd3440209435431188948430971314503259218000947017313792606877671898206409451565012973286001955507159105859339870759867882295230516038868537170153212050793379461226777519357293643497314526390096376;
G3[259]<=640'd3992414009695139388722504334427018301946317537694857987032254667477902705318430703444266175471483911141646701419855438079654796651941481931318508935371424570222600708975789683440173036300353768;
G3[260]<=640'd4279515833227853320754312173279441470766168297365251341850503429990885220140610612622533145656247677669842113566937185617773900594224831726392160223811020552335081369163074372615631286235146176;
G3[261]<=640'd4422092102527708609811687467353746566219968060476174648260805501974955167496575315700687400522652863405462981286973409136477749107731561014451977547630179935182820196615028111773065984841224712;
G3[262]<=640'd4495607991387430336331140035108455891896630187738243567900042831809157644148974486609193772047600339769459855848940927246510675846814586060943436405005203809973146088095426005493993826820949797;
G3[263]<=640'd4562440617621676529689601546910839460085632390086854144939485532399224136054044507341927369542305818900951849451557784105106008954980771888450810362914823912228117322089701813882561988966417057;
G3[264]<=640'd4562440617622130382707738005972697419397848522733565452267273565915365815801814471848437241097971248244031520096475515282036460781322609228735683040735869520145879375253083951042875772975230762;
G3[265]<=640'd4562440617622191167121864968067881935308085871745071320442208264880143625514478813012357564809930550296276454380771473022723412995657199314522254484369009483391201517701078603910625539775598071;
G3[266]<=640'd4562440617622195218641171604030294524358794009950068473617220210456953225738861729106248581256636513522134870236959170320072560139148291429561762867742997751675270621133198541734768897418199115;
G3[267]<=640'd4562440617618175375433818141928977339530384456485100130332304072440959580425971641910998512238993707989880486421100646601793273211814728039499461665750065653512378906951925364531580709852547698;
G3[268]<=640'd71288133853656020111308584941388209256825390836822307792393877301700733844426791034911562463703210116566474331476726641570427634150859083500962950383906871830909965225323631144112187415497240;
G3[269]<=640'd8911015769017368360160646546553737683867911035503069664704027954885064002261280594175132843783416929024860231218665415969194268147572017212555960943210828570586628275592929802396163437086081;
G3[270]<=640'd2227753145547352099710641783617313568207146553186695738450110359128603648475383229004845048122149604842936027283539382527492419574601196517046670420944108849796568891493093658636048518106816;
G3[271]<=640'd556938539507287672081756338868209631558028939075896783285733745492214747500732491189103884156935262033825126194322848152983604019289545917961068394872965584243341735537675957053231242072320;
G3[272]<=640'd1113876738754298693023686937456030681919329576932212014467462830078866936264165478416205265322942821447448389653044613286535991901495278801994309885152658107234637780825395104353165212135684;
G3[273]<=640'd1113877070715544203503123618448659777212221657927910593862237378871029579365377372941071819942486826902098928988282441604732334186648680968344834141111773657906295275156789320074279322365042;
G3[274]<=640'd556938485563585275179646307075435524312177016814600510021867571478544470950276214273085723923648761274596069283395153007572251742013709472057185716228955975184256448737616564182168990757196;
G3[275]<=640'd556937489679848743741336264097548238433500773827504771837016771276461821721463184701725856275901739511016692204253060709483661165659449354660665807695205138132030200063534497355127210055762;
G3[276]<=640'd1122788118618410133320407430081953242025568443637327824507845509920129589546582106949355683224938151167537289756294184813982947693774620713075687485271123782852351821118327448644954878127084076;
G3[277]<=640'd4562440209708216735364039812096548692597322718121045516218678383956075203181095517474840123429735771569035882235445557238851565732642405702081365297103707546969467231316888560398175493739756948;
G3[278]<=640'd4562436266539758063685099140593703247070233423221739510733699005132526136233466892090694365198792638643328874570260275714842350106832721056940443363529443781325243848154417995598913200604644528;
G3[279]<=640'd4562423213292446598816881745273939013601248171141278251197177879150284619730151202409917169939499282776492590088931076778936021896245650234736953337092168312979804623205015729518585557961002044;
G3[280]<=640'd3992135540419420816311025154987754909281574943842489939256795981282905176241031134269118925096931437235971067842226520809099879846619513107286811508318607210812993019504037413996418119007950555;
G3[281]<=640'd2528027624263871750811061352159185504521249427524406282906752694972657907705792127830083791760066799564105281543653249191486546905823;
G3[282]<=640'd11201238980536326930839346002165040276420308822459498338166255815180541494759655844349372168708016065731008579066364098707021994933009;
G3[283]<=640'd11201412272392209481768069653051549219151773599528047707802558113652741637687566073992302522374685173014778391756136761252455182351490;
G3[284]<=640'd2672810262168494886901410360792305454429891738473356872898934294283234058334645802185486838497612693700987808188873414306931438686769;
G3[285]<=640'd1253203378778637678797262298511046598270419659593006709231977512630728594937092620193813796342610456868324856920550976777750216491044;
G3[286]<=640'd10440834316923693455599965912163799570760981380348891016757084477522071484533456758582931760230361858249557448153056285766713529076;
G3[287]<=640'd9704343929422852008524449644500792962028548280636571540147353759566486197510645921382306847260085146071884617487627724899332128142;
G3[288]<=640'd1469514937884031875576559517595834362821311904095228008334455042792368248462826518336288032359497489800904034186413305747998062593322;
G3[289]<=640'd77634751435382816068195597156006343696285438678793010630253794579372475758653095231205201302121502434664298658304078486979408750141;
G3[290]<=640'd2053841025846363391343146398072256870013777038110337978848511808032987745030079550327283119831;
G3[291]<=640'd69205835565255538895077218036211369237781781017298580756611900516745245762925047474464508027768356907891331102569792746534509923012383;
G3[292]<=640'd22713710134237715329666368996500141698584636763344225884267085246733839474152760287573111449662974230669259955255958731172043457950716;
G3[293]<=640'd33374797374098815486198883889476470772314653149266802758551412521172336584716345483841862382630;
G3[294]<=640'd1419606883389857208104148062281258856159651337987634679598807612930599538678993046955750681714133267569325316143490126669919354364312;
G3[295]<=640'd32592547224047760504488882911068065920727054772575055348171867893988962720477326549688868211;
G3[296]<=640'd10086913586276986678343463598954567447797588287321934925647664300666215145465152696923824282042493262808325452864218960;
G3[297]<=640'd80695308690215893426747474157622775116888234548302890633390491687411790602969535466686764030419403916951712921057289320;
G3[298]<=640'd12032891116593492437478087924137957161487158124578483025065002626101472008876912120433510;
G3[299]<=640'd956156419055637128563609460148423571657506200435434046979890293285861219973347761287;
G3[300]<=640'd571134909255340073692148226186575962215210052602940331762285292541089263254459450982856662750004379649175;
G3[301]<=640'd49947976805055875702105555772516416918652829119596474833244372250674846925174151471551193845422719610786682514264684853700641444542952368466643356;
G3[302]<=640'd7566108674227999500707800769729103490481092561748379876621915702025242705325857092779422415778904589511235508176017658;
G3[303]<=640'd49947976805055875702105555796492027848746154610993183464126809628206331789046119782412893891812730962796914277907601209667826689199636264685160978;
G3[304]<=640'd271734629868605141094551964136183353817308535315232765835625488695230408494541303770177647280275498607052652741384257674;
G3[305]<=640'd9017105333094607225022266872455560871021745788125938405691018206489017193899221229655802589429295944751206263868340358320;
G3[306]<=640'd71330254592325858080562959707944973942752192809188920584420469758125510001623189414792595801926336881488075851112722215685;
G3[307]<=640'd109049149918687624569859440587349555726332451463749367841173256151082429178166345335526150549453768865676659692492687500807;
G3[308]<=640'd5546561151626284839170564093712640451913647671679825021882645404581251112071013569861703484178789753260372497876861698230994;
G3[309]<=640'd42141753143201884772499671022941400190706469207746676583854771990908990138165003744461350600945716375620977545174653373311010;
G3[310]<=640'd83965233429217149251021628215008191255949715673842898137720331896124302029233938902533136848286106069094779099296654782195839;
G3[311]<=640'd26154154568885032141741346220922316220052106733347710958625127554367254025338663757398220351497601632132008957169949327579504;
G3[312]<=640'd10243715918836854696465735561857736611070100400916787077763143293721347381421633609908101006410840127908990212770985194053196;
G3[313]<=640'd439347050248359204673795771218878978693669461899215576299324491654173956184091799666310886111298625230318968582264926404210733871180218422747911407521470354585;
G3[314]<=640'd40223423789839985628269908136626676077603164223156013134620142804416910238541168532719155232655513532557680833630096141594702663905973282402251521997423180;
G3[315]<=640'd10404458953625931580302056102642482414543257554838990594679442016718234550780104515268958228471636381815689006544147472762279464999913810997462847341084298475;
G3[316]<=640'd14742034351427755293983378491100207006376430851424754215514237556955767599165379520821893079561312951392691628109490688327446055349984393922168671672852791374418054736;
G3[317]<=640'd2265556412037340780517306777925002060311064427517752279312640585699864020698485367256672490821466313702492029912197153208975118272956874158303875210494615214547263829490292583654461746914976768;
G3[318]<=640'd271942652322184750755106736933429847413837505018877975965805019953230667823069094484133450866338740361001598563095333368143429786751135598643996887678056929681503358158614838856863501963;
G3[319]<=640'd4063423641076936139638052847261902944674294167422105827947077766749235226028686014327205010783274488814562373025665664682612619556286819954874849473000619897099067842269614870997670318096011830;
G3[320]<=640'd10830740992584322679696163104860307087727752005555326578676192217374972059055152928874537094267529030448639010021050038926622593;
G3[321]<=640'd338460656019375671633736840851799842766387917017410441472616970131959125316384427414689757028078659920244569904023082925822305;
G3[322]<=640'd338460656018682755428141562246537451970514292750665074519302380460273099832619828056712532749900974419647474732203436480164455;
G3[323]<=640'd676921312039290038016123432967415997886266085771633623394591486546386230323991919138462461968980090381474177584423966434815564;
G3[324]<=640'd1353842624082429093076842346341223688317427764460626568455744220342323290708393550440120879484292438014942765600173513114938899;
G3[325]<=640'd338460656020606719013161331925791639848382890583691438329236359190793886582670284411105147824350865230781061755439170349851248;
G3[326]<=640'd169230328010303339543968475616751192048579828285566520692316967088577214931718159500366398223643929753418100103626969209774723;
G3[327]<=640'd213864403951040400873804919017201155854370086277276246745899649276531167686781913486860363044006514416215304017516217784213312791577594009785054442546683066159739629861433204549689991095147531;
G3[328]<=640'd71287845715177044676327586121033818201595692588240075963018350283599424236978192743352119159037774926054715415978117474412209894577596309431029624910254811234305277428681752528381490661034319;
G3[329]<=640'd4562440616559919232993028384168798554702324582113172130787255397408790822182428392453384009211933469214623818356773907777723894685539899922169441491464323345634849039428203355139346909539630871;
G3[330]<=640'd2281228468152943197180176869151838823522374151358654827229265984752460062704108103422229457399258037077434716295385005078636097602778661166271598181027138038727563817523895720619065955736511570;
G3[331]<=640'd552478692457750547301255022039969164030118185495126974321314996881759882596615796514220023189877564986900704781014117451281633968037169583319976212018435325520495720481943078095192952253465352;
G3[332]<=640'd31205963239275344766221943317872263208106571294452508460038695259220563871268827088103240556212758031892500136607654635579799421997992462000510816131395326587871220456970324717076547719418510;
G3[333]<=640'd4528885069866856197410320703693035153955140492415725532085719256639389618679231580658429451161626501752120007798507749874998045874111802794714855045578684959168390480397369335617245958491751662;
G3[334]<=640'd4010079404390255959676466725246359945859910242249024453344081568143123974714670304134015260796251516371954340633825453387807033295777520089000070180577125237023603999437544217862149504913122947;
G3[335]<=640'd2210192695221675462024156344768039770146988214304393854624498010409472154261200617670456106232563091295065370089805738962696364719472219563482612239520007942624840944383685335095022603615083234;
G3[336]<=640'd3341665848186290526668424386952241617297350714540957383975082664674615074567548521060513871479682459142010273864975261788557245567162090619269464888548903969095512318105964938250468266380645262;
G3[337]<=640'd3350472745238062407584621298524526788013691612080012822605375390908915403285560167089390474484432352157811102010458769220521109370031375551864044038986625446319395148171561633068436944689067667;
G3[338]<=640'd4544653341628871469656954315296979568629644854362729357792549605373161891518810676117258361199738449431390458206788631163281263281168346613026053167748714021502832724371002783666880766492678321;
G3[339]<=640'd3203545096030782437131072027614975693555824818667529865125229456257508182001332370954234170547239227048861460390195278078048902715743232991679775892958417658267043895559959527443012560076547125;
G3[340]<=640'd4544613162099606363841967550401356243598088597926296113902734187001608002277509016762981369722390850521662700523343418793417195414801250724989300278927805893629680906178963474029153634226296577;
G3[341]<=640'd926739631738550213174205397630189654168309257569231217194606992036862573565748907567051489618847763186833893270620599921989541266886160291193910677159460563102911652480120924353099969786365028;
G3[342]<=640'd2976166629467458079843318232497910576118059720128586562280621542848262220531816192037735164996429111798577518906845750140506568517794106869171664821214307693790796599069498016138881235088195623;
G3[343]<=640'd249464977447998684351052758546918699359342717623121420178406597249330777404084139307051101214232264094329064472647814231861513472176592504874268799400186538487867724683566533203906471327302957;
G3[344]<=640'd71279440983671708989163203195674406550454198235335965018233716339142827105544462266325666649720191055627017154942685015416968165508954178192295933303795089360179608165631905646684469732649038;
G3[345]<=640'd35639724740944130256869132715602438406057462986815841408571131061094578900223763031954210286567985776335275460650458625410826175727015366537413578213651782047122832581235005667870740813740816;
G3[346]<=640'd71283792066117530402503285885135964381785810699695215866221072604476298832133130614173778206302242547026063120398489367368893137817568293838627086397117097816667860524534251655131528075151686;
G3[347]<=640'd33651279004888329698218381625674460192366808070697736554220904886077460279143230898551547578187780372803928001342661672225009983592447937239155601961183773280044890262089935933343726399921746;
G3[348]<=640'd67041478191707876731845707186842223054994081660031694826911112681811630627360982154523055699420764728603139471644279907106133880545968643768592762208759858237936643826755534824036150519277383;
G3[349]<=640'd71166193865404462166329876988640379737873940138539744891683353506794610094648187786713879655191233187282102887813438003570581178574211705128819394646948583512408768595038689203314614981639505;
G3[350]<=640'd178220333175545311736286394272080041743266229346347775060443655435934189239989867892564132994271631949159322164725058682877897722495846948542745485400949945232096998797962925846569697211986780;
G3[351]<=640'd71288096422935635040444166389074914129622627809842971212633131216086031188489739822428453970354391226490752121700704382717096340031663401324175694642920485943871173299735250735265354058172745;
G3[352]<=640'd196042366836058773622648864419512176806783990671281627412855733045007866856197007893536689795203225883359479533569366067155719222827319681745266881758063026264512039984068368638986534984627474;
G3[353]<=640'd71288134384777819712030450380603577399793098737638377570595973298441290705858854856310451257733039331455631438008520550815994507756626010919951102181130019452192844748926304229278315050059406;
G3[354]<=640'd71288117649781514647668804808122684532400752788935302670863714179787346473892216802089070161936515049274869125301857171574809931592030480502415504376230523088652600283011395146509103414651659;
G3[355]<=640'd71288134650334137778657454970525584776473023383860521317853372292754229740613309421312055782255899032319773411063250503992960046797600449239903173364816521859624441322299169927413189512804993;
G3[356]<=640'd71288134650343507832892356304362275897385133601988884507896642716660955321896808392341220848031402554262788178673550526757711450649528031339871237586518751208261333099519102162626347286404610;
G3[357]<=640'd71288134650343634462348134033072695198706321996882153195416280338134218800457918679250993833372083368233816123688161731298801599993124201860684036907886696256390455463127025104948830922212128;
G3[358]<=640'd71288134650343760106456495612370671864195569938359215177239978160892102279556401847104065241528644206773234906745542364497574370783289753701945957663450491041658413495213149321194552460735921;
G3[359]<=640'd71288134650346800040072987793342755656076638315032954619148124083538735622489257262472884859280013220368788331124413614800642436878582115254511143859568264663021474132693295242751749884477696;
G3[360]<=640'd70931345890500093893220496600449357815648441525514189493637719088242091827002298085071912573926502246091533122389792288682041618475753829510985895401025894409553245604119379332108297154099200;
G3[361]<=640'd193447960901429092628318309658594446604597253750029233101236141941493695956745504306501933247232638704482436167407509357306202285465001332052596592639859512568520583296707874914717380506821641;
G3[362]<=640'd554715674789845581526123451172175114393945828432129554996405161886489075713511484758736622259979223501361621056421923815706735398544279240813551713700933882371077194152545938676087445524987648;
G3[363]<=640'd31188588653254322866387410640281399597629491456462521446241227572971888162684002035585712637114607094537590389659725270372960667686380361992971874327900601408985424702639359868117866722492680;
G3[364]<=640'd258419553437480267518200749298467468854697241668030895267970866839897584680007587393109390690539870245947896449671823020606709706293542926673604508124785962234888595072787895458248047659714572;
G3[365]<=640'd338619466039864124273130016109817891986162508336951123855135959216144421013848670893925327802405379072859607809143972212066981001798590736324380136678138971914054488490171637130773505366819340;
G3[366]<=640'd499034348691365009895280934711231503313702443014897029626671417072266306260492287079463632049441488590999599448368172526188654654275187570460772653635763989001862178315888253739124134271914018;
G3[367]<=640'd142576286954418571302138561579312821529821468572898790231391571170569710846343915023133163201659099697479101969872872307930874586599515494061605126554755606343891923902559352314435004507881568;
G3[368]<=640'd8526826473950867233960534416005637153767390109851011615235051743317578214640535170327810384198982419184546941880411106515063292166728235366992363206422348558154827537955664652464173224;
G3[369]<=640'd531300843061631497974444261755755270255821890889958657922715101777365801621981497476911386604735443218894861577635466130880042511418685126555548158447678831291417223402825476409925772;
G3[370]<=640'd464762197892187142823007955530456766278831820546215329500298193100713560086255711977474197253582983971437171123187598558436869996180257809161534273443209791781391544136535447262396576;
G3[371]<=640'd66392321938966852403975175368934541704013772568071430630608244217872310513003911674735358512629740880030718553997824626246659050195205350627517912536429442424194949110730002708824300;
G3[372]<=640'd62242738100041448652891096009496082698826816660132368437470658258201459969302151390314343484406189501115526540204214389103414222766653367015762346133206913031682054748562534410747912;
G3[373]<=640'd8558375889623703165594610584159609104842031944589967617368779783675046627671258368900299429803476804535531047046158763873822777731551354027665401728542697643640473938542853236064258;
G3[374]<=640'd3140502506481669842888628627503057488960640301524256215365128450355261630601445515639787628742618126357594789819917812940845973499620647371599224677666158135480499231310358733914124;
G3[375]<=640'd389238692625478844767987337327074816219204261875049091900130718144646465854792784592840624093254694169674894754690528041344611389792122467918708270947030700521778610053121926955008;
G3[376]<=640'd40019542941241796825060852900435620876294870767278627752083506369641411074148998542459739969150649191842330732287949323893692463327420366708400206555257254387173758440547878502405;
G3[377]<=640'd8100595259213249570771893833968173755217539443391894596438244113782689936008346388211115226458228081364014606630767454522592090005852726738026159999952876758608215030225665261576;
G3[378]<=640'd8104491890512505341773940075008431180896307255991306951859961531470446449828779267889869855205632397295835495064317372307691253326399317471244480831401402622361223524606772510720;
G3[379]<=640'd2223994850104913290802109145568664867824852588380607443684729227553319258979719174426475274464645820133425626788937464462911184265674342385540038258879950539379026207576472682496;
G3[380]<=640'd1821464556267055605436303995041616111866918434743752074986177800213890650654769940807000760700598069846856288987138065997685103592476523605855910362538164502942276455664459972608;
G3[381]<=640'd253235599730691743498971730638001902738519515088834041132474324909371767262152267661808015457189319081055577541637195669137707778445836683878621236584631227297309093473160265728;
G3[382]<=640'd57133088745352532673844106783585111817505157805456090352796181309172493282131429713681012087473276488920237670490726393674386856268199717206540009911742992055642793695556665344;
G3[383]<=640'd4822941704644599461036929724283335117166570206286411929560405510517435811941964369624106069403225810572316138820081878520517015019036986034535675954091147416088889277145939968;
G3[384]<=640'd7682700592511893175438537723492716751164179870971476260178566511825768440591211862331185281420599629744652322771505087315670343916625615837426575154127805552957839871630639104;
G3[385]<=640'd3208562470184392903783903725686838814254545065758831037211309958253338331315976859709827014898547767295646292895306250865479007007717191552617800065592489311517712386512388096;
G3[386]<=640'd757389089048910442786045294867758635833905383445300845058958624668069322918882659561728940199030778717673265025467738229376396533326401955093669214787503950146429785739362304;
G3[387]<=640'd193223103081022580496780241245319789854739702527253766538136702655235858028429267470879652948141453345274637575209477135757840245698659286404999584546418342987503134813716480;
G3[388]<=640'd46615982201399756607745501450558034649439314258343908708807351223350545567964021527328809344185925056577550985532041900292611411765007946106606391118118827777751196050128896;
G3[389]<=640'd24168455368553663301426449526016037205486595642910670908959082265420070012084717162926529721188651563461591553646838995834596604121202902873276812244813412504430398104666112;
G3[390]<=640'd243660616480677552557424261981559057228901483219873176751196313434447744201967352805285725009242614709211462868522145294590022789936617871808432511686992730284362374100250506983262356766720;
G3[391]<=640'd469916903212735257999798064054023455599795250129312590405375869322684436291132168604047256452439324521226351886286962443862771508587587838835843899147710447084289904481201914577160039825408;
G3[392]<=640'd452512573464115432034519556348422210881742960090186569390117023237109733048589783770780591337334703580478142451337388796693708213682515708933722992373609145130759205693046014607046333169664;
G3[393]<=640'd261064946229297364530943515302414239998556033412123151539101447851426995012658665075381505907956383890068278948382820001710651280255216977250612839919350557612594201918707566965660535750656;
G3[394]<=640'd52953410273277198886398791352328419946400183190438283073667198945323699453930673465872014370588314766190263151682376189410574267788045767106274627982136872614849029341184;
G3[395]<=640'd14860178599072814191473373993085029054649588582035265300219272090140679359770571065406896299154749216710014267571874969384934790152218839711777513250287143355779433627648;
G3[396]<=640'd7544239683855775337795377917806896496380455681270550169254428821158286307262379207902893122844111644282356234412453811055266780310660454577182400388685037134720746389504;
G3[397]<=640'd2889022485830434681119458654133688238475058920286748788686656009413802924274152040122423547482115525659480038764975060420827781106471789942117767190612186253574784679936;
G3[398]<=640'd711303239888837388522913694981354872928298262681108167181448019332685061309419666763810723865390529711055247357931190845913871779340423973015809472942901474177398603776;
G3[399]<=640'd29944770216479456229327313172476119009841252804723261719058570341808774383371488628000972536953389749848249207920366540520890227602216821006775377771346843051495522304;
G3[400]<=640'd14742968619450782166232813614510460105444165883233326108168898056383576836015011298456688360453583435022974219885734947424758859620755875931667361111620422570965204992;
G3[401]<=640'd4376544217596750645509148658284628571040223448411471599732506522148417397051114813172928637663470691943213741683937568824838036344752131819928438532198569724004532224;
G3[402]<=640'd4603288594576598948065190960868928083280166674126938165631889236309399486514709953402070572391878988496585705599314875314760164751652734125516518257533146055187628032;
G3[403]<=640'd978960127023453462785620045920126369142027252992703484265753436245087207682680638315398792353970582470519940094704304481368362779578198484471207837516331568179707904;
G3[404]<=640'd233943517316246199119856158129874941879306640763185459565591943469947575157820053153404900050864792760358924104499360176722707602907755744769182618175345054957174784;
G3[405]<=640'd439347050248355906107363437128190273553454147162376012631129013466754662613927236408761422758269768677039827440363463183614761035254661163160980961300465057792;
G3[406]<=640'd21594789538943760409946711874170503507600229169405946831490779314522931560602594898598986502043739673691035576978538172741176359764589300499356820335612267627282432;
G3[407]<=640'd13496741383655776295147015549762203597613146064612363998752926907663625153374111217022722563891915397904195821935314799153816748204572472910220654731205889931345920;
G3[408]<=640'd3592101482840595334357322074606400322668447918488516356167429257486150762510527470311050388566648172458698785229038965179247222391630901673740746430579002958675968;
G3[409]<=640'd731066841314349010841399535193939640803215803175671342896074412000774197781991736778354701700383704349908833536851352419420008293347002601007274585146336749813760;
G3[410]<=640'd175738820073130910476197143470589628279676642272197411269036041146315715817759909741845927894511418902027637222673034305040003698658718630039866535784274257248256;
G3[411]<=640'd28123252944483557338824062499965576239726203107809105634136904145592941675353680214738956062691352889046325857358889874624273115686583733171619518312043562139648;
G3[412]<=640'd7029552856347994074527370401756090397946322094774531504102720878462084891672634129440632025000758038127639344399432100681824212566436504457676819071969982939136;
G3[413]<=640'd1839765772915402987429677045029654876682615131026793874009511024348580554627769485879876361190862232202804158428492653771780974552811458847363720151645120626688;
G3[414]<=640'd1646746975888570173312338604520828307354603096455321629424306630563379214967606806078615443285402822633782108104629852708827736424777737375359224406837819342848;
G3[415]<=640'd233403120444440730309381173442670942288340938638863677673810018388111123949081460168103330771757656189754284665957589129135231900054007378188401621975292706816;
G3[416]<=640'd55133224033693294838227895393028010912096256043708413640304867500214022391359976852609843413665430330737061120513358423119323770645254156227791471084922994688;
G3[417]<=640'd13729595326654560461011682143055148355095464330907537366817450959589666964400825960457227203379131911077080840044954161435114095864038934558093978111796314112;
G3[418]<=640'd5148598245097963216682221373110197253083293600833743459671966370117169486391185028582758415215960318303174090103591166260925237384912904371218311063611113472;
G3[419]<=640'd1715361427236810729233114200184566611333605641927359285187156185443641111606692317489511189882079264041606344346863342672730503990665982499917893423431942144;
G3[420]<=640'd858099688333327704932091237594649562170232497843844381224021211989291285185416061149456135623613902410275213445584777680315717226166441367674123051843190784;
G3[421]<=640'd107942932198943295772013626627130543668690231930582013315689936161326648298458060278350396587994791498556493699443669757881873785864105361673786977301823488;
G3[422]<=640'd80446847581996894010182276105173899509887951880157537107433901714973497119759623286086184156982474075603083324142255559138751371573739479433049787718434816;
G3[423]<=640'd6703903964972084304444329394137907865697011498020617277819589604705314099405126823175488774276326353707547525115231375436848561970281546235407480372854784;
G3[424]<=640'd1728396392948460652065717806898792129680038280041597752106748871295865513669300534814567660446543886296580115629909282906053924698204102920207653671010304;
G3[425]<=640'd782441860459485550617200370085792246483628056346420134024556384480743668709614161409800510575070584452099094067084246948499606683323089775011345599561728;
G3[426]<=640'd207973785551038058991494870959355599831302692244447733711452202561756660910121408093123629659807578366597920892677335704442220137507340238086739259817984;
G3[427]<=640'd78561374589507410351481481445251920876562635794157582087602829633157702695156188093285810309266139262620745038018674075336555016179099005558875549073408;
G3[428]<=640'd13093562431590475225203833485405224456977822722170167466002176991837940223870527359136585929606608120951561030915981531172763869553153531947123115819008;
G3[429]<=640'd3273402905925811461525605073040036832229515106338536067968276141856064033373746252085375262473473416200934628328173352653341958408567743169008848863232;
G3[430]<=640'd613673329973483650209606482774273721675974295881081398296416767453812513205115704551655605498484359657287215211422166281256901285552339616714897489920;
G3[431]<=640'd409148851998615217169591313905261832330168018460958835367663961895676667274919611673007775975904343995500932976849925349353571761218345308513284128768;
G3[432]<=640'd51146728248377943552135045267726611194459673367514770261073588651859569801663771000565699584917650656302394472707181635687147848685206816637644177408;
G3[433]<=640'd38360046186329427295178128340773782251481344631336138134705937385206582689459611784450425328090818803417482477962405950807559911382504835453542203392;
G3[434]<=640'd9590014429177527664255916412636661806565107297923344643655704543488786608243785674058806011189852227760407814008994936287031473043269595157124612096;
G3[435]<=640'd624739928620358526779277573156337513077547430458550740652843786757894518385743111066750794362897597584988149477604579975591982691134322706334351360;
G3[436]<=640'd399582348342778332455754676126389886903675427395692094269510996232265902141208785169789962044512404078753241197437445938301678555910476806462898176;
G3[437]<=640'd49935782474920325158732071436355059122548416680105648572168864907880081938239319590568352059953920679958053577725703953425035847584055251104169984;
G3[438]<=640'd19462151118739661248309895708247556465518132771345689047008424633928323007594325128010440329281432997148301864402308121025453604007356792538398720;
G3[439]<=640'd3121801580462928607885077351021721150607061274572269405863020863054012237966910193571005355611083999539502318129786245757335540684696689703911424;
G3[440]<=640'd802539359748163327689260311423863158027175169711592391627806715538873655278765110137867486434833977061674703217257531869914482162255742684364800;
G3[441]<=640'd597522020647046145821940361716565272447981866829427749954574293999208878980252147350533353995482147746593728634374748007871963359490300700524544;
G3[442]<=640'd158502476519416262053257214082897353471078631969679749878524130565705230111084879399223990866355016253042408111935525227699400593883614796578816;
G3[443]<=640'd46871956993269902888175837312568294062930229175698201524734364148601087326091243404081695017424015789948572451228441204565482102791982901362688;
G3[444]<=640'd575668152613507949414316044720823822139937812281238562058134798686150309005434096918067140792954997073510400;
G3[445]<=640'd165131900351285148835979104461750259737352679220116240909106396435912892257078256335195475761118132345765888;
G3[446]<=640'd98001321673230277477451886940349244899328;
G3[447]<=640'd11062536532739110488009448639031640719871705088;
G3[448]<=640'd42307582002575910332922579714097346549017899709713998034217522987550501117627444157351697997348884993457647787383615060443136;
G3[449]<=640'd19283256531108031685905520106503187384513945383307316658438144;
G3[450]<=640'd380768238023183192996303217426876118941199950765270496889376095317801144174553956024494079992962351879270972632155196269527040;
G3[451]<=640'd1057689550064397758323064492852433663725459148756203305229863589212498879646883676780226009579936926179414595656755153702223872;
G3[452]<=640'd5546354770209691541004818510199305743190050580588329896987666356028128760293375879179037602135581912792334678361185695975673430016;
G3[453]<=640'd83180090823624445787352425524292511103093112261640259454036872231629305081571782956297913362044668534862432343562883328876474269696;
G3[454]<=640'd1402970865225132318946677577176400353938837160140895671129614992565268876491007300892118608916612028421939449460596041762134546186240;
G3[455]<=640'd1070250501930634535797267875079230309526464711097493624448968042441444083337755136006831519620677963538782382338307619454349454868480;
G3[456]<=640'd1219974665413158538214502241022956829512602711088837038928004224658959634486458063495704777936150632168794167025186123707634002427904;
G3[457]<=640'd1064705162542392907155527584215794212024557387286894654737403922334565790178571939293621698537778938553211662670703779607967512395776;
G3[458]<=640'd1395778701641990866386072804758435186649679595635142245072070185403338381176021713097924407841191235977602865823744;
G3[459]<=640'd214524926879081553593184399971293538039670478706071266883623250925010598655258237155382526285694039142163389877502076510688686582322843141964855148516737024;
G3[460]<=640'd80695308690215893426747474125094121072803306474696036089420079018466738189925612158059773535543835077331096756476182528;
G3[461]<=640'd1716199415032652470425315005777629835977783264565558370323826052049952644631219512006228833730116955053100286462387739118017864391423477517504773370553565184;
G3[462]<=640'd1716199415032652470425315005777629835977783264565570984566213997443266504146849636194602911733567140092564497981158150485253760812987134900390890515755696896;
G3[463]<=640'd65496891123725728121826229445925609628091459263756273002009235179992668192975383308999259342957664686854211027901051591182375130774535929856;
G3[464]<=640'd339392981277487863901329194950510354511573079374880173308919576323087284342297930865723938631813177784100747931040120097024002039536020357120;
G3[465]<=640'd224945689727159819140526925384299092943485239871677629023628611593455036142505377466086948665598580264318402403056445517839681610066962320580169032978702610202624;
G3[466]<=640'd1651281319149134800346780053861062781479533630301536112715191682996610221063765763447006003968665462738814014845777660400623436593511611610159856116252391189321049178112;
G3[467]<=640'd3864139372759631413057977753218770873889721541916190777173327378333147255993816818434414541500779978312871251351463669481185685161985359311002104320827371579203742750212096;
G3[468]<=640'd1913378901959530117815133546959568265000980558321701472704871941919668852843206179338702608568225292789300491372639460528863957349746577682571910836140829321298747741285363220480;
G3[469]<=640'd3939602299666928636150625149954920152238291268578738450048322552819728049422934582433546539571322914737882246610632577898775409714381323153573355542615759575628294034556943597568;
G3[470]<=640'd15829144045001524653361491407109890942897037631523905776740130442954586989540084220486652497577376729212770939578019621395916541187456351813746314449417082766060819911605747712;
G3[471]<=640'd31658291386907884434534552357652578632842525085376274317999933824659231673730204002768985549085651482316779909759185205964255690088631312669673213666363826272153245796930360970752;
G3[472]<=640'd2263398275169258487092172797364911742431599947187545896029356742903170185581671078580786622227112604302437682492675137032077317277667233984563710735144467008576617756316513869840987190565799936;
G3[473]<=640'd4553529601619897275850267158164175404359575238086240971849579403808305581562424344462208303691390627882151265105458088642596798145573595136789841342958930633308892338793455856311755853159989248;
G3[474]<=640'd4544618838117437112529171454213578855932330062482169547963159699409196979681712397062440329627247352418471288819081214293449947359873158275609424620308749591417412018147782656444444316643885056;
G3[475]<=640'd4562440345430571962138054172514418598350069414680478102465712188963951028974607102312319037999427748770961265882982724019420796479002673305267906874977270928094784372557602142373118666189307904;
G3[476]<=640'd4558542047517832474260735488533852903879377797484811763920043113853450031751861116508698214504297731808898835304104489853700873138829542162905723470650960049793538823672237648601947604586070016;
G3[477]<=640'd285083176120547359810464812557766899017941406342003020607259106537660034422762627333091796610828604793841183653007400460231803232571391042545068817666654453355077902006545705021610019853959180;
G3[478]<=640'd141967117501994982305147074331156634102946390497545076151946076353466646350699117098736675190297514400708036225255127281452690638905520474762829346407226883460917077204260984762469059356393483;
G3[479]<=640'd570305072696287030467030149544274941217903985106871080018058530917686698836791191858355398504076280700682226229009759424848749122053695298129194510133749980939558916898276353669999985770629632;
G4[0]<=640'd10421331101413813803596711331166825599489479307835814714861895713002890260109422257172279819960802706900034613129770465881837764607;
G4[1]<=640'd5689498613970241458896523958356275450623094300856173766079306130438018304114199615536995419568004011301259593956463594783005287186175;
G4[2]<=640'd8519018875525491819044984452552568333857550074952716703340668679476291434057964833270190735252682708050575030899011000943297699577087;
G4[3]<=640'd897192232679394129379940783054231956470636747636656473208040626701630583430445506751910328921780382533779592537475850239209239950031103;
G4[4]<=640'd897191588212624873361807847245006761852698659066916035595632350660663166727795709689316709607155613834764463357063978048399906961556511;
G4[5]<=640'd8517660338758791174041520278721313155958910831480454081619331344799522851575977742527775536935452110465623400474219588812595464832799;
G4[6]<=640'd5678446656594251311025234864169772746472099173089781741059833211505526614248275394844029080062083412753356723227550150330157891618783;
G4[7]<=640'd112472844863579909570263462692149565626502124196680288379808915104014456885178936358163550718014629382863611741809548216426483879235421094579557281307439728095484;
G4[8]<=640'd19875568780005286327789819845237159855857777572457261163798119221708914048404947174636500833792008776254163748098387255279490523806783;
G4[9]<=640'd2840253686845796746226799192072993702451076754770233141357070411408104683750020033866792842711781784112767733379346350301046355605567;
G4[10]<=640'd139121482864854893833005534005598992060877995902078131581451700631366487922613000071878320835075405355334734988921397198330454771564671;
G4[11]<=640'd136282269098055165719377866054843306182046777790271598426031046403698384719061460478951659836055647110618565164385991185382700742672739;
G4[12]<=640'd340695593290091502047727835756147379169375558041405677224095118853581695630577735935114285257500027551432616262532094558691;
G4[13]<=640'd583265691212880477688530742976180307114222295955300860960625182158618781623054004836971144172151133280047538776658927419427;
G4[14]<=640'd363419383893735330606559209959822594363060096279097972758741013261377208079112497981791819188148025088287170958070638435792368496017443;
G4[15]<=640'd741991204453505347020035855568301662764170928814938818904983470010204212503387910018700392900343534013449147058707247038811668511241092681806362357127236036368261861859395635;
G4[16]<=640'd17822033662586700072817076584766790447054814380439422180230060330815675613941106438145155079102149781366412990435675186245913501083742706593641494775911372185533492479985548758944192013994112;
G4[17]<=640'd17822033662586700072817076584788290993326343448505870469730906679853708377534613601450947257418319779114962418508944811163249522356184258637241967456174841551933864111851828569390628336568320;
G4[18]<=640'd57607624575615083292041076139287019460227858594525444645808495902062040262644458596262499226672734223577376012527754420084216875845569083486492843561403931896579840;
G4[19]<=640'd1817847433583843407427341811703964634031992846986580797565714117635941886924518727065731912430010302474567270781326330431047398830298498138704747190699331519720845347349782931594638359529588494;
G4[20]<=640'd1817847467576674947700438014761236165874308788125105997578251633755940347372309477444100122821599986506592539634985643968277660810448817397789892257176596254885863479034870665316475981075055374;
G4[21]<=640'd106932201975520200436964729888659340229124844999661420074577780703685780365873888206598724457031339691329057302693656945379288212955181256467414669256175347295333074117178118793474640006086912;
G4[22]<=640'd2423866331402111850292659121768291416954879754873609701292733046031037797138598778787643206637676749651432181276670716161312849646550277893697394066947232159551975365076545405307205227733286912;
G4[23]<=640'd2709158107828316220218989128928139830622169758468468652963572859968957088933765537637023946270253353354107643900475319272291276614336755961864962846258961294278698701207256830939295525143363776;
G4[24]<=640'd216057349499382905895762773830269598839286565773390994278586285722975572687153168994956859669918611056646215587036824416476952442312605770310199760312729221969262017687276293782636119430529027;
G4[25]<=640'd4435493436435778453063730094981223730290508775805705302078306528766243644310899617695238661653284780696224898579929086762225657023957537801101345524754888187613685609998172558998159482414956545;
G4[26]<=640'd4504595152161454919582996440443124594507878524695965860660876170924272585548250608039143656497054705822579857068009948213755458728609692536290479750416596003787455639505851321498682298816528416;
G4[27]<=640'd3698572359467029294103792421851631630399595756888883919649033951185170850191208946863185799459503332874337730870795901171704849843700909683167496635642088190543983700988212494050070939803058176;
G4[28]<=640'd2407941506184605137340167302741040222082903040941310518444562321919961390353625681410099576397182167138451421824688836595985666946442936616352136006908706542476428568923496418385286776294998017;
G4[29]<=640'd3439148044055906765861434160232094348277221804132450676008916833627612601396541032587764246613555245673066062060828281315398053121216407264576626732023771985041934550359685307406707920251912193;
G4[30]<=640'd4507899255387169410482723885826790067063768234499038515922947394394753240619866991535968464681854448898854256909735092414967854127480155714548411049728263923203199774619522261758201704650637313;
G4[31]<=640'd548274729933485730669341054163530196841695809919408188078958484552768763836146283952071830513488542596123536207267137846584998629226733956568045206388675447384742260870401646659163695968419969;
G4[32]<=640'd1121681074630087424856190152248791720050434431556126095465533483953928801111116829977470311990030812544944890558436892874030404667899941291675264699831978152941386249280591700976190786262532096;
G4[33]<=640'd1072914170281056090366764770392284944816445341810818174338293734764737109998927493055135210955038728027889800082649936123767290336788617638707785482884696468975897839286113363429847147032346624;
G4[34]<=640'd3476400074031545523998620987239627422017673248339503037102213895479810257110939812098707214469179481658828629626209211474382959246906155251485983026000789233678692142814556111693494124122472448;
G4[35]<=640'd14254657024675411441544508464015423202205692292838236736859410953091313351113636088686383044673908855040976220791189364952546652354417851642962213260469925846854611852349052407145558521675776;
G4[36]<=640'd1085806035223622020202281947073992235070229173900398701079724114223302168395454827203222976120486664992525543484668199908121048450783718947711571222754716437164729998619729484703050908670361600;
G4[37]<=640'd1087032845057766078655222703969381609255059243130387149520206179161671694378658289933328936834811880421374363795674429750214824272984569897294154192478229296323051083855448469803864960043843584;
G4[38]<=640'd4553494520182737231407602915217689183525608374770263302162387196757335853592241258979971201411822157822705179426540441674481818800759780061542937183563996972112851714896094018925897990872760320;
G4[39]<=640'd4552693917632648903704544652736997502551134326352204382799634751643180869778168796136343815214611806951128277320674351588534236091505397410596156484179429001076293687924233784569617326603763712;
G4[40]<=640'd4553494648724089610927321786449779744620520941425775595598444900700119581866248262508644099307355327283817250428050070355566657691522767307862530394371319684422548159506860622455091256155439360;
G4[41]<=640'd4553525045749400714225684209020192334555103099318895019906085171848583354436273407121464416212011671220842904058816076339332176605860490279946424001963957988750872178357144490514241191220871168;
G4[42]<=640'd4553522666253267652893522576144283194361526124913541462601605715438830061551657174714204104939292880764524621698118940672589964923972366038602769497036481350304376366549189142616520667472855040;
G4[43]<=640'd4562434090994389970638180971533479442799636371199261028528066965895783412984538102400756141683026831629790343265738746924542179171691173147795233597994542058124431247424964383743635920420601856;
G4[44]<=640'd4562434086749435543672926118466117455722964923665761779284982323819643984153701652906050059068666210015066696779868810387374083793331705230829513397669033686494250050337634592488069220731453440;
G4[45]<=640'd4562399146367716022149523145532964292100651932480566562074292660931322224845798700363474457588692604549816948341587282580449296319333941622152717756499364742930892942707621467007793322436624384;
G4[46]<=640'd4562405808962697978992589997866374291538536884954658526903350985614132166024817826311556754097457438744099271193407076740863955932754204617220114464061781582168185856177494359563643265715535872;
G4[47]<=640'd4562405808962697978992561693119395081693372626800248142343539356755471008298632243740121784215150752535412367194431981802890309275960561248120861432557263237219816772931477787392411982465400832;
G4[48]<=640'd4537514346939980861014636006475301849436830685794159317502047299591683186321149847720109952763976423228116867881544857554928274195932365430698557123661848297665572528886773976279019345862983680;
G4[49]<=640'd4562402409679543951682918737887876187858160745888624622955106891302841322837463361485469822119185405707097336817022982594203975880384420747308750652273745852329838203504945104077017562977665025;
G4[50]<=640'd4562403497446003661536473084091250079966921694958768964673735140133123787799831420662579000960953833761525576019460774873029026082656068360833281762858175460393882747047907242593066796602884096;
G4[51]<=640'd4562405808958548463423710891888961821600713093973404710046028872529313914696602045945182138604282797903250171448166057638248936921597127422940430830607678181943226599987945686461760290160640128;
G4[52]<=640'd4562440616559919233007607216621603866611771752247527723617322335079602538743986393714968031457849568914661848975565856906620122923749751496734421937778096379426261308677833777003460190571331712;
G4[53]<=640'd4562440614435367261740327479967573506931873283774696178242092688639743397109378400859497650452214272398535421621752564021759104673593649700531279266436893757578034406532868684577756161253572608;
G4[54]<=640'd4562439528789309944268373512741326442046051175479423480010248170130307111825372255414536003815040936509920947102729621889703905869099618093299283456666632809318307427994744963191217138643763200;
G4[55]<=640'd4562439495858746285106368880873099869247167493355812558096161682235633151431879937642239424565669023669997992525753407246537895200034218633324121757447788780931753349109976645268826883918659584;
G4[56]<=640'd4562403633421479401390875344474926883612204652154501859214141185021710129332388318057138013399639940409245818045011939870839541175915704149406857968712864934308316046760125743888296547092267008;
G4[57]<=640'd4562440617622195218517479987197951166697624347708319351768361621277298461924054309625141838816674138378733321303144645700715711365442209788871854125370560851876707893425829953296501072797368320;
G4[58]<=640'd4562440617622195218640205470398138263203403504968352370311341231113217368242651445753143148160625475149609047373222593178174814950142054964855056756727559972911638523019875139530846901547040772;
G4[59]<=640'd4562438985966281285531315758793677419004301031594534688569685204357312058646157473825450155436507726294113407513902253504325511689695956368754516580559508774357398825566146557013303097320013828;
G4[60]<=640'd4562440073736890574270685091288539848984700063936789220475912438799756476792398481490351804549560245495456802712563726212659592952601757920669828780722154053139709712643066950130598391450697729;
G4[61]<=640'd4562440616559919233007629860367471738597524542213054901654108795021853340178978275811706290712928060440753489845447225040149217206722908387581032485137973825724623070043086488596133304082628609;
G4[62]<=640'd4562440344617266910822037510286051935679570290916125617006239612749219682764603995980662695186725646845536855590800722787951944076806360553985339910069396849261698170791743918369326340539154432;
G4[63]<=640'd4562435991410277784408424757166463278772081006342328619155119626040472957378149957844041903001204831530777831978085632178664187744918362797471152219983072119321246500280507627098056561820434432;
G4[64]<=640'd4562440344617266910822826376234675989039276743935727121716824666365802675806451833894693255198095449807696031193520100995570704591699725744673839974859426610265321713923833284810797737148678144;
G4[65]<=640'd4562440617622195218641115931519702308747156833245033847315202872518694895453406442914731260824047309680861977763017963944861558364974835296143832872718261801978877333153778589336941838129430528;
G4[66]<=640'd4562440617622195218640673331230994947078198305216223429368604787367230978996349043099328035485895895787078647271575997772903080637595590509203915802965700995620864024520674538746567404441042944;
G4[67]<=640'd4562370864331874578220959235840101066874550711095284419176428316394042917908787015456235491836754272819009090948157718879160218588494843183825278103005516331364804862550060403522443503646801920;
G4[68]<=640'd4562440481650869057547885038202936559126514654590565395706997599374049495077591261849517639268070688695217050281739665071236486953360554902885113012409300383273045909355447119265041043154796576;
G4[69]<=640'd4562440617622187114118146794197980940644817015450381387136692741314153909770749547208481857911291903447104759444421214828291994815754046191502140096461299345289428536190762717839342967099228160;
G4[70]<=640'd4562439801794238252086712668374606765125307376200691753829374703028319925030138414342113642548761764274060206798863189131168137286550936164619912993498154080695909010203758477907107696953262080;
G4[71]<=640'd2253651033599050095658462413916277544622581050584695412848374732252271720447904350561069816685874496822471899770594016258298654352575526629077010298646570356409531228016559377800838261686403204;
G4[72]<=640'd4562439971293650209613313296716423494022584363308356431627530639956353373668786028876232757481339259525229124145477381994924769396743423974187829527729664936429222315340368843355265439589466112;
G4[73]<=640'd4562439682819327861116557606366435212953007745085980185125970946434131203822014483580304638058493263487597594550032553697060387697752023706051926698861485508867607550693714220390133192043003904;
G4[74]<=640'd4544600775433847365172680663396170127047863463219753130256947394239081974618598102615248599273720285692940487190387374560754425096901142338206676453496133028540830915909519365940855993729548288;
G4[75]<=640'd4544601053733557538708874431962708775350873387240168075573430443535087821420419889878554304037126759314671755619263028518851275450287425557741793650562235326881297052454983062939375433079062528;
G4[76]<=640'd4562440513992193401400113594648971288066817220903290295736839500093868061610022774900812140172179720847463902946834301903697835502673108037016029623676863076093111752478282442314898935709171712;
G4[77]<=640'd4562440548516162934469673450353167140073204555567080105218765865549361978221894573911921705475676122313824822012750463808180481777807149933580319692651125628074354133255079133613291994951450624;
G4[78]<=640'd4560212795428708800527520283922465055675840831263957993107839499098716658863826276115696781211657318936713606303852692448257105279262197359268929364961228338755366372786162457654252799227068416;
G4[79]<=640'd4560212829421540340856564507010621416528702090179209581883086601103376425490372204910091843232848224349414297125089502823911865505918351639974620375064567476820550546740905462095342983408779264;
G4[80]<=640'd4562436529453064507981522096741413316129145556871607970352413534022231484430622927355529707945811872679704582140538032580210568311624212190499280550615618354053957588481192981632026105528451072;
G4[81]<=640'd1140610154405548804605815753822774321150750535988360042282156390357206053849633860713455717340683032556755597287531815076160233633555129605174327097183926538813128390095841337316460329053454336;
G4[82]<=640'd4562440481251737496837818358046205598770146057541489439131682090367452612380107503741251749123273235948461547798963843793815238426329710269301664124327442807823791413596525513884442021542756352;
G4[83]<=640'd4553528648575889149897049805584226318819194643197103772596229290136924330628119133433156260800054176329187867298364364599575375311847658859880780796871334694013780089199658553168316553056223232;
G4[84]<=640'd4562405672700905723934055057533815259434155521413124376758714499778545804841818400203809532927252189614251538160092025809369739956780512749238944233602075116887593333482949472563249887873859584;
G4[85]<=640'd4562440617072384405704723687773236352894831704716917203368198533082974454093464904852980527235727600048133589304777442784002812238966172424071636236182296720893077588566105753505976328503951360;
G4[86]<=640'd4562439801794238252056115315578080899023151481683196100276207278050154518466585490753422310871326416908582575888312518475584165509420013068630315388858500608691342344072228907111750681634013184;
G4[87]<=640'd4553477251759788083242953193695071247858654754653975578883792422930001910332005698154553371469047805292485648305649895422245813467083649406504567531222033875990787463543967575574137399425368064;
G4[88]<=640'd2798058873858913221905184521181113048903238911568279146560962110139106089393519028825832172971109418191462601002720243998715169237783744763348822543229467977950518304885003332496038721426030592;
G4[89]<=640'd2849819731954779671100512488377875082410030526240605723013366844713779545776890100810761489702057540304595959765911351852789115115962906666550385205500889784202293607987201580213014610566971392;
G4[90]<=640'd4559098956566732614387396129929684118097131371980150261683453667977128731436743779929267229961639325759119821703932895719248051857303622216275147502759193654600255337033625086454416882926616576;
G4[91]<=640'd4562440141523376907260413895410549243914311545769567482527518173091876049516413575698209611877151922196392369646791985507562770092667223491727445867027400225138061394847898263276552588177178624;
G4[92]<=640'd4491117469226693638960351149109588925630363325473205947095156911278637879482926570658390981857608722438544614105752334892864966711185343503687351272508638637653365958877571936978154674391613440;
G4[93]<=640'd2138609196326937235949852192854939305318862581871024567039793357264248670014234391557648522182639579519249497577799374009320895564045502209643931217825119083328476248118931386414240907070013440;
G4[94]<=640'd4125522051130753803479234453640085662991088192200998848055899519433655862312113964752517410290109940345240567192912510096733215664607436377115971967793473949066723287730726036834531142960939008;
G4[95]<=640'd4393131025868371179728936221154845370124702353391142066076897408292574451008415808944003767531408550493659045474179088497108732786617130746460944616843431475799426151274218538923364680873279488;
G4[96]<=640'd3970971590356781464693701043149532634436083598262228920629455242754222221594299989868131474199767165479765390995632271863466335839416002432687189294121994261704575831915532621255481993598074880;
G4[97]<=640'd4558542047758504377984785660829977688345982085741203224426371875700827229093904409001536547600464650827695350623686052763968390284403235620852230244780358690110969574929879810354803774855315456;
G4[98]<=640'd4562440413665205974019184621142503058193302821357388813019194326458213559744376281773772910769147685037338823045571920413400754939937443518105306909577081701701406232793239065191900127420219392;
G4[99]<=640'd4134711707741619793091823865486632074458191831053544227229185504791184211545523582323117172064872518753470505219633026667155850838420979773740672474637815111729385344982028223871561174538518528;
G4[100]<=640'd4133597898623371206149097461884576632923627510031812597519415198270839682976708901829466949167070969472691746847340650178749062873287531891044065770691171157037880486900217191516082391744512000;
G4[101]<=640'd2262284398044599238543564124818627926726723119738033051217332714924839296585326297613929208398461211646869101416349534817914857028005513058830477348455052086069928702544542668672867121806442496;
G4[102]<=640'd4562440617622195216933053538967444955132362858152807974627709269666284046964332300908282738701128082933802197457999239690474770224754749233316668393453603806929663045072471214363445098274881536;
G4[103]<=640'd4553107409823171609800925158123567459879308792517145189868408090518384886612637235905527452484950767816691740432676419139654946038124496240263514692175238596730338601903190248595633875231703040;
G4[104]<=640'd4559097898539844809754648355724594492254694309776111488948093753513228499731256989445469767364754932945411469945536099775454641547325441722935434371242832608827848013936343461455379503238873088;
G4[105]<=640'd4562440039744058978720258381857835506662018142803181241483402127025405512654525185009803917028327789243082645772842429418593777162461557610044959848481249172765315239179869529416041741573685248;
G4[106]<=640'd4562440345679541780672218301591622011564509496913926511306997987584557115953656648542065092843217402930800770848020996241583834370206962417253932967076072198711369779534459327167690907681030144;
G4[107]<=640'd4562414511127571180911172545893551663334236484614447516180835481745210914790826925460676006601532131595057519577185866455101544265257758806797509002851637843201535775437160265587745695801016320;
G4[108]<=640'd4561883543098904992064324145835287702133227232209654051187752565540155574670424179580903726720094840059606582527156732511888481762036777238550370429186670318737474004445560530456491661976403968;
G4[109]<=640'd4553528377048966323847046472582926694747533786200229191483520143595584401704982084799163359316955866155950786449031864689090377966769309413395989752378033336179335112258377312662293533310320640;
G4[110]<=640'd4562440617091053965022328453394716594999495552503342806185238967268099196000379108109787633431385691176980610632106354739914274481675212181097590225199935700629564618569163344597269544217608192;
G4[111]<=640'd4562440617423014957266506858174516670580133203194043355249135203393924237550523814303358200556725296470606284567212393737763955731668071322212946520891149785150982833495495025040804334529937408;
G4[112]<=640'd4562440475277212637230397354492401118276999556156391272899995438809252428879728692557677769871508407490594092836817876764780485404487726282722580597941416047451426010589891049114406337698594816;
G4[113]<=640'd4562440616559918726474988400257175715893530324198142649562097816059764691053174594168724986152081921031466216444801635249737661592242391102388144484122423260176746413901918996604997081831047168;
G4[114]<=640'd4562440565554072847755674755886579746508346833335054623621017265177093397851709553852515092526901449403224647105203658616463067334557289594822267323612799451404405042831230388019847646146527232;
G4[115]<=640'd4562440565570667870837159581911759661751073738126525320864329869942545649074377847272336384815823775474755593586043979411511659360797094516691155693305712353330699310322092272477286696841379840;
G4[116]<=640'd4544618580772776509410321569581581392017644172596565906946196065009228810367481100485767678689776905741633158053621882201827298516519182457795714318805449274062834173455051483704229390085783552;
G4[117]<=640'd4562440474015756358546470033874591509113217892451176439415789799036458349348303697893950743675274920780240877242516971982685259094324729058313232254101290573822792682793787133659311005933502464;
G4[118]<=640'd4544618347138451919131027137152034779306529738980170422150945921648284038555974767468256592265191529615157156027705373221269785358004830138633974487269257041682105889248223017562460903031439360;
G4[119]<=640'd4562439531179426859682879584309306236098265382996052708542967538567765982976859239276642486536328955486212575071749094001858906778855528283783220877833207692817706953786877060690936223450005504;
G4[120]<=640'd4562440175779699014046812079420128790173052247916580121301381565995780315125411127517643923225654818898661386892187133995403287170607101666644649547005947547566439255431590929883350675514490880;
G4[121]<=640'd2263362922632747593500527085114093833775519039206755308989368111657483690262548560478640589559598614606759898798076296459118029888304395602580706141775241943607209394975713943220212351856541696;
G4[122]<=640'd4553529056934637260176313730102607762878536248707475812852084141605370770497007255861253212058945686814684009253396885054294589582748533562982945786167475802236330496364378402402019549635150336;
G4[123]<=640'd2272305756758512090910822745569339218101352324022036710324692183139144045153402205280673369514487645681998656105438395827615760695919984384853782570373437325671098676759580175075279634364907520;
G4[124]<=640'd3546517121138839303265849175957097991536299401739342684103188902660990191944716758268349938140522077850952831568343403634668984714898629849666181528239176368732471512360149862011537556190019584;
G4[125]<=640'd1122666052497345478352101327868776096331840336156913930240227307666701204141571109407013724415674963778236361373351970165397307892721982794060934917503086156158790526085813388388497535062245376;
G4[126]<=640'd2280974506658676415151613032771324381273608565422366459543328622424695759338802971854538722658731163525658245837396394227564442132935453542598196360781546823548280758513341273957241270462054400;
G4[127]<=640'd4311820206866598844675702821626503636393533277811716412570134883604707516631879146153117901819303511254810402005677443186866216073585954366848949737158945560665469076758810917980917985971017728;
G4[128]<=640'd1005136042458255665946159887784204242288404538022804298696137358390730281192622608567180669712596465752286393788971136378865796430625421001533810693677876404959678323640222384068932569877454848;
G4[129]<=640'd4045603511281399723429107575686769664331369597312838205332036474725950230060401476041889311007120772826280550544565297612077469749564314143519793038555924134739687469308195701287967573797773312;
G4[130]<=640'd3421856705738149601418856461534980606581562073137744930760661079705430555841083651868461176440577898714605981365166863674293459614050502630747322459858167277191489384719158305511780162885132416;
G4[131]<=640'd102000926483082155158930838779477088751273691944642846417569568920094957100171739856353618322262759054586989742946500939869708241990013758261141466172406502792756367674483854606361174144;
G4[132]<=640'd17822035789196776863056003088660158586355922845658295273373186439294714519348303858389039340511319837832292815644894833057870981206881639163974749592370923084458815278588697136016590087651328;
G4[133]<=640'd2027256329121287071214445897228575223308807596857807370048912039134674739479193723376496498272993123470323601879591173049717197230986530025285126490015073890794835910215403174539212735832395784;
G4[134]<=640'd2270081554970125857553049828819279709376305931186998420322075168094083366542479334467166378285142191387988529702065685629414139394546846849650407495689632632894403028373661750979177431445805056;
G4[135]<=640'd62359935515543997092854801445964750530723119669765095655840160895512548964601433030724677687488099669398139495511714286470486143075011783646572807535119924096909669951356377922332561948809472;
G4[136]<=640'd2415355898963853765177740450585951167394151314262764998432308472724351367721276877426062885416808812757363888279005600972267264453934252579075431894877776529932172042588883134654498351137948672;
G4[137]<=640'd2833281654248596449256911448061579349324975305075876671195715693796466895331710257635241953584189755361983201102874636932074486177375595191751213294106757110993787921772191799748710937604947968;
G4[138]<=640'd552472981529364577863876048214053113356930674450120610914998211262459301061876208545166993689469197814163163542943100713002851299927664104493188811581345642778740526632352276355358091789844480;
G4[139]<=640'd2419271150557985915335468467239324153155805999575302912979588249230512622177918341197012309031161753691065844062445672821707796993756996825071899181113890192474890137503762524919305953916993536;
G4[140]<=640'd2352364568789015696232023315263800757887260229738393355001401688025573874611016995955598354446224125185696636358518265137886218415546251878146868784602270797565611337997588136415889692536802816;
G4[141]<=640'd998033477177391300805960775003309468312587585544442501693322589126500416382818976149680236359042125238739941406407841339123937074592543706085320294074290495300277424563937959233383590027398912;
G4[142]<=640'd3270343041105099564686348065228532734460658036994175456260274548870507791355713336491233166351989086626797722410969967141190997414805233245247884841723126130289605404069446636145752105251556864;
G4[143]<=640'd2342895525646033417787508348473280010368621136203830768647261172508694624742081235067876791562392377414147916226873810310649134631450091283817798081329226517783165229987651189267507495017436160;
G4[144]<=640'd33388030449761208033812698614806064685464614912160346136524755391381195831823832124283866644823210464800224130552345097657089329684951237288785203510385769454001343539968024110655723946902284;
G4[145]<=640'd4348576213669874358375174928935841630028956272699301550066379944269694784470206107026373181556968664055868842072487040187168911400622471604628302822186872109724271410021877947298799382712891404;
G4[146]<=640'd2298955320821051264025330627801958415034056840419690000221450112065917229577694179289720271397115373399635259517648663036965624609792816594921372316581783531734892150506501226272178839425857728;
G4[147]<=640'd8858803306764131517345359213383648569979200039821428509121230404285941966707321051056595901337378429070339993356900262447279413781953258442782295153795448131243020583241436519983082440016113;
G4[148]<=640'd2283378444631944929898371580713313416932313670422218495587005227025565373581639302358726915942653581601858013061308420483560185246434596744916079588665282961327071385550168326071696336539665393;
G4[149]<=640'd2283343633850229861062117832169542963070796152642646771693108856646943107995080620937463829226644857378857293196423798904556991939144799936810713484927064653700274965637376152950223737781632625;
G4[150]<=640'd34807568191044027819260777763758229695817220886880167663379798908923304803464923219506464948613111385807545232334427251504431542065479292659263286855723052616541140928132214411408917871664;
G4[151]<=640'd34263284552976403442832645728844850517537068985400222999510591232804172962167820450861350083152085366681324112872024323014402546324147240616697550213762752863766802406797806298272945324040;
G4[152]<=640'd439015509137198729869949992261592248365339577934793398907701725680769149537594309181585889205783767849290329484412374551426379427770451765753551816582305020211056055500359880163700810610368003;
G4[153]<=640'd2305734096918028746711020747810821193246378032331294703899035702134840260329546312936389401788165963828596143314656688091463676411649252790936589728333499190750370392177509776307880491007002608;
G4[154]<=640'd2334725325212130797323992770028894166700584482023004349349710322555462769076617459270906013506734242673824743287462317271295040321890622707198525101799633085031325643968860728507837411332376560;
G4[155]<=640'd436674773095655886132651568943369543321201108506023305100832285628881038315711223517264002744671380712427890871739623065392868595577275664612393347445679087753082245418654013748098590524231439;
G4[156]<=640'd512418487855941981675702105774793182654778475915365851801630130447200946025100006934795668760230397478828230300142810105395159302015921160511998420725985255563264234070710596355929028373249567;
G4[157]<=640'd454670714668446940173548937545912760692600569932842245802477459281910223291467853690032134952952357756316052281931630193879547813679500924542928141709112906183792173603423071299052983824645886;
G4[158]<=640'd2765165101801220919340555156046354469536707227274783748058271085861455889756983587822636842996882511549423943076897748178750746487790675164552921728538341409062975599125677901756221273774489336;
G4[159]<=640'd444489195243125436271667155866330004609767523753627962081750101419774805536427901018391847825824561447898093835769026039773050753634038148237038325185080739117067415106080414371696555323219967;
G4[160]<=640'd231151289528966182818414055140347380076197709492355668719293069206619229608322369428530171130751084560419068652678545628158093108858264939380566458393565005604443193949879372015962726426681203;
G4[161]<=640'd2423239639563984987058918032484386949573833882624046647019876977954146620046856417636146070214992802155331204844206093609179309110225352837956150515215453521169770953440683356352376822766238065;
G4[162]<=640'd3559394285553887058825602097967893488625333999448371263405420282296333085755429227002429131897094306396121712207558612001604569027754604564641756337989470094517666651878600434084038370069051440;
G4[163]<=640'd1962324038138964466979930467207622818718539094738074543300082872030755075681661652280209401923508634818034901045854446225313385587822527459301595252056959227376097778392074904327572348332931856;
G4[164]<=640'd2254715691207444180285812202081948257886910296585600694031977663341884351035864617497913728111281720866007467214171929378656819038044364374411592645234836066470667360327909116716368049813323544;
G4[165]<=640'd1844652412913428400049124825875824859284646699261061718142100169364654358002243844853035020047054137073100024472555766537321392885618012973443262328868271443094869655238703716756677936340271048;
G4[166]<=640'd4055628846859080221179847098273217645220329433318059336651892556180008334495574747163268528766589363643739579934893448921771928795045693005105887157692154811006362162607208216792819934984926924;
G4[167]<=640'd1759916132605078341232292308103759975515796315142373964368805265923162903505023409402519045257259451351267553065691134465787545977250271746175456856493560445925943770852199091014391020436584142;
G4[168]<=640'd2788026504754511278883896727880122360643774191309844150922890797837100490990074823443349240460198810735051845983605806740208812254975420705954220945792668404450058930786419023836106562901901304;
G4[169]<=640'd2352369072853685358294400741888780040464439383088420188415734650455704806366047111214811269335356754282540322316466678402178068358844026700313664279479101916915718739145907921699702508898680831;
G4[170]<=640'd2919280386539026784044869535485704138058498037983672827595069121117750183996014890597796017326839745751221526896449424723921528084356221390657012160151831270066012115052991016894527754158997443;
G4[171]<=640'd2121882792641178108236941072183967318338513872833574952172235837936910991367243760874227326873830008220451471953772046261512377317109734719027677873721034249963463490159491058291849739789926384;
G4[172]<=640'd2108560757521521329614385382659707159692967671960926034207736820627333208680939836800403282967931818188207652660165092684546956497479251868924146857091589313688995065261789464562455645259825148;
G4[173]<=640'd4330606346253728701063782886267425859924558073918510559007022897011320352945315137770627030459254379451569161059289885270978316037085896227238910606244278112335054742280481099698651522855862143;
G4[174]<=640'd2325349836714301151986768699638574964630958239353293794134808787425418662645073194215012296624794972549936960701933195563295267142273793983686124985608312710232178509683068435640932566170599423;
G4[175]<=640'd2751415422106139819407717497491833730651349037441734908649814720411935737336107304719688441679318709937942524012087320751833521841126385026034025102553943383456558806601110643812473431375478783;
G4[176]<=640'd3853023584684560651920799971087067765306885375567850562642067591182047792101580316832333879694121884275106686041304814219306103081008769385656055635777209415645851625169705460442243841138884601;
G4[177]<=640'd431074824305682565515953779615552887652583412653733891162926662850284073218331863860171744261366597562371969515170800245322221033607260368969503621310115633066176602583989804172599995211448319;
G4[178]<=640'd427728875904341936654749589007555724924558330919792997332288530708010026192511322513421838163872964033783154783080510629463782729354470799690982871420383920205214809874014754256206513540431871;
G4[179]<=640'd135975475676661258253981353653123413936637470996372132539228891051269774224671475379162924319728681779482672743592126560140863215667026786534232245931855315521042073857850558995233767414;
G4[180]<=640'd2281220308815247123405484385554785059229930272747278534579435849868462437639028846903227107843434582681583096546684262442004952722838422315246035452195147481928623857173710238667856384989593471;
G4[181]<=640'd2299042342745477578165786312324280238786610391684070808742671644259340561929761139187273046079501285330470816862230529020734458326620385511215966871398029198261237651453068135797706564002901759;
G4[182]<=640'd2281220308815247061572884018634279713598342612546004693622897752746257431412729138039974987959596603300055617082750258646002737542030207992340282850599496640643029426318360760332614323773898744;
G4[183]<=640'd3707052908080245417408670137762781022199851648771424509938719402250774630466437353435127260655308565876755663842816670033523024490567279480312506284617902922694978020973721642768460995266346943;
G4[184]<=640'd3421830463218721171641608712463327461829467954680725971992951434870788238605155396813204728542136098014121229517482443251895971090526774547538949872609506350762851609308366380520177585767776127;
G4[185]<=640'd1037378768523912313064038017041732050669896923101815236887104251053202151906331979187535223251789180976230326691423973519993955088382050779498148704985596538401888988976214767042559;
G4[186]<=640'd17822033663105389518927200704579080877566000139632344410318573250652249441143698499186176158911731958497789183414058924794783793933768655305402916803180144200420207805085256716087565603567615;
G4[187]<=640'd17822033663105389518685667109377078092359215931023129894307052742842033424840215632281005551887249952157011475456520412608948949343720639631138019405945104321663178665104709398566125971701759;
G4[188]<=640'd2284566291205529115247908381784193313443102966166705685605267497219488604097584242502695353888192583217543106438181695791960282251829298612479943438376466842596951595381658004139735174961168127;
G4[189]<=640'd538002641214484278698953821133287859241946280977049639746910121082937938402149032933879465922288586589359562873924794751249048910781336492246641238744220671665624469656106431876897300560215807;
G4[190]<=640'd2837086458600259140715742347862948988593012649000421834723650244464245027690614829252946331501607548374977535849798714844037131099023660376318744952201744532002662673023441436482882526848745471;
G4[191]<=640'd4280688871135818398889449334900841950085059490616813153090184323310008962574198039007422864988403410938292525296862642999009334847370197966210434700156644663672235792177249980859634857847816191;
G4[192]<=640'd4278283937260394111099739024100570140208236615301599029041475719339483773477261163285378025439479377603889949226343217068256676000880831187106586236136745505187709783347572549000253886355728377;
G4[193]<=640'd4286194744768627262357361633594658291784316457494441648075172543776854291933512737252539811575646280195887401550050689228289568532658008683263470236614753923008800092301678902245555180809486329;
G4[194]<=640'd4339658670215168372546802436134284259646904598498452975933861363374381829147924321555084577480985591708104447223436209165639150575018131998823216658188695004517447139441939890648797898925408249;
G4[195]<=640'd4316826365127170298787497889913909528258835590546286750518413047076249724620351571770339156626852914030788201282481499898761292726581588684348779197990857131418187720221298228804229639155154939;
G4[196]<=640'd4330754180008503284114619597568561885500542007310845219462448898529120604984073021196254765172737298338443527911192732188329432060866055955109244470453542475446854797724045390816704366160904185;
G4[197]<=640'd4330754171526955766876900080309884766450090818826796913791079813313831001800856604928432491829986290628664343110533816868122268019813385862425267136782441541236282701367129289139785256558133241;
G4[198]<=640'd4562375334397520696102036272509010599741635643251800679196180816419139372509164095554041190774597732275212125329532941536792730505122143068612113031961370774457302682392647203815537471953829884;
G4[199]<=640'd4526661649750790196705811082999966006354051467525859325674863644076440073052157302958534929800308988972642600801128498429016672830946127931157230522091306062609159940911930354907865996071010044;
G4[200]<=640'd4424120080866396825674352402007888257475367288396124217579754963055824239819616180634392605187332084925022588534977990737205840035738897182941592914156762235018747708591285876701548890556465150;
G4[201]<=640'd3421856569711277448232294052862296665079565974124974203983133122823568224355182038493152773809505134806934577282495322339314785977706787063929678711840832637654206006444233959551426505243361207;
G4[202]<=640'd4280923324214302551615294316661191147261649598408750636959482841024498556189559112968866675554169431501583377663378583025703621707985247617032230042975445102738228553150926950201316675158003;
G4[203]<=640'd17821901907168420525996187229149973741157224851932027463816651317022955038780822373471470072182219006291088620231862489657618318631993346602706017295375621784871760635273495507339395779788798;
G4[204]<=640'd17822003892925643463733190928524404319241712115108450130735558526596565791955639953314449974271533139040748213592861678991124724651098653595943852429139585704890546314557315359955824460955582;
G4[205]<=640'd3439652496878977014799591666685465986650891920261593562561408024178229983857585011631700658216905187988138034578337710873756775609494477528700671053691580373734679761877913792138608938567335927;
G4[206]<=640'd4562127305693770998285741497635204942546923925633875966011093520745634638768674312183354480685356665282215386946073026641974977354500453711076128249903745884489889005413128442552715706846150514;
G4[207]<=640'd4562172628761038875701985514651790172125110432611050509941285788345013577035869370997406685647942304041987679813854510096501101277817319744579684942355902701775016103324267914001692393612509183;
G4[208]<=640'd4561981306503162520980442974768784002756737583691915695752319407444659379846142882855188407281208620267028684816783944254812348581115947047125058830544411281527549690295348961178429148352217087;
G4[209]<=640'd4561985385622726190444898519205592003749602143546676913586553831746929195920092184577311471673528999752448866388254315641370004279090642249957413768952013339787770992457196910492423503329886207;
G4[210]<=640'd4562431915457563854348875052905473727670989986996447720388618322609804950512023186310160447672068978014134000283218390890934020523191391443466870240973157012688735558989998972621736366607171583;
G4[211]<=640'd4553512196461164914744902409657627379343117579693472329304378212680116177724410815947156310805729267646817809336884484473629333284856669900991393263708682579168897769706387744630771564819775487;
G4[212]<=640'd4553451285506342842897795753429688938897233424032608355098103283547228377049382510338136727544353870461484666393941362581170129161865606569175458223813043196255548455846456444644778636050694143;
G4[213]<=640'd4562334020351459196286425426657785597516654104944041902114844483790297758298464718639069309752920058127020238383140172435763712266733389494378676418246302306293679799599033443397439513197281279;
G4[214]<=640'd4562352563407987830484339478068001123031395668439450840887828520224249577092243826597269582012473721869699264357040285120065880602530345849512749051709421675611858798070277235706738592576438271;
G4[215]<=640'd4562408052240608576366728675987714764100508872103648726902779611091101150329094571846481549068509994818409643010615845927263803869215970883471739726138959212829478566923974483973706430069866495;
G4[216]<=640'd4562353662900976534007766817215106270742865951843571284449124422446712761353687392843598023193937771166544140722702143703013920824519637578233659557671056565275388560231691586729076487656570639;
G4[217]<=640'd3778262977126535769658649087496079864082646513954223010232351406918058529710162679043825379390604856514920557867210484371863625370201049543725842814124766137143668092764478828396357095286112239;
G4[218]<=640'd2290027978936300889448976480629086367240717412585814662645169167072152999651486204584225969058409304938534017644957338505888786376733480232397287616668968144363888272976712370023150388087881509;
G4[219]<=640'd2662318694869290108471443348721669971269780602118580100992211379385998649495041789717231464211563683391313193890366445083136739946966334353867111348136433772399238895654469895662297965854647;
G4[220]<=640'd34265836339031228888610571608339072627666235332997393462396141839805954789687202621348432220816516538804540033767589993618910223622616672484888504399569215654006693848590305699841541373863;
G4[221]<=640'd27288902337437808269747315782119288325835870698271608462132465288331649539682256020894741430739004569090498083967350430406164138503741839142040546418555186743790129432022120822453537665187719;
G4[222]<=640'd34264779503967166024652310526880903736956888590342110710586386797303956576862406479373733651346935854963603246388262333059835912726808009891705862709374600841399884246424875122641316686200669;
G4[223]<=640'd451750071758515069137498378832847670655163755436365320833848361535765382507615832837488705678166719589574169459869492631149943523032681580150941633461834840786850150632586681132786893325434756;
G4[224]<=640'd2277044357427060483109541763292104280505918006622699955268345275548598016999225066243917023766388121048297165756539673398143010841326386136845038408268534055888646601974382046492348958303915369;
G4[225]<=640'd4553531776299507340750081119979379296732611192425423289220276211117174358880813914812813665710518120812765149091515407302457692977668358001441694363146777179241022903310544582616447739726981614;
G4[226]<=640'd4526831358923354338618243674984600896107249346957631196099010891521673397936884018781204996530537541816747064047894122006944708758257075729000008288065413823686370867449731911527284258816528215;
G4[227]<=640'd1817986668155464371128114779285940807784491193609137988530343748264391920970458704141540272768343635448886532063341709985196179223090047575435443992515808528835659137646321734975434882069792354;
G4[228]<=640'd135684154653864109144637242180230680607523240620098626297295082433248760410475133343374487713011470782133387744972076815671214868087820414803536423127369165446077165813555969193593001100100678;
G4[229]<=640'd2283239210929169219778744530037993454971317114944248043573634617887478448956609923235529570865928523470517444127133744149250504455123143140183071717713339382314009853023577082443909021824746534;
G4[230]<=640'd2227751021011589653449886338708061768800982741339590563188725796882525281028724012201656027621788445191595143009185879591817939974655992125686498368037358059846416303730831941075417745429717;
G4[231]<=640'd2117480373473810369029222140704984105473486547410863797403039749121018947380441028430913690207931897916753546613287786906145795362184061896101633126406674589659667398183381078008334415481649823;
G4[232]<=640'd4553529599197488903215680366273043417817602916755745601571434110771669243544001780882000729221241693558237197295238655764626487522460604080012762997341768716725713904306161570945755031478126636;
G4[233]<=640'd4562440615497644260427713280067462941890065887234248945827530657189237705631302428803730794113610044589621759055651636158456981694880926374862390128661536569701338704769223007973701560401173009;
G4[234]<=640'd4562440615597247830072425725318063931079709179521692284402816508123822637578684118972190373220897620421846195902607707175870523550276887962585877534786696001600546563650190455562760290899253007;
G4[235]<=640'd570305072953800132157532948360797382849612100602692889761711399170136446057814935254328919794985059792281259131254120444898736458490273953738948342491960567404172209925942643875863207506894482;
G4[236]<=640'd142576267719983556275441385264006773869786551475967987321781002222002130562331161480995674922402797907333522506616275232032497460797587742373841507308508114103660425227316115107982762522837893;
G4[237]<=640'd2342622749918284661827177685471413242718632326203557307559092780357135506804493510599738904180872830988440210224450209837605967991181360299839097342997557468787960329400913735800124755436824199;
G4[238]<=640'd61541709990086372026867064455696316358790492885408544847826208489122730885523901332752540422369669436501723661403451472723262901153670845941042868514681234901750611678850268671559531664125462;
G4[239]<=640'd17264619210731919932255461988798928799140840824286606146111751467701219806852840202807525043878514669026863853637810761468282554259510746037706069863828020735091367258172109838822494111215135;
G4[240]<=640'd4544601188128067783812308056029940383313149827652028930395112161259799895149769063016899925859675466611635066696744517290574548343023763265300341824857076997271602276046605908086058404671202841;
G4[241]<=640'd4562405953428082509583606942972103047113909120616148838623380357439767099338881726370744160352457082333136249589570809502402525123992783286548354288059566814883724244554360241401819013389191276;
G4[242]<=640'd4562371969094624501396256784791714879481804284260067991767484926697703523194886202873616162209519764786443103498494720433969948907550172879328695366459173794066079932593926227869049686320587049;
G4[243]<=640'd4561884103980633605957451034801926125991554765292478551233355046819756350142632745106529784720527538623553719744036589948277203715632204415790835276583412148266403241166444647252974791120085543;
G4[244]<=640'd4562162692231521898319147664088838281810601990349363738671899103112426928078467591577931164167565014114889969019617800284431699061779843929909690089734391526798784069457847434737112428988170851;
G4[245]<=640'd4562432459342625547158752882635187068230704020136681277146256155682197575526315326246561340673352462235150944690187951985553584048936378409196509867539164119617855222604927123550249050042141165;
G4[246]<=640'd4562440617622195216654810640756695000772190155887603845421955724532840542953146223655782594876665143271779039412293308229980172858251599623140906681913915774447071270521553222654599381675494346;
G4[247]<=640'd4562440617622195217883724138170121100317407038058689959358376767089072339697720001517779224351788674944477848430802155028128904033420703211795056335686273405175778958742778099058063966251799044;
G4[248]<=640'd2157579950276900857596435081079805831215185848675160707590802397475528857511977768021039970982702165857252023489082372164235835120266601983927696423275361454528517556322480519228318571977021468;
G4[249]<=640'd316898036062862162625741863929584510239008035964697361546851190169682313318468731454079619878566791409413576990997143569708159778621795894061520303561983836496939948408523038798386732336308939;
G4[250]<=640'd13432131411812752122778422592921983202024457481286982692851972692691343411805410224722915856481653920106860546261973967862397390258395063451472019678557725618421321365696705897892744436288595;
G4[251]<=640'd305935483862456097726637788193631844600457245256065886401793360351591855724164847515377732629256566972610356733325453229398546238424813078625047546197052821003010090932590499929142961256;
G4[252]<=640'd1670823622937395383327184457454613256134138749886716433807302638824774567127552894050032136967358899979496929279647509244393896098345546017498448921065272551150222420107398257748584958624998;
G4[253]<=640'd204222558238046945436311603985194308603201545450244569145809554161265507866338126866041900161531840168048562889706807929812909014227033044051245603920244900229722175047522371156863354920;
G4[254]<=640'd6224273353309224059915840752882569843615705300619366067942018582078209504202758497347581247279211825547852065533033564472127365818694997873857197663653101620505750877191006856559718;
G4[255]<=640'd17822033662716372434331398747132250343398222056576552584345512874835371078952519428455916289280049460299087282524528518779269868985836111062722171842992182237383669668176741413404161010729399;
G4[256]<=640'd24281909467732315047631692352532701332356148713125808186366020754367324806879023339395674870981417261296404548109647844158464774950977702843167440105837719413727028293521331823347;
G4[257]<=640'd203956989447417447657075756019035488526595925586147771611818488383471663688066354002805314887222213367025600777068705469861507238557914363053856174653674435197067275850524295831005109427;
G4[258]<=640'd1122231182191006272188843473958475707161133445788273370879384007391952337724932271348240373540039299385034802833365532732707630167811490218481529974162908807702621480368161448342144299063982277;
G4[259]<=640'd570026607927055878287218898300298032298417582460023802792530177435739070637621168814147573705541990118431437580404708107534917299914643824762457936423914005009254616017468493057324568695908507;
G4[260]<=640'd282925023340046417195833250375849582717621838582919767417493544120427349621237318518111686460746811380254468135419578207742636483674706515835900244885723538022472258386723403011790173893623808;
G4[261]<=640'd140348727533085673693629496034268028317852634285358670154114761305841881178942975600103156287585125021447637498879029836420262651278178992526285502217804772108343423991766470953200335894910285;
G4[262]<=640'd66832643222881621428617464923317064418374893379515107302610735091879906262438549146349275475766606965311298669742706240535085554651018882116034871701250958553907645192392422128338343884210335;
G4[263]<=640'd30802372756785855614779500151741228235976882708707833690407169234139705817943328609083350119116935821208353271405921486702983186337960955725044906124597775132480518589865363403551875588;
G4[264]<=640'd570305349144454181563842934944256881609352521880083291730179610324691186550914572671314756003668499442505764484257158206149892114458056497300213255450011984336964497015590826928033132169315102;
G4[265]<=640'd922290513981453266295445438557218181376419009997265384751340902825076483651743505889270742182960716571265608609127928892634311372079512629575190744804659143525319501694488992697022017161421075;
G4[266]<=640'd71271002263242398130103637003262793719292665680829682872049013871369094487883888759083827958498562882250475740196768943984888000470199647399913048500642337261306024400234181206094080282567146;
G4[267]<=640'd8911016827273344829091311212049885998747442180453186308726484266912599206912084573510343429123544795195011214562839377291645714836586684403294827363529589975415256467554486078862337873842688;
G4[268]<=640'd4493380236382980975679034390656116939076569498750047995198933903827921467912043760759329645104040842946825189647741232030485823232500324668799268994335565297332597703852288578559327251215688117;
G4[269]<=640'd1131977605787957390136274238214823384114566064839821762686684381796778285186213159711200538148836491136317781368572427689641856310162202214170004978534650675271161891622755085676230582876456180;
G4[270]<=640'd1138391101300323791653944204304467657975614650217932049207758524268004473244638478793959820778375972214028407800567531427727067065156852857945719076408417843715869991310627017225543098392192776;
G4[271]<=640'd1140057566923581578533896055591179458062387792776945108711427686146816986850401737423024463192298550296310462873826957106470035176619283048932639132584808885697911472132224951296585622922277446;
G4[272]<=640'd4561361548812623419473672878978541360391412924102773409105951147274172559682196697663872054821782646401861779521513237570640866007955517724518847364722942377035835223728192129585920250585564056;
G4[273]<=640'd4418759173349268134665180912698185391173643108679521955872334675444468301485868052813315795394997692304758797865655952586115541428880460521288294780214558507605244087851758326426034233928419757;
G4[274]<=640'd4561892381168721445073945115855372538499235960651805739564952611128867304896054188432598388189703942960851313768576732825364353213883434558875152777225258270730005033831818836535436168406770370;
G4[275]<=640'd4561918486667460645327869584217420268254234827796202851180210139836962103268626814410840428573986974859613698956540615948184932204674997701282929601832169996934639452500755007796667923898585912;
G4[276]<=640'd3439791729392670117203178064628868036898608551097692698309616073544543827707368874242126967635832721088615929974793734458491972546056155822849504590317894896780538394470893072029441503038780454;
G4[277]<=640'd4455100501668286713048238072327193925506811962868713107807280739512410172401065045018957594190288837671888064496713420296956974303886282709808592271133476361942131655950993088231852316505606;
G4[278]<=640'd4562436266539760089815748008266046270706885616171496080405572040318183759671604945347303006796828086952278923895105800508650492560752213620991986990473529415869970728184335550932829313986106225;
G4[279]<=640'd4562423213292448181731451173142957000817382696883276851419837015255583824754232910622469474778682465482400191691079493145410591103985383270261464324286552801593413209767577842006641260055810132;
G4[280]<=640'd3992135540419437531888878313284584854283955535678158397296102969015944694085657507951072118611207521668034020532414805649572677725023758128724280694686033473082377931166958870456868847990415891;
G4[281]<=640'd16715577853158296829945002380591835669988284856679170857158391960140427802050766013874821194684573675238833826283035419612192686043341515350374956614183810954827702525062065190057;
G4[282]<=640'd4052261297735344686047273304385899543241119491453011979113099743230133502794433833560446374520932030574254743728157845406220029925994360972626731463365514111102714891850282728641;
G4[283]<=640'd4052261297735344686047273304385899561534103469168309654632373577643359105626082390345900893900192713311773158670380778237087846771288833310067329852761652592013888768439207925292;
G4[284]<=640'd397121607178063779232632783829818157030487646181322939856337426513681768305559774580265488941160438928445745730877150352564233533819708118865624767931542355694836117689886558304881;
G4[285]<=640'd2281220308811113818365776744228889851539831797222526104680560794457351146588431286536936443516735425852399709295044425369012149444726275626121239549228123815932735325074051330755110643090818012;
G4[286]<=640'd3992135540419453234401407037745243287468010031038933399037781534825472787806973871021383170349660745662114378029329606171622937198727379552640889458195737567148694057980830653611906294114025734;
G4[287]<=640'd4277288079020872853656862145858999873460271899911828262115287151771994062962890206364451060145880639999252368991112152128653993743969900831705744747077483442268970487205193198993406607603376926;
G4[288]<=640'd873279649466764512613227694032315575498562062563790768946417098976343450501370633180074626168046368593266664334892697183188862718452399405095065733618099848926975462359187074741884355030852432;
G4[289]<=640'd2281272521800359677838646325507946785415772805544371098169766596323198100454662434197334871231535092856090067592103009798649179902736578342576617512723460268623114010041026183980873477986980087;
G4[290]<=640'd4277355520802490299186238461773487894809253535135537513924922447887409406894256569778036809201565801129966129864434349487469379077726825405723243936349944324793690021558238749679174874804382659;
G4[291]<=640'd4286338058563914498358663184471531447308872376194451947564046547428696024465770743071120939206834100429862962410863943263951883021552060874070084625162738159376671875938814169461280537757611652;
G4[292]<=640'd4433509070934906631010010687055702120122229318366916596145165298327460567747991286034873718555806809902041386180648614265900103482910695713252890690111884079349908725373833064042658310059562678;
G4[293]<=640'd4504797476498882624061715563578458438568476643687870284322697898998407680185861106312202428364125963349376526996490359541829640046338324829148654465539948787735604592524771572884468943788967360;
G4[294]<=640'd4562440616692703731211829182993511963426408409421674419914690697149900640301748301407472376423702111208754103792538876652762591669396196403277263051734173490394600086819566797693083887338004558;
G4[295]<=640'd4562440616692703731211829182993511963426408409421674419914689277543017250444540197259410095164845951915934359366997740384796089985646793626153547758351170475616310381314717491252493735448604695;
G4[296]<=640'd4562440617622195218641171605700291324893228507248462375936995143142044492365873214853201634285947885756364456862582963310224917574181929621536224445542427205823523536306028209475426150062868446;
G4[297]<=640'd4562440617622195218641171605700291324893228507248511153258093830520659829832972393022172538731837966017776751185259276294953497502160654668430403179375101162769304709416363865597409717434008772;
G4[298]<=640'd4562440617622195218641171605700291324893228507248547736248917846054621333343800729470741821433876610884092107238574733245229424111858150087469745059182630381471672390733819708371449171149887241;
G4[299]<=640'd4562440617622195218641171605700291324893228507248556881996623849938111708862191068576413787552810635659319172706648275819918243578664206617000380390549907690112605974305649207535780193773825871;
G4[300]<=640'd4562440617622195218641171605700291324893228507248559549506371434404129736346216205902498586635396280447781521884897932654415176401762599682995689903005336831868313782737953621109876965805663834;
G4[301]<=640'd4561605209794261467075258305235380382878172374049091152898874929944610456253407879553848511089311695425618418861775877352087388577361291747835200478295443469243409831415115589812538415231647240;
G4[302]<=640'd2262562867320577157681855425800467957443693946618319477185509587014713161312234307552742896988154194488869251995113197901164883525658384059065381448714012988313194669322580533609264009057474850;
G4[303]<=640'd441234567787009785396541528883795874285480991755187526628426815379840990259975127238120739393760786691194563437661656208635574543194526740765147495808583222922334042206643610514320448687780153;
G4[304]<=640'd4553607920274770657814067439326493344213207932803107620366996023071195242622219630167256978941737597693185467054857520840833515853995870185591604256400600678807025153625027184373376311542695270;
G4[305]<=640'd1905723118226560350098242485110257434858580106380773491617287243911377458927351024237806561034264177250048845799833213992580814005720876180468788403616291439169796189878098739273385955650;
G4[306]<=640'd4553668835428890827199081950818726433735139109178593516066992420346040318835742609189521188574363690992116588359360145860156889405896380682820507447826656836163620720393958955330083414324364463;
G4[307]<=640'd4553668835428890827199081950818726433735139109178593521835184602859433270647109833042596653481048942284992106938261994980941515239879142109240160635555228939152976488533922450032210517003089983;
G4[308]<=640'd4560769801966327715509345004770469440863116240949518709898582999399958961470376701444523883678333442489421511681357115552207796584090417970959165305097192891513380015889105322749481304853062950;
G4[309]<=640'd4560769801966327715509345004770469440863116240949518709900036585458308782808001186404587301344821576191501443878243491119572454231144286620101616167238782588697654700551103389149351507689785558;
G4[310]<=640'd4560769801966327715509345004770469440863116240949518709900036510531432789320269632797450435304223442109753435427931654546499117196941369895712075134608873068172287639358760119801883909925900704;
G4[311]<=640'd4560769801966327715509345004770469440863116240949518709900763338165115382154672496769578513694241728825500850392476890563022187936719351089064696641318480854040213089101054272945609410255600845;
G4[312]<=640'd2334721014501365707549050856655279257846214552844405178559204622728974418899162114952393443215090156342476248566437953919196154010777077776698923757924001790274462219921396495369504460997925667;
G4[313]<=640'd1071480428586683184765721817022853694994299053081781079549073810061473068479869316567734126931106753205162767229486164160708550824581828972527194008819537408336116877909192717389063196499030454;
G4[314]<=640'd34538841396888730893586541895693889674564991419567803629074464187631166403139227035348214245098771983037298385216823472145030310287554212323545866233132107657796282947468719909013250557110;
G4[315]<=640'd3439652504842161595258916738934668031223273621258934689343904317300254552903387374599587911262769463996575830612688928831019311989680038977191854020575029280042255487568518113227548245462579242;
G4[316]<=640'd21891383511935872739575325486914906339771635607365906622923163046914852996620366677127819734922301544820100516878204229496445951758064674735864361176377202759199507950434518459218129601730;
G4[317]<=640'd2296884205518464215136959658022963806853643362450844356424102666464635237029968991928720526641429045726387757175419094252031229484244865969830599022226784727441168689748757613977932696936521736;
G4[318]<=640'd4549073820432602871463633095598409324431306097036649037983762530350237531856631869536446567395335237870755745722848964106883706222875470209439837894584632028416538583541699234298341327298234377;
G4[319]<=640'd2780306834689947431797730432786559874608966337263879994279376880633318026175471849030647095560751857754153443488882327825448483374523102467809591047269944773309769316665585857691172911079117078;
G4[320]<=640'd4562440600625779954790922345862061724792056122714607125115127864732716527962274731878735253370889685272221910668357171336326953789955572037946859484018406141491159979688534457575445414156052121;
G4[321]<=640'd2025883438293191539926525358553244725139734811822453276901309643784133928642923090796030030197455429060063608070335818537648126652753730451423687872325453204443489273759574542542;
G4[322]<=640'd4052014023954421901765105302462429428103783664599590441403845944439988784128469128723854414201679514210982510076248977602720594301718796776728409569561014680097378178200122595984;
G4[323]<=640'd1962814092624445712724953861417646091867941005556260337439421015173133079700949796198182587495005977062288289460019201099085352949230298293022920577325917048416339264539387275973;
G4[324]<=640'd55282765180607315868479032839477138785811839307018050282199269945272493075608087493142786254338926167669628956305058111046867039758060180197297185665315553273949340855;
G4[325]<=640'd107269004826365920536733424261934078083215578107604415325129703464288809840758564333420679439562473016787000015061065932812885672994862628407763902066501814;
G4[326]<=640'd69617318994479297159441705409245167921747307411202582954538853771640275015646533050662957429758258300535139540516112604486657472262300626163471410520829160601040448180100038311111696979290;
G4[327]<=640'd4348576212608878832133832489303913755933921365402742316526157313450462606623736656889419605906232203686153505510502019481461574452172432002587511817058328782817084880824854529911896599349439236;
G4[328]<=640'd4526796261361852062881681702283640178689715249638604259891652637992435134218328527609558816017892065238834434447818861452412230665862117079476987185757867204436572474278301486414504710369579151;
G4[329]<=640'd4009957573019715321719726116966917427170658797847641409961351305328159542544339597991545174061251694050231205689526668312821164686511982795339757200674857219926385544441721072538415395606789550;
G4[330]<=640'd2851517226672026423783419658297048956549919686194047007672347159110925179737778738574980631066836918338412900278377568221406499214821510355785150136201888839700896326600259438596073221510578288;
G4[331]<=640'd693949786819423061403159216138348882319006736572539717777620850928927692759912815111927141809517004298433834719917679373641302848735130559081432753719814197231217686636421152531110057676913322;
G4[332]<=640'd120316131552204793240005193160664089266703555481977607299945297223012792327883786122802479921287764668194791645444281275641248978894691872391739499523424818861703374062393967441789045252314967;
G4[333]<=640'd4529442220874009158494435712998780724929473635490963723197013160225724646893082249832687964420251389414272352304185498123431911345971784833791514775460984168916294013495738661005727991479170118;
G4[334]<=640'd4010427490985228356162263933773407929087717957131473401081091694497911485396432514715167646260145478109917481056179608261178778570832583567885182511330126721873867851359921020040826511276132941;
G4[335]<=640'd2212559684067487758127577362751954215693076486984457690294989112110066319637721896083108552660471527316081504634380443858923736458965756872430863643849788657274740491812243183008238746295999696;
G4[336]<=640'd3342717314451494254021811032866166819304899469289108612213482994936156865623857338313388096097097947261063109949245689079071366040909787796496806239314239813723892196037473950878807316489832585;
G4[337]<=640'd3350472762234478177721168456591349411422283006888212019834198531410591296266706950737681602122702846274364143253272725422380300864391174306120032586279207767472097009783755957572964458863405323;
G4[338]<=640'd2263433037066877802870505301963539565467577279505804049301109531100470630787135761532749978673294719755354746736306311244020852659376179764676355559560005366422350202976162443937583719512478115;
G4[339]<=640'd3203545097093058422764606224994152110093160903392020958070243702197093067016683312386674842661047734405537095852592600584830978511784690486051226011449782244606507174668566342727481601324364144;
G4[340]<=640'd2049459344035498949713900523591631300141338489388683530688725045038205525596176592925648696722335985930485805537484470182588857765880590236266045973076089299926570031450722771074699064899667911;
G4[341]<=640'd3207960246485131684952640045683142292553052268071799422000066213636672064758506288326294287420336271962373470662080423061510656219978594403136875404468190695547769889443814310082935926458566943;
G4[342]<=640'd374150020665283731669873896324770154969919386450354252015301172748828202580313583136613988283601385851002225048947763701525238567110026200854363737373432764250570107335165935266999751888096073;
G4[343]<=640'd944524298787087872259192324386233761154593389055922212921460028531392728392806497679907116808225666290274705005787882009766828278904561123004015011309884813133913282410272374908458957207047426;
G4[344]<=640'd35635612670595076388723460340833829199015956769302164824523239453286947485764951171995366988021619639350428516230366660154447912646327735008282475044533106905277456048469846088919162102026047;
G4[345]<=640'd35639776792467426300044804295246680574798557146826572856847654597617760983585491905419815577537794042940200944505085783159715956383440010591417635770978784771629402354666492693738072454477559;
G4[346]<=640'd2334682186720676823422869217307861382767161830474950129891530274685055526969358766325778100475028837899415820428272893565374790020303077823122941370728124596024875768326874366186707337389811796;
G4[347]<=640'd889109967712001163757364481528687664268853345053073002132428877876157604041789878020487205431015322755938348654387164680732067075114685635005127338309007413289119006535568381681411638578816002;
G4[348]<=640'd1207651639933551738329618277912521388739642753171582408555691039977009319510427729687694626305290285618439139606901112814542826604750949596680896082255163938659025336239856013962577463079213590;
G4[349]<=640'd1176132280945786966052832509236725357663184594433390964886210009340666215068459391734171790504519039649028643755836339382767069494166296160522938442012796604271721695869065053577804215441595713;
G4[350]<=640'd71288131200026132279281215738996065570488773658962090745170423896048561054977384423402775469943090913004255388183931075204418185857773372565048823120351540571807868726859892317761872114760718;
G4[351]<=640'd499016904325030623659882501699550936262968564047308252404441953576482716103455261753264063391392405984786239122792297214045012971211712150321717153507953864399271545401017526921948123708918677;
G4[352]<=640'd267330501486425836681201031182533998113902927661532100747144789852714257126712664552136956176382787935212838788963885607292883863062625277702047704735591996127295584099197691460963224489715861;
G4[353]<=640'd142576269035140797513863510277586725731913226596842707349511868621459037553576593316709397863658823114777274383438951694237700022674436924238647181961858517290427478274074187082517578642494621;
G4[354]<=640'd142576252300128329903392534650768416642426549708121627717874436535380577516180283399586061732776600355038362827550256063723535771670054012570842345107460431211826761417503078952888511185945130;
G4[355]<=640'd142576269300680938073556195283531719645978629169176695818518700403331553401241705100445181228165117208049397991399352082084035942271494533444978793464722425235020762416337133071368999048340268;
G4[356]<=640'd35644067325170108554720830790054341618686335433207568276590663454291817001292680807150044737756496926335483868745504223694863022512919650675371029462397063667868187142460894903252149781728328;
G4[357]<=640'd106932201975517035596866469105475718495885130223272993093866612898338143021001325399219949764422423483143191637697078007775656394440043520107569541108984183203638888423845358739962129323145538;
G4[358]<=640'd534661009877597962060574443234781015984353864504456564179517980166139278981163282509099703186784665759011599750238476263017379814680705728537158929924470580329306996257273455821764075874827681;
G4[359]<=640'd106479689402056084754170771352460129891576021517737245504278158258038436687667399179910979274523076180400585513693791199021194249759077588323400229735071644454122012727560298411718090774682007;
G4[360]<=640'd71233669635995188680603668828874832973487674989476003712133206265027143009818029065269634516020914120350066356169790347113211114233925879361489955648274608806914388814837167101081556382646542;
G4[361]<=640'd110397130727266688016622045039224865971735232330372785685575235679522452705583688988963193138724444741987802276786462046104323233238339319572972075086152883392977303109097052325308409795838276;
G4[362]<=640'd2375900312100378218405855554442456293971881425635766192043881250625307375632357789824456632218128041835186036751650100323691667051874168093557239047660168062326445037615478520008233056102014505;
G4[363]<=640'd508069218983232766809728823652452510487402776904808828103223354711853716725942894782969233498850738969577118820376838466723884240743692466196323010041846504248864397127906338414497731674182148;
G4[364]<=640'd2673592817296823171252796013099797443990742865243164058969397841328843716284920525361939209831830598007369055129592928893458183971793635421129798221071916827485111368222251930866881221433127688;
G4[365]<=640'd108289880976673550568556283646990254786554273107646374370505304494467449979275463127169581646303443145010934958257081503352731017222912271778792764194597114262881314541886433418688193033011491;
G4[366]<=640'd1141865450497895045918305905916946843020742852257230793132238314764658081232103768637173193160580885227431118911931099177725973684392394175939941092769323716358089487975185666244247649184126581;
G4[367]<=640'd2424188491697529068574055289758970461523982941440679379497571184247656458753015688605608365482201560991519126302333151908838890451122716406133506257237981673498664839484228246229057341040492641;
G4[368]<=640'd21275603336633307365040777354346570749342001974680003355507979683916761994834928136584367981041347315571178803328948102444419986052423202452748222734412585794587950883230353195457843341;
G4[369]<=640'd16199768690819136939424503785515530487516520076308209404913605850178271872599843545712032294569765631477309972755922043355975416414424993333981304149157003341359296114893337494857912392;
G4[370]<=640'd1626610897589940525476514228200661642001802845222399402583359688738560154649049151083112090715802517930513581992334734393694219487539161304805943547282357828719080588651981744896221636;
G4[371]<=640'd141213216423281669888747491516659633656902150876828523490923606547886978614191508409377377950512226921411398895487338289529809488973691725801458938654179952311341101510298247511539840;
G4[372]<=640'd31125420027975374321531216839711082647328992305826595478164811361062957513677363651068092241342095675746710244269203781302901017191871260571775884949345691038488226431690426079645831;
G4[373]<=640'd15698618646883213845914545081714373842280405340283227262326773561300722564086573325272892914305931538139540168055162217405924413683981896148179813157754989028406098189366407214858641;
G4[374]<=640'd1251642270552261650429908955186047638579310948310342598630244546619571517593887633009571245300078967586576752135436471677979371238881439303102024510676868255073436511792322329380488;
G4[375]<=640'd663684420682663716023888626811062160939023231528502585896944665948016157646655861853245523065769614854505550629205475962740228324634358693229409783690177621137632274544773017256524;
G4[376]<=640'd461454594240625191089004564653316082097912036265398300753157123123459507874882780958211379488429839800104919663369993846785031345182581844334471157738529090730885073155377013326787;
G4[377]<=640'd24199324811460110424239146874803223477296658831062432069930691274575551990742959864291634652202781316075614006125877614054389317972397079115623981160128712575709952698773388853757;
G4[378]<=640'd6316046225432151389907509664964843904214212884949955045675786161147884633684159663713830109008601234312228063057614878091673937708281096593905598981880748208146797382335791366184;
G4[379]<=640'd103530281912283366725390414586043268613291535275936364817305673609110554264386311513639268821356115488221316729192705291792105876970380931323943395384419975098640229504534106341410;
G4[380]<=640'd2834514798234086169140494586677614339679127331332327578814386439005344636865599097104439162147233329794496794795678419495776740953639784521062571308329368235131144708981849588770;
G4[381]<=640'd8227415066106621454531530875555864725392024909625844075956444809646113419125456276534590752447277103135266632727824537407210043020446055471256565458272676244774293037851479179298;
G4[382]<=640'd56944689744492567447247010158339256268766174977335164540174583165901460928216298367151776668042782442173152433789837112609855541144753601935514589684172033112736198384722903048;
G4[383]<=640'd12737031483679389868018124338485577781997637724841140889821541764611897229906246101210096701062803995012746276819658692259328189675892387631543288496861972035019744208815652864;
G4[384]<=640'd27468893063744592636297556318530339517329511957398606932749001676587093050824701304338564767663818121226538706213435544007548496477881936346806072340240918777716308201292431360;
G4[385]<=640'd5187205623461754731428646321284957602523181398509756098326167411785196965074467371416581375354621337580406589304911404814906671290726266687431987864767800380812997094088376320;
G4[386]<=640'd1251083755947123970194059640362009397966086746894617272157999770007994766240323160123308689219825237948192872444812653072994509080155325880971380674253415421855426033160814592;
G4[387]<=640'd556938551955834693982687264456496189717539542392023343596889815071963528647637928539782063715103132092518320792903233625223129986988043502277444308911708229168870881243320989248671581208576;
G4[388]<=640'd77520960498263255769286589381410756895321910443893699090615336453548978239131459953155159795365232658824707293640632986416686241615427720626756166742176873783949973967077376;
G4[389]<=640'd243660616480677579684649586799958509134085122749171419587534643310411039123090094215453872612400401486560870252177762621378083292304355009554202791694775266951558002987392949967470746140672;
G4[390]<=640'd295873605726537017697930494948728257096494790616466305214476683477334781324946027761676339187551760791107379335741252548607642784709755521931921888269171459261309301444654126859455475744768;
G4[391]<=640'd78319483868789215251900895948478360711824244661272768904945789168065918581841831138838815001385685801740225270696570398914227634986991699938541339893293359179633188745003214965877080326144;
G4[392]<=640'd652662365573243411549064655791435825630079577811031974498823365657320347812199504111965928640720003220695307658651486662673659568943655256170835704940448438433592472408922484594703511584768;
G4[393]<=640'd287171440852227101086500952425170501057467291579354474328978566733963053881359559984692309127838149946231814545672642521283439161381763314660029814523879293299228622239633196425509060214784;
G4[394]<=640'd261064946229297364431051493848780313660889181346483963948028162043179839521298084163613342329810728358218899484918786556094174814248020986561617294234115176375481119080088240829671357284352;
G4[395]<=640'd16747159811483584867591753731593669707597648161062040271232323932144624254131551582327614702622366157481518305398864336725951415754548292513139430467052953973964715065344;
G4[396]<=640'd11318202108679032889451266385590182130383912985986647317318305148726698780785562791991616075597215430147245010162347482313829509322005554588766381431772058810899574554624;
G4[397]<=640'd1903598566255293282926656016533098753955839099296751920129559552612183202158304160570598781925626121799521947848127141567210755364734485202986670410713272250836145715138509957971174227968;
G4[398]<=640'd1903598566255293281957784109791306812410962508801510983710406423310777570794734659503236863456770823237442452590949605582545256125166580999216466042460597147609214095435955531884542296064;
G4[399]<=640'd483167159839152946254246528114660286344628635943694384289378969441728362500724427177376647653614010878225202282971681070388629100394006851126929298830209278589032401469440;
G4[400]<=640'd29830525920830742443819109121744974386104590997379351813506704673190858433074060821245156750907733956572252755133182829053420870143929552058185684737776362146859319296;
G4[401]<=640'd11747564578576323400912357590299760508517374095111235893309935440802772432084193108023201000502713334748318999966913737550402812491042594103818039279980322803664551936;
G4[402]<=640'd745020124376353730166873135837931314530435641176727148991446548117648558245790110139580428282663818161224622639093874093474316301756176169449910954214446292495499264;
G4[403]<=640'd2123483796355242622572621016596219506946743862684794763661429181262518017583058841881978727869516257231808673849590487430486843464176213368397443081510895123160891392;
G4[404]<=640'd781011434732649778410496488980455048736990368886192859169916460324172756697477148609767428229795061225698110049972351765699358246816027650119204556433496836189192192;
G4[405]<=640'd185355687682229939327700270947803963396921513628048803897636010429466502601313989524027857120488685846200702469433200962484865269963803276298489385561832706682126336;
G4[406]<=640'd36230318476817095943765771875018711424381748539017293263597015050760472146019584448689310861665424693685894136253586352544896322536716235956075747660515414640689152;
G4[407]<=640'd17095872419290333401386300611253729616782973038185735789379641662191248895177973165355676607859281954821956144279234292480506702120716097503159451640275189933015040;
G4[408]<=640'd4379411718673045019971496703981511819602670817887849773487270951731675493969951534406593854932315795696944487263370850249217596221547730563282593670023361981317120;
G4[409]<=640'd2748548496054813638758000385432603913599590525851874189730626639513880772732955771322166299998718206387838319448479752637109159442574121310373884563671071946964992;
G4[410]<=640'd105443292033393466994782479344084150401712558197316408808313104478044073080427914448956428731072421384232796188404532754538807073731588570998651499495588357996544;
G4[411]<=640'd108963110190181617342450926305975038303332034198581597686922127902621378687822665360455646534613001423184674029099595371718872187051655382026814680017999646162944;
G4[412]<=640'd27263543959582966209436522637557678587742925269819914955474353391668403865671664642451043479384741882682874965175613860925019371431623479147784897417851283963904;
G4[413]<=640'd5354542279650774614176950093926980762464516861380714350767405930202126461373658884556099551958437840470504410662912100792617802755027259554260766069063396884480;
G4[414]<=640'd768052875391852129794655302613760135388306845562185656801924969318120295964128117444801353957183920965345745269114609149480745755221985738204147894283931746304;
G4[415]<=640'd672750170488212839074620922451162023448184514705989606288240376877646612298214370213209674449173674452939291833598821222867291260581539643340231256312125587456;
G4[416]<=640'd213023570216697318282811613794265535059133618115484370240260569227920686601955131320867087529072932044726002143959209373475780187818591296598181714726918029568;
G4[417]<=640'd32602341970066784625020103985806460510053058589794790938943033443375674425382634087979539551959505064539596136303914111517779644608869129134076258208117162240;
G4[418]<=640'd12457526013783672322559558143543383195256403701662277819359673418173925409813500402936714087571057739454706889526616256134228693801128301586113011457619656704;
G4[419]<=640'd2519829903033366555207555700250209242611676464458172234782289467070229634173495616651784610755579582324601828269122177083598209164669707616034542200498946048;
G4[420]<=640'd1045808999352524064326127587748238761429090563193629372975284797304159207333839524454782178168370916660792475634644958786323077592555563017668099211723276288;
G4[421]<=640'd228613203568426669668179851654983335252401635150541336793516469487423879879358531705940199031193551462327459822979375495256733203626970706103218053847187456;
G4[422]<=640'd29408243517145892475076075347867269267788137947020641438301024922072415838517664888602577256597527928977674742364195291423502451212011479695652982536273920;
G4[423]<=640'd22827195489516828745737442149928633814870444365953796331232668284826380039853260180995772136556989150266073104900457646534026384710235508398510213225775104;
G4[424]<=640'd3428922813750506353537569858464404179802310127295858975914382453991631229465683254230760311920851495331676893714016872491501729225796070468927654371264512;
G4[425]<=640'd2851224724649847214646052431367657558737221747661069783079147077282966516430419803605127934138494802759673560136185200841569160301351943009530517871656960;
G4[426]<=640'd302902113180027475716871310804516856624526481049563403153517107864557305603597868449294846343972878675351525393817307708774988666019550168738188863995904;
G4[427]<=640'd130935636705285239338286684785587639069158814065531452890498012021667402056042750200939159358104031504269718376002483914860983869338575492429363797819392;
G4[428]<=640'd45340576003058991342149036107767688235546099589617510532763941037590189631521168857889023011708919235143274785879236482015568829541156127764263315963904;
G4[429]<=640'd6751380426815462208351912664032775385457847449485510749554060797946239084301562084475187121456104741725039775436130203810504787076011823434009835208704;
G4[430]<=640'd2659542459908572318967850043312675919772991950551070440168228541318590308101763305913554049004214686934571023067152227267717224786473555099271972257792;
G4[431]<=640'd613735764992682296185674696050295309000672380105172194022014973861022783997080972805929201736465163836747230339479659755333437087497984519285814331392;
G4[432]<=640'd172620208981492296510143224881498259110754725416505235779663621569813715432627627810520379944925986113234951696793977203333890810306584708572386426880;
G4[433]<=640'd66730503113231999152009404114068876034205252192051295652280992115205022166005050131137007093073161187104522630081973110266747376598311991168817168384;
G4[434]<=640'd16601461673187246215938983328509217327976364827967683121869150307530000551338334954016208076708238711663216889969689318361882433891340738092960055296;
G4[435]<=640'd2622659000822593554863480960128871706064276281531091443360469382410596409377172323492288970098463591484594238144663962054921530435039472643544711168;
G4[436]<=640'd599374255563001835223434697364690244287309846990504909681922750006277054328763353573885240439208809140286041693948123368094992699151737573506809856;
G4[437]<=640'd199779712890087942192459615293172779003940244208568772204026645530595850932884890304208177071859086795696695155309455865654663227902544874458578944;
G4[438]<=640'd31949145320002251810414594817343003847459392222076792580183042577914214900655818818414350283379156323638731636314024799623717493105910428408479744;
G4[439]<=640'd11706610093798901384145655552874357127700541152224295823184624489455815869917079313501447793987167806496235115265731977741618233285325045704425472;
G4[440]<=640'd2948741488079051131696989549300920264579713970695309974327076087127656829657556946607185809941542229648988157686135168679782100604624770720333824;
G4[441]<=640'd256080352843451852653795427206780234660939395740833168460095102064989799709156891309645381030064265469913007429018319562148175616290633298272256;
G4[442]<=640'd60804559872708354792317217945928300926239460270666208163030596536589610503757447105304796431105789973313327357137630625101170531790183683063808;
G4[443]<=640'd50611234050151699002730515410558527784104208259007735748771330062393162313616557409716246174215153163878555281677080265854830450453735681294336;
G4[444]<=640'd78803704726418006171874296168754016141478037756952908607091661793770611377872294561008834799613866783508431256944640;
G4[445]<=640'd1270714133064343971129527093963571898162096781825370531775789043678265951365152049462376573941033257755165670705725440;
G4[446]<=640'd1566971440295332038038869591770174668221849782225455632366147709033185726320820524508398182758571431408692120572230097205390901203858902038347776;
G4[447]<=640'd21153794784150514999395140829342704729340093015017151453974913051894131968142324062235668914358170301614211115854402989064192;
G4[448]<=640'd105769120229902789671654880153940447387269557791036995820670002718828757774216759150436477020572590529007738366809478501761024;
G4[449]<=640'd1248073834303992834218352177499846022937900600971767054312789627622044536054148601395261668858427263564717380075787743966265344;
G4[450]<=640'd962497656362244724973476549272884374902039883874734162406343758312353247833970724281215380625003922233228979724121524953677824;
G4[451]<=640'd1419607168966040138518167307693383792482361358000437758132219103283987904304989097970175323448752743275640499585343388885182786306048;
G4[452]<=640'd36046229096524580899928849380246349128058229406817331195102246352550694547397246991576951598111356717630188669483142464417298382848;
G4[453]<=640'd623851696559152669785856769581375465907218416099166128936049238762724292537864986825697350261774992221492483714025887710881213579264;
G4[454]<=640'd13863348470605335162090355544050211446465389986334208464876654390306269085976336047654529146378274962415586447084759934360191239168;
G4[455]<=640'd346583711765183813620190273534647003336613301613602522874531954825454991532090914859701532690689085232531678647003944041068904844800;
G4[456]<=640'd47634102832296441461622142397413642652792096015678151040817319912458148615414649538833487005447985527316047245563875884824529438431946736128;
G4[457]<=640'd310539005742503392263323841578453983230443691912630854184481678507379722933718159339190798287655796795539095300580958425695786106880;
G4[458]<=640'd321787390318622330389777931184977197465101717118842651540282283546573485294876009058557184538553144412398440615603353886827151689384499964401758785779020544;
G4[459]<=640'd536312317197703883982960999928403075583218447438381686647503464840874590484491677725705309705881581604521607089481404411748533713255967801503461697825813376;
G4[460]<=640'd1501674488153570922414252019487275994054211391988426447769649278729105868374218653052330395611085595291733064761639164698899579319699596154519076184656982016;
G4[461]<=640'd858099707516326934745504604158345803236713230290546241466667594168962738116972065170320715258375499189018161662922120240470150107637173889578989185426528000;
G4[462]<=640'd4290498537581631790747889298421141770536016341751612764853882571379652473791352390409835713124373773753836962025942455815699706081962999363770465049987519584;
G4[463]<=640'd58350780111110183273901873188593332068820496120784297216497686901865835238317939595734701451629386272171241998962954835099551138897975352358369309754058613728;
G4[464]<=640'd3341631311736019344490509168790733904223082318629744409692523706374659927910685049335346400095887061575604830134967172653259845792909490492222640739254489315261558975643237420551329305080160;
G4[465]<=640'd53674952944743729790990935350249056517713115830413594793914019248830808336080207680404049012238144226230511309371988018493430539698661427393345087700988750394797990594721308580091685766705408;
G4[466]<=640'd522265863792860343908621928371536887475784639347860688904777305241098860776722152142188867072100315432910856311297101831781098867589038255537544593991541048915609857141706883767486499524608;
G4[467]<=640'd418791684576164579972672833486219300068251403174741547562450688643861984146078290512113259369908075063164202330068575819892989415112409162646114044095238041520580133573137732118312168456192;
G4[468]<=640'd3263314034435248753559818495018192752802077807116086245735449718819186028842442404714472594700619763806432237825710137449538595673877979767447538642323756009323366851400973719808990511616;
G4[469]<=640'd2296818939904734499603704203673980547157896592569380904417439099374105720626964548804676055353487729778497299985601848603339533641993895461512776899339329332780125286080358549906651867727003648;
G4[470]<=640'd17804629881027023059192092395689870802214244306481771216976300657987343050335123309733151808442165299117743802898042185156993808621322214884866723022602357166049577501952484280915318431286272;
G4[471]<=640'd285135338229633622725908053163842416103378590834188218391918525541689738552412756505008808041296742047621025647961272943976414818924184381594581735766101397632120613794300466077031156213618560;
G4[472]<=640'd231442785542036358624748140239900543204947447344448511896656661845493322130364170567090047998919944592866576107767192133616241562230213654259342751033832133453288195666897743490833349921216256;
G4[473]<=640'd4425137861363093953023398243794027686279662932491438724129695385767665815708509668112967467046051108290897414050917700066722243973174640625941746759650327768704108339181922426159598505511944320;
G4[474]<=640'd3435462150915356477038430525918236375705544695056588894390239376461924381914692728109980729262625566480327406797274498931354301165314086765765163834963709592474380385125008490977956872813805696;
G4[475]<=640'd3423083302759662132581089490098269509683789980375736115854345601198960300046791361884285265043731899092341047240688805526302129346001541270639988051927768471914077197946416286410386309128389632;
G4[476]<=640'd4505073771387207291176823329627627158803896099808265672985841448926210860776758053989518401361889808670405122895120150178143273580638476657731612181457637167525489691166259773704235362920962048;
G4[477]<=640'd1996137132856141853635860079356895338513280266948321661109912714589571075840264834530615920069157322315755483444826195588789204536473338865928054912966456856282274100436803106844448390773211138;
G4[478]<=640'd998643563294046910009119405913368945133727360199171721477782487497213541357091005619880765189737931698293667605088051148136365128631087172438910935701622798067507279236498980745358435096725019;
G4[479]<=640'd427790125949152152005368619886611144691281805882113493878948099330855068163903803364934693101897661135467739731408515674968713183180603809865500504144772487372851006720027314703820385879392776;
B1[0]<=640'd0;
B1[1]<=640'd0;
B1[2]<=640'd0;
B1[3]<=640'd0;
B1[4]<=640'd0;
B1[5]<=640'd0;
B1[6]<=640'd0;
B1[7]<=640'd0;
B1[8]<=640'd0;
B1[9]<=640'd0;
B1[10]<=640'd0;
B1[11]<=640'd0;
B1[12]<=640'd0;
B1[13]<=640'd0;
B1[14]<=640'd0;
B1[15]<=640'd0;
B1[16]<=640'd0;
B1[17]<=640'd0;
B1[18]<=640'd0;
B1[19]<=640'd0;
B1[20]<=640'd0;
B1[21]<=640'd0;
B1[22]<=640'd0;
B1[23]<=640'd0;
B1[24]<=640'd0;
B1[25]<=640'd0;
B1[26]<=640'd0;
B1[27]<=640'd0;
B1[28]<=640'd0;
B1[29]<=640'd0;
B1[30]<=640'd0;
B1[31]<=640'd0;
B1[32]<=640'd432184316317727476765814107180594002455706216018662415299005541246318057831290728995189006540805689236844046902967438973766410505833415513506355613293998804941839339270454785310584762351484928;
B1[33]<=640'd0;
B1[34]<=640'd3421830463216646413980882478237643315211273621991000936203285305345676791846936416085734854112190941982833818306920983141784070009406609262534395760376290565981628567204450145258199293580279808;
B1[35]<=640'd8911016831293350036421275415735863463291272039286074215957554315348540939336539590523968275125258426843632233720365200848037239317787264465630988430328755738645608177296297149060374010527744;
B1[36]<=640'd8911016831293350036409953528296204348341164383361784948455708905306919926988762470251563033956241069122092658306554949352535591781721314493607081308633677841522742557836217644132033089241088;
B1[37]<=640'd427728807902080801747715516353328220175381850296128668213085038939322191736289270550722963600658550063601553601241770495091063530756673809088312459555963599037764396116762340596431251572785152;
B1[38]<=640'd4491152482971848418350018773766368307872483353120702148115563274434200191710983786707326302496028678652033036407568550867245623290752265482461856543608500061709577932066557945629571361512882176;
B1[39]<=640'd4116889776057527716820863940370128183316443215537096313996948523659989822462480715255358397874835341714800510891708351652588895628156532959370058933543617913917330174413780445153655344632692736;
B1[40]<=640'd3493119685637602503011647814747384772347064941980953578923754351270953312159183075787494930335297190172606535235627953286926404037956276696861199149844536739057758347149298573519847639503339520;
B1[41]<=640'd3493118597866993214396293026980842151195517381439756530179208983395067797816822258906603875894185566902002450999709158167987268376038946421399647683339036237611658386666659525453027809456816128;
B1[42]<=640'd3493118597866993301457079655280276503010001327939758443204583252737234299787853065902069769082110946504332151313658393490129955611275758782922080457342748713341031294929579861178034812820127744;
B1[43]<=640'd3493118597866993277596458853780761831985900110461631844549769072908587913286282232381244983138694919296911979234761361350093050936432149687204636731774105124693718742924102100129359127266721792;
B1[44]<=640'd3493118597870105350952672292121874614500188281089057031078973998856092143047211380520024144962507615338516611692976294528150701693593392515937752645246995954290007799915157923997319304751087616;
B1[45]<=640'd3493118598132562217084069235569208826973957216232649828027388039101534461105636061395762068518710898020126119982071773785071735386934375049890298137946580555922263108067652888833070967635836928;
B1[46]<=640'd3493118598360801814091464326501622372399821596535484903120512531581387818148085970645681106765935652239713813380830095535613226401471537731650009779674996246953176739293553633423933098575265792;
B1[47]<=640'd15560784603270524606087740364428845719116524268442300074893753332590789806737470312653912463970909343603369590784004412189186482686156432927584164203691432118032660539637352649195520;
B1[48]<=640'd956425433090495723230661295613662499049485884813463160695377940269080751918794726504855658789788380652738740528167442998919440757988330660062846755205928267412583112867996783083520;
B1[49]<=640'd8911016832326706534348914427409405078084777406267651070014606774186188021844199939928720354099689679176496872283011835973497192733289040519569418161350745789944237768170724721898725797003264;
B1[50]<=640'd2290200942961628635887277321129949205448335193237819194617113366396476772779209096629094784446000790040808431939732797489707633769088698603226279115954453702460723397859278721760530457943867392;
B1[51]<=640'd3450234329366621322987825738108271114270064286274936192463843861204005953910556609596411446579780739383271983229742939702956661345199908310412049375117165846447364955700356431376271007614500864;
B1[52]<=640'd3441323312538440111359390754860900301457938073133519616402046117440490068018288304190754530769328567889410960698475494622639320773837100193856939151422003722782721143988971943450460764709584896;
B1[53]<=640'd3423501278876351803826558530827910640916303122371587508579187949845970869871917227072664298997879861577234563617555485310689369641957822432526832408401756329746507312149223542589624227781935104;
B1[54]<=640'd8911016832077873719581773014882326530628256929668131224556947080299950080868742144298944073323118809713974328461128136706561689240467246734122502581681302474903855220374732174679881199648768;
B1[55]<=640'd294133172752459642450266801742513682533128896385425630755843210657089999106783976367223378559295623914689379843290286016113435964444702227862095078414018011525510247936725976288585777575624704;
B1[56]<=640'd1078729059987452400202691458407775609321886826142059655889870662917349032234920964759148468057408290183693111391083485506009406687818725204380409278366587083052513327968528779874561165579255808;
B1[57]<=640'd3477245849136261178709963460351904625872523290975143482178723422332754469264375216522677132861200486467829272303457753787520219713793611830132291557917091276716318997923917078436387171560587264;
B1[58]<=640'd3476967379860280602008434953248592669275926129342865271383774263335968591666260634553711103498815409324480124442767983549830762884704290910663294299839331354792753238476439992343235065811042304;
B1[59]<=640'd3478673004175645344665176074467325199005965120355501718744850916130541363085014506569934979536049293824428127239534709596506437471087170229272377245987929532017971773709482210266584433974837248;
B1[60]<=640'd4560247672073875705558405586040134166040799339774773366290286137253986698175922010824222871662174582784280293277792292846363501776179380534260129488808616721078764593656846975178230468941185024;
B1[61]<=640'd2259186427349345101696183609294298175197266245948126300659590175376675759097100948855704358903014286966100838834494269394461603279523988080473651662545608359299691080159534589227897842011471872;
B1[62]<=640'd4558193961163533120950147098170846753006223284446678873092425884959593000507504884229244280526353696925188249173213615892605949326479029978687345883225660351502033319428684641224692410357907456;
B1[63]<=640'd4045601641407182451709278328301898111784284297631378957260758130070092090368352543760932382018333231370300341430281569996640246848723348894773977815611904523295959888441261859095368436717453312;
B1[64]<=640'd570374694521777001979047057380609238644893187687296872951845770016546742252022848528932713775246877554838270699043627619620205475751969944784668728067281718885717375783452963490176327019921408;
B1[65]<=640'd15597273442897654679190440231779648681738258757075500473972049310718091142953842825061798681045414900674981694854956555875186130477501940502068410810995254260065781262911012864;
B1[66]<=640'd6925251241246926953694070588546999572433361782602549920363972404295373704840227309618000072755179887969915034308331595398774728989429206947969885719957560725985701334857285632;
B1[67]<=640'd69747173215415478605061710927518655350054828500922067675157229654056777293043331743973211000553161084894804982795709150975640495876385052692998169378465737522728091748789125120;
B1[68]<=640'd34007930202551873433319096640078959999230657806334900296914288435272735975048531618247283235255622845321004020487497144615570632349155084324022386377863977543121365972174241792;
B1[69]<=640'd17822033662590279933047998299792754701353412122948367871649127788395254650166838663585427475178643273048156086436050535676625421298186546413581001973105578527731464829339042912057535844319232;
B1[70]<=640'd3073327568704796940235804326190026722177281084203559966869104774189639718238771707468071529093419189029881973342972336717172839697305096592467479291494783825382980660734015307776;
B1[71]<=640'd69617319006734518552434035071943067837867575904880798982487054339874774440694298581157184383630358364099059654418946448133812234783411225189216105705982601991156100492098690258943262851072;
B1[72]<=640'd35678875984670700142831833459744459322251769629945093947089821240657595297412667743350080813876440562692638780732292017559692592368375849506698960019459234454173892685217688899560194120351744;
B1[73]<=640'd205593396224518143937791044621579557772139381214447730607494704374423124227133071741117036112295833153145094958918223891546638708886154238270241099012963134594558566143908380672;
B1[74]<=640'd8310301489496312344432884706260084711083682167952205879966537717978384665915688769985189322097053616901574774484549935833196127059269224029752683382277149206472241422632818311168;
B1[75]<=640'd499607410975671158802215092458875669247883167204288701346661150068157759198101479184815749334208354226894157219321321878693249456798082442042877511353007725514930725560736808960;
B1[76]<=640'd4046325368099990177229811188024656430409640768827992304940810592250715528538164501851466712601572562730536885000188653603008802556978615620714863433610465001608894859795102695424;
B1[77]<=640'd34808659501181105857596246559410752135641262235781812242199980816416479870276330781881162944141814886396946256217058066136824695086662158957116131379591941718728368521776506910860103385088;
B1[78]<=640'd1978643211784836272484020168157127572304245736933992613756827758082285823281972297824117461978590353968960255158207189817161904402915452448842426734848818175721985564624692445184;
B1[79]<=640'd506532662216918085755902459144097802306544816443961221788439128436891881291037101220160712224654180987133980445118675912854776125132331043732705193760574372094057275197254270976;
B1[80]<=640'd34808659639290402040177818378795359873012082138135202633684965297895566028195328623558254826702637274002171971859581758331759509813308575544249512272694286479059152345518109293480710766592;
B1[81]<=640'd1011086681222051335239334305928305140509103768453915898339221348485649689029701149612345104605449951674261518374107321230236120650002773237105195204602612681134786350863605563392;
B1[82]<=640'd4046325368099990177229821243881428016780418596623981047159707418800242720912399852121332763318354342493209549764914585996842616869492937451995105404472351541772031795132853387264;
B1[83]<=640'd4052261297735344686047266600481931456294161645997679646797351399297256209520125090181547636904849513427732673176369769583170141122416046411077778228630495556541377852554612834304;
B1[84]<=640'd129893969567250931616030955999182389827021761897027149625758563693333024506687909138405361658860703592743646760671441215608015863993825802769447860535043420128427901029702678085632;
B1[85]<=640'd142082411751845523054532520235030603375591458213570427336822431815438576347275168758758076815967852665231574289998591040167234770049652484819501845742638858080474645231387281457152;
B1[86]<=640'd12409864726513388272619229117791052671518465345348528399926469384148433369900686596926643034406662675241608507855193461780269881152689413323309557945848171221563466573715064487936;
B1[87]<=640'd16630448707614466034157649896877041285701739307118983963374371001832452771027417266649645524076140476498943231257192067638378927040066408672592807711215284116765543347750744205819904;
B1[88]<=640'd8911016832124095013405271037298898205151365833520962950340889415332613955984256403787554762235242500976436303819421897075437315589023036528592799353240706677975366387930351862067491472670720;
B1[89]<=640'd572160300265397535241659143985674709184416542193334336574852604251335371123609554646285406152826495830795074913609781435488470538775219630424507495856086777574140220274062248640512;
B1[90]<=640'd23173869296424002423332844209456863117484032782751707659409011618606350138418209587243954955396075642849351898630984602538112502733154537310049875843548584914382539482392667619328;
B1[91]<=640'd4173702503501850797107252526226714489020266528928471734458175303101941920320199310300031461856408920930072010956470367606271257715611124732241480739281759837961919436430558699192320;
B1[92]<=640'd4656145184615288501245668743727638297898149413478340452309590253022056791759568847258462555848853319102119435804670176342432841533802211066111906753319810004340487582470221424754688;
B1[93]<=640'd33702724487134062438288436529263243997266617838073456849605976904540925483078826306564343784645717672159314180401498076475265627238773021660886571131754950652399870830924119914053632;
B1[94]<=640'd490845978833887903787655851155087341725800520351183675832451054356460712240207356425720125436701299254561469055487719209003823193505721948689606278812008684349199679692283945418752;
B1[95]<=640'd1140610154409897395356332789594080134293905657397944476455605037528365744233620461994873608419575297465868063021197257550749425504483153307417139800192192135631818493335782500880973624569233408;
B1[96]<=640'd26733050598396037806320008026860273279172847384051880869425933932121603489796526013328776899245876884257507688303393568079087077817191298920983327256673991006556619467396553044823405567672320;
B1[97]<=640'd33455469521433407201110822461512507799675892034879992723936451361559784718002424190826505228403551258190333988796134842768439075667942183471835086920295037760704911148135586084159488;
B1[98]<=640'd3042287603319922321211211259802170041529188215526252467844377401638676444474589007116816700268848831204006818122909908961233542473166490227346666434665067602730205364285882761216;
B1[99]<=640'd423251604306480934754796056701357307133183151474652521650084554859819926690596018904449429087640843043224353816056298070191582218241908966847674597815422874443948168684648214994878464;
B1[100]<=640'd398450750120372979655178959776169337181590784844788128274643004382627335835534912095147946940959881073467750072834260684955628817508806370904700560950626581092624211357104959165300736;
B1[101]<=640'd265666282832481389120848665700867307805871696942027783184107358397856749058912139262712021041448860929444050023777976447014284721597520090077656318568476135593731525376713985573781504;
B1[102]<=640'd66489599832098110119431943974347037664958359075357329756010134748513779582043213782333144102481120943531486393537167422336931628764532463566092598310329467353659851506571532629442560;
B1[103]<=640'd236594381596129397268504249606727189594412068694992068391265866688084179710562908477525824109176431217916727267302935182439938583947354471108886916182619707892791126927422915189145600;
B1[104]<=640'd6493783355877096094025523940631265632505082920528851541335707946923747736730200341457355623102089252865079671774939550340778986561882459880444485636223279721692415699396102979584;
B1[105]<=640'd3717973476352482119607745708049748800619449915880657837908293784238094086660846537430400281864128039925378267541718181682065991862114481327056587008031018798148359945574871327202869248;
B1[106]<=640'd531139631133346456534021823321167861372683956826976618222460617600725517809039255617544533113884622223608038815778398175993887784063303310659621703690298740983466192861719684838326272;
B1[107]<=640'd232374518088487810660473547071484931178445886034780208363657722789707143814687725950016308329756455240680539143694303873641009535922133731996757520376188537926244118719632089664192512;
B1[108]<=640'd273104525925692518016207701002039687945343561985935003079156858661102528285938494366939199526638742866306340434955311359228276011771338393231698037678608196427343358343301053579597447168;
B1[109]<=640'd324525329060290894915340009758787804269598499297258567395105684054643093587786996741808087603079330082094505905593775730684842887962928402736512144696045979177140119759944589593416826880;
B1[110]<=640'd933649075862527497797283504132797340237109160539255028202424916360241826293408654080412866985318178773593114612939783307426611902751419153213794880900834097922936125263811988284243968;
B1[111]<=640'd4232513984781208288372028115511593145706960480388967969094530725477149649339392586962247923837660635616638509983587730165736905986586761045236798501144824932934939122492515198271750144;
B1[112]<=640'd152328720585867091092243109689997048831990320943615070625918936602229448468920408784636528902565080531845835134018761911942293740702040254131854739337637752759072140850413355148735676416;
B1[113]<=640'd4174416714547847576562133841457221800031560236374392696333238828570565614451182582794594648632479346859934112220911886471224836605122118940487623626685925476442957004720383721472000000;
B1[114]<=640'd52898040681136224638971902377083444544809332683815731398020962919188380118953291823678074318229211298958556484701868912921674605453793901231487249191324721812067250473644615754590453760;
B1[115]<=640'd54823415905095073102960150818179056479540910900924967872069252650884631095560253748750138691601516219768066514812017054969751113254578166708348205038213543498866982430293335216075309056;
B1[116]<=640'd3992135548353302688530214624829833374917058680566830150444000011973890863597883958552744514754524233394740980643553569749952229385974575618600964443328667958159448463394733732632527425236893696;
B1[117]<=640'd2299042563364854692157896510615291548698134326299833734975314137245209329578276195551940176855035729011754918831826863399937225625670037386393819144439958244049568564269427707063087800004902912;
B1[118]<=640'd53466372901373917943634278803231482280286152431964348184003529027957354122112672907836619102796353297982565542518370028172299357208289794388373246473799222425311839142926249236066853783076864;
B1[119]<=640'd862151756100544587906850240265121171783510181968987091858927676374949238721166597262462018711413168400810152732723354115873341915878186375103778864963117391944170068361726579519625771763105792;
B1[120]<=640'd53536806066998183855021776029348779249786308970305871703536266682961979318455084862514437309836768714425839215728180224456604154449057237360662415717220492351403276041826712561473259789352960;
B1[121]<=640'd4045654398277590009325569501890266427908052804726615416936425447695871935339172282571836327224645268162465375490697564714375624460972072152973852037689844563954672013084285402772181714869420032;
B1[122]<=640'd4026719031396395267833502172219983485708293893928514409126059527910639876503364595607304116392526326565704594441246067911527332536573792938990677479276438787673908483227000607881796306528632832;
B1[123]<=640'd1033625739432486752797017796862258974790418851077796605214463173922922758815664938616922645986960357594875517523423318165061122449329920076335018394996274994707143129579270402508030956300926976;
B1[124]<=640'd2281219492974845062267245920222411751710106409625569330193356783124063293040566786187696678242443481866883525852899126263407566530808233329845790962708271480194517112745756037708149659747221504;
B1[125]<=640'd4562440617618045734618751828790521148404017409676876617446755122886186159388687577552932562464651777037948911502051646839694883975779587330490547292188238676544152843867244764721900104668151808;
B1[126]<=640'd4562440617618045944343327048686025788774530936867371943536302368644163523287933082492957540935526376838315665455514492093484781850140452362203138528345124653658189349051726620542265857549533184;
B1[127]<=640'd4562440345671243960480042253324288950095667513993144718206422361746058301086273089640145227784833777011492127173712195055643376093099646239620884552748462507177190015721160345285039519273320448;
B1[128]<=640'd4562440617617527180079661456031898746913126777523752126151216763627029799806105931794641984402885982093261795969453997304740656541987788724725399970213709376637682481457458902166380758542843904;
B1[129]<=640'd4562440617621157966382118828154578761293983499850532982613067776787793588547484869219343240073705883152794090860168997306634449754694433545401325517969927813151027750907830326222331615712903168;
B1[130]<=640'd4562440617616360089994949125046487405755112456030566630471271198255431440528351645538028634369886578156136253114804796180725676987910453936772120888217039203381831615322968360631292835418603520;
B1[131]<=640'd4562440617616230291494917019389595098679598027423445374436471219930233735325288263837349989183063985794507670359291229306943487983970941432252519939848955398098499411077122657848387100462809088;
B1[132]<=640'd4562440617620120485358087647960248704735128768100217624473781293296245498252205813041359546674190913373855223871839376426202443986937910513268428185833846866557407540105360129101678409047605248;
B1[133]<=640'd4562440617620120485403492232255048985621850039782359136798448180064181840066924827181484839589700685128290376410609187343495790941095713562787349659298355304462705752612734560068083997174923264;
B1[134]<=640'd4562440617619601936626545627770561507582200324041313885310421440219649560729615387063824243473379537114696427458017729507855541275721637436593686280495542414047256348756191612010193992797913088;
B1[135]<=640'd4562440617619861154222075529131258517840581263877403876760259173019502416667957823428022480703757208973090735512818712612722810864131858405439686076017939246617511697408634579159478144637861888;
B1[136]<=640'd4562440617621563311213962585254572846374920945828376865879631764597559557516155376358557388714474035578127749271917297928881639899924654315694589528507768754325505598291320952581927820622561280;
B1[137]<=640'd4562440617622065562107732945132884016718940292287908278176691217704410755390956550642093644216054523766095888096459188465487075878901470182698654451265541528571856863173469722077752880254681088;
B1[138]<=640'd4562440617622085712487593200487769241420082654575056126730794253326694584661808671681481812599913252104782629489261824559965833012119202725178409517694167549035051133410213459701267620738105344;
B1[139]<=640'd4562440617622195218641169718684437346552546375629724296536109739453864166920423498975131016291735378621917607567735908873346430504157333074208778640983416638662445434966480190150151284677672960;
B1[140]<=640'd4562440617622154696028192365237577663271233431654226215634264648775334547470598613276272558369676208512286506287711590579356074831483045048923583548205411843033625841323544899375479207453786112;
B1[141]<=640'd4562440617622195218641171605693992914228844633618722135951029592363217047906597286281166020677853208458106412844046869858343127448257806524630313150388262696662156221909440724867666819256680448;
B1[142]<=640'd4562440617622195218641171590957463320479228181210434048706595352485905011026911591363130075627422008276137885292496916294494976346606744161159150656964801262400490837236739210942564441408929792;
B1[143]<=640'd4562440617622179009595980664321491692261708918780950421359881758593316812445105155489220317950353194588899011563170274358932417127047273821306415793772019321777889324739248425372926443178164224;
B1[144]<=640'd4562440617622195218641171605700291318028430847117937823564340103033119262052151741528161198079068738102258718974563916982049999734771683384230099944285843243322518923985959676400021239073079296;
B1[145]<=640'd4562440617622195218641171605700291323177029092215901404668216562844452142266476188184770788140415044359507103276545589167884711591862390108113608370303217938912320542871374288563761180313649152;
B1[146]<=640'd4562440617622195218641171605700290444482928595497863984150278753449789626114143873309584302296827310044009311347374633075880506542970427062789045005198517108243431441639516051161476685614809088;
B1[147]<=640'd4562440617622195218641171605700290446199128010530516412895594957249198266426716761858390949727678401360625113445796048630171094493845429809707352208260930114378874749885631710895374869398028288;
B1[148]<=640'd4562440617622195218641171605700291297434037866726121070650158357835245322095427945071324354186465491479083439644589270478161244261104332719697514141133624441210656314540806559841218472450195456;
B1[149]<=640'd4562440617622195218641171605700291324893228507248559930577738840450683953619230096503885624258118126714181054201977627939417841953140885845436344597541032409195497168432308899123632519698710528;
B1[150]<=640'd4562440617622195218641171605700291321460829677183255073087333569953378280803215820758407785440408795119980044794042154924823854239611388793483419870202750036139279381478820367608494286071398400;
B1[151]<=640'd4562440617622195218641171605700291321460829677183255073075238519306812082261428275405439356482152439012933626803176437468397395180765030041539948749290389282318500942287554647515450131928317952;
B1[152]<=640'd4562440617622195214682919047749864465339014332961471893084440344170447134602154464447260981860810859363509986865449821564194424198717858602567927079470780323083436683180137768922180393214410752;
B1[153]<=640'd4562440617622195214683885182130618779925188170934204890005464351904922798129754412750117674576773738865803085509867580658339275472179337975566333082502745372366724572432895718308632622465548288;
B1[154]<=640'd4544618583959608514610977530447656299944870199767821484329077763244487174450404438463096149086722514482894098804167956337945648216151831377650527419978492835045138078743497244785718885257052160;
B1[155]<=640'd4410953331490208267527565651783564771375377987429528209061010213228794689072239450288104752026933274213120169462502719591560481308166301440347803909508207384457131477885378976433538210031730688;
B1[156]<=640'd4121345284473174391341389754138841929064063648344184301086208696335355290011203270695926365316622368985009718787400549611793387874940272552496661181688713650722538579710343706773636186871169024;
B1[157]<=640'd4393061680508627087782970527298317185860533881516767388220145101486820519297856951173252051054063273120474648612438420598546017711496453491291435010862719407599158859920847873484306748733915136;
B1[158]<=640'd1797310324480472013775999998450177553578595095204226726542024485886907961930145637747163818754697908003129356499110824458645851793065793007205082357478570038968547541492042816594792658266750976;
B1[159]<=640'd4117968844501942144937409526061162388564330336160241661543487151568171223640790682745417823876102527194358443614127109289694312675298853658987833862134146677440032867201685473851028570747437056;
B1[160]<=640'd4331293680237943790985126909213918870740223336467619475852421657326477835724600920238550785969172270580060561283741847934067631810963113820761074051921804023173457728532171277774720340770947072;
B1[161]<=640'd2139183573728461706732834151519215075260066157646183816064514079265306442073450260676659797819595546324215998931894328044591384455533743317485108147225360127282153414725784720721330561968242688;
B1[162]<=640'd1003025664426731710873690226919786671031140700889393193275559067048007953687570550103620273559028804063872871348890634045263388882769513125409849569972088294844890328215671377737306616136466432;
B1[163]<=640'd2600107877251964224057742882559688251968728426180501065113945636037435675948865962543472878910671997737043666924421368863223088894773224423319022484279959179754373792912844351467588094307336192;
B1[164]<=640'd2307675705856956708548107308363747873266895881484646303402503447449111913787679243080404649776558538021513109926263508989123195977915140585080569030810072491500952308461012807302280884235796480;
B1[165]<=640'd2717734631475137564331077254546363688247035357349570184984135172271787427589346219963761757962812912440725659917223151738942432675955118536814296623177814432068442923797806361053010946632450048;
B1[166]<=640'd506675527494301604849872884059098471095403958853651308383466071619030226000839180959384452157471626766642755112100147800701482265376722204011665996217981065906008263837425617831173320637153280;
B1[167]<=640'd2802515579424324821849565642255586690446320369859612673303313045953877502292955130314373723090745149786452426528243898836291234057439666137816928665481365102645637916374434202155693869778337792;
B1[168]<=640'd1774406294515327460852328177740947440231309797084234214062539470643869662628728285757656659605859770241651938204379788418712550151648368715455295939838405442493434538491211915364185207889461248;
B1[169]<=640'd2210071476780285240448707719924809576795896298118346431464907249509004946702512914334218017622101940922512800599284243872148793109686719595277346734937269428478151736290596789637560886898982912;
B1[170]<=640'd1643108018017537268117704322313699253899846761371942031437239296172741317305971859106527540798599358209484777510714841071409883335130752084054629954508128842661704794113213270647127969200340992;
B1[171]<=640'd2440504753662903409034692659049205546111259801585916132048798007643721354073527018082504838217918123792172051933664121463684968762226357110594264849993170992325805844161405278368586339404742656;
B1[172]<=640'd2453871274772672002869956023842968848180398875287739332423539803689244254130711732662588947022397233217544466980537801387099694525592185614747344703040300018918884249203738320632155919605563392;
B1[173]<=640'd231825839012347773388577284368489446699460214646517045160769738399355523086560609474402361948595317746395579217799950059883540187062455996235107763402619651387400811484624532222684434144428032;
B1[174]<=640'd2237083081519741635533191601035396717275868530047760267493715518340324459219384117401234941380751874975796352604619121748827278452269516110768194388513531007036039800402870709202571802915635200;
B1[175]<=640'd1811025074202487759083350550174354569458920637678190897078538331143967401217084020968897040282908805507913617714508010957304355032125647524476742753185573352259728355080483008328801890101886976;
B1[176]<=640'd116678763440126092476681147493162498286780877339314209473837545976703665677058206738812943415952201684703796452391379139501669439281170570093820225075206331208492133779974671480709261587120128;
B1[177]<=640'd1149939827580818524596209871417401909684632153917815614656213363631551250559488745200352457632070452725053408804485916805371079788942364713834072798486608333038268672548924747014648253890166784;
B1[178]<=640'd4041686501199978552041746562476018651853406255100908388201201358345758611071255917797012957531493935636828855846781170226455244987780625742020158167021761173099248149727840586764707163558379520;
B1[179]<=640'd1844579993140237472088528519003410391513580679081550028367561816905008430459557305693346941767184994145123006849170280299239307825736720836567882381041038375011967479864606247763841281754660864;
B1[180]<=640'd2254452297320704754803766974212999276417410275865672988284608765530708769178620972068144173772599674365355949646353771308280171217617940268881906157135776357068834976668048486561059297512390656;
B1[181]<=640'd2263365472182260981640421460136316246364964554630931794063758013870758984911257503239245587380270840089656514552435753685176269869974488979699988446105450602268451546991953094881412359433224192;
B1[182]<=640'd1122783606169611535720280794344849384845406364198754715024666072540070865385173910086361796342194028392443952533018730034325760978543990530523370545243364737621310503622350927290497474507046912;
B1[183]<=640'd139233625386823835859052737994112659790545081695524707545315734416810739455641484432544833121329995214094875119109646603510313551413825860838138521324925888427080514337966992386290546357829632;
B1[184]<=640'd570235316713044249932086961453523949185023878144920686580513370648198168309042822610138496798842053354126679693389162428809417707457784756014417458291300466337685037329450634114105089456078848;
B1[185]<=640'd4562440587849421011920047128373764957934790993218603883634146603436381479429105937430361264247916617681775465682481350246456271412512338409365551030779963449196465458751548472726146522393083904;
B1[186]<=640'd4562440587874318105333333086124839350359450374238989729643262577486513144551822609228376529546853895306787792110791146539590725099159272015799073211410262822564952386525625208176785271228989440;
B1[187]<=640'd4562440480584443556346379150828021627163021891559457856472107024852573716833341269249408417226602109492999263949580883652722117309754483682045479523934554975637085754600968476643724291179806720;
B1[188]<=640'd4562440480584443556346379150828021626519447110921432758550204947752658445539908854260137638961904635011417284129573662300983689749725089899048149526033353489026332040999971646550021284370055168;
B1[189]<=640'd4562440617621157839748951357460663222954121332819716466803710654503467533844272786916062368063170369664562828718531945417682795676808334229263829655392061883521058774350057952082206871879942144;
B1[190]<=640'd4562440617621157839748951357460663222940713524888023983304633348727366712445881087777391605802003042818977028290289823436680316866392453460642139000252944386354193944137131973537511218408849408;
B1[191]<=640'd4562440617621157839748951357460663222935685596913899193667085856963453148857811940323320397450501414008575668675320426790009833099737922929052277498170319393214248964737068763623531037648224256;
B1[192]<=640'd4562440617622065546279644074670337812154139688171592254814043830707024227089818582816794608286456675984587682101361043597417117299111217094430708544831508237315863467791793921749962144142589952;
B1[193]<=640'd4562440617621935873918116543640384299408360058698328362166540165449354721059880121482409709352605101106911484366678557467361897647643342705495099665659496187993789687697491900409430669615169536;
B1[194]<=640'd4562440617622130382460407840185314568528541809362828745397702194012267932553493871786070051675913981201342516417818270903096364361887550848267949769530592397785119121992925503418639144254963712;
B1[195]<=640'd4562440617622162832209081111500183306458343667509881222727411704569335181046864873814713555115610907109204586289297108486908128082412969270907249535016670650843194263182165814967193804143067136;
B1[196]<=640'd4562440617622162801478278728466944949440879176663669819528466994419540009906071393203685192782836353144302513954756741962509402503281534660050900952834304209560544207880837303589518118460850176;
B1[197]<=640'd4562440617622192690893552250387815159799965975118124840372591431741563186711097542048700826540254374167147791930783953762361182120266839555218440077063348849600474963264032542224761628036956160;
B1[198]<=640'd4562440617622195202796567761329532111642442877576174648203798104825231459574596464720774768376571539570315132896096297313099583268158248683323336144039417449431512938436824036468477791020515328;
B1[199]<=640'd4562440617622193192495064587935879267879516710194804584029611909277038747128215140079127271539470129210131869881979318685127249511507024060426859838016934861932998634096398262898163707554037760;
B1[200]<=640'd4562440617622195218633442530654256808204335461132552666209270105986468791627613453972687543483330028341202797863348854998183169202705377716031343121827836533001805711920593446337556192188956672;
B1[201]<=640'd4562440617622195218637307068177274066548585529607354281504813801604887204124465921236596410143250302482718608722926703654137920366563878678931236731071670472388291484350967678215865809003085824;
B1[202]<=640'd4562440617622195218637307068177274066548716465231670127179614329192591077762544283878365165899371413337764573588198706989236989486451612603825782014327662441131142193209364403137947263272222720;
B1[203]<=640'd4562440617622195218639239336938782695721548602987104749848525744932574779936400964833390106111344956956259371365810472167824258416571674011016581969381170170551909171348954244892078604826968064;
B1[204]<=640'd4562440617622195218640205471319537010307827189459290423224440898835300202386920600663131038312561251796659344029539176309476175958603988414823976157886154203262588376721744735478757552962928640;
B1[205]<=640'd4562440617622195218640447004914725588953794532205483951464337260406764866595562307401213612644741747197867711607825109966016742331227573221562576047529153835360480599772879847923142392411062272;
B1[206]<=640'd4562440617622195218640205471319537010307251072712300702261496706605170872977815388705541615373575206841493397814537466496642128198520983256354333006364724405502684850631737987734369256033222656;
B1[207]<=640'd4562440617622195218640688538509914167600337991698667200673719362727019322228253029605920424900328626301989767152845775136798234486024456609066095599381790092859525654965351468396445658821689344;
B1[208]<=640'd4562440617622195218640205471319537010307080856400690102971113248294260861242544873895427289749097904584539290910386891061920190288495299767080531548906603760922278552947143600159180301250068480;
B1[209]<=640'd4562440617622195218641111222301494180231998542810643239868819482682155126456816513794448463625734775724557730065320876991949949417961680567068084236374870784231407861596655154201816612711956480;
B1[210]<=640'd4562440617622195218641050838902697134251501703254072466244387479767973232729793002278339159624592878145334343126670277079354140023112030716035578828356275299287706178011194363488309972530364416;
B1[211]<=640'd4562440617622195218641156509850592917420401184506215685394133271379586457337464418037803875095164910840808845078511106484612242810527096697005407443481909226054080133318859759898936131832512512;
B1[212]<=640'd4562440617622195218641164057775442560501639188623040190350163518336093477747962698823018728333237737801186090953222615685257352915369817645060821019054904855559797642956281876667389657602850816;
B1[213]<=640'd4562440617622195218641165944756655849966415806118374202493898427061615372789355067325023673388552155940722042035562960176110051946481635714486786535486555173687963362337882767739232173284130816;
B1[214]<=640'd4562440617622195218641171436174000195775855393252201337432003139435463959124609379666786377089784065911402857094956602354169587625231882551252129981755634228406608795265761931133070453462007808;
B1[215]<=640'd4562440617622195218641171602201935958256432453193869396207375991710073706962672793738998301331568248108013808146888559152122706572386971166372617454748780696840387522882632590335820684410748928;
B1[216]<=640'd4562440617622195218641171605448352152398783322686306608642193500754900325703167607352655816633617902788827778952455382995462561063678188835740631220715384894791316425751698672551420208779100160;
B1[217]<=640'd4562440617622195218641171605700291324893215413686128381737286602504390961397914130081981623554144100782224030343460016073119212148417887254726809435978266330991110736858462503961919173175541760;
B1[218]<=640'd4562440617622195218641171605700291324893215413686128393645813680970497647306644255753939538532832851780171616227582294084631198140836081779839110110648521468372766414874264151756078072754864128;
B1[219]<=640'd4562440617622195218641171605700291324893176132998833759028630821089810357340379083071211412506639522867694619471417988653318175197462942490324434963866026112449755396330183383614470702896250880;
B1[220]<=640'd4562440617622195218641171605700291324893202320123696928163588463783529177902047673768082396611437529216275806724851656302782327340376573800399215945974648036667212924246286401479143042546925568;
B1[221]<=640'd4562440617622195218641171605700291324893221960517295544755896565821842671855186828546780694017080020574351848672597862777896904877895413976342466166121863468132643448629188847321317500033957888;
B1[222]<=640'd4562440617622195218641171605700291324893215413736082419981905665671354723789264883917763562768465330763613734839215187575588891286050242138489645027612257083850142798812436873089413323467784192;
B1[223]<=640'd4562440617622195218641171605700291324893176133407788749565804614006617544456233275064819494677795890343106580446800091264305117252745335346217801285598556549598195340065746702187653011651690496;
B1[224]<=640'd4562440617622195218641171605700291324893123758798762566917815847259329109660127969277967141260265303703088575002334348707692694357420271939862133759019055637121092904233280648593042766383022080;
B1[225]<=640'd4562440617622195218641171605700291324893176133198625499529495809672542698248550935309859996742997535592411466680527774277220054663816494395780663303203672545863501337587894264066332957138223104;
B1[226]<=640'd4562440617622195218641171605700291324893176133798001221190166318097814660545956105007707702719311173680881308373453481608223371969660225492023959905253338605878340272074761567750975536060432384;
B1[227]<=640'd4562440617622195218641171605700291324893123761945777769562928140763732246375665046764405182966912738183219869201716888661120829792642255411209599674035271821378035089389414235746534560639221760;
B1[228]<=640'd4562440617622195218641171605700291324893123771535789316133656275567998937268615642306697425599829768373970139917632099930692420091181951708932874894276906442522497801085528556511342668657197056;
B1[229]<=640'd4562440617622195218641171605700291324893123784322471378227960455307021190501424830652955417955551602293077046543154742136452400103955749856995988764928016315804025180840437086450111872931987456;
B1[230]<=640'd4562440617622195218641171605700291324893202524710609754953099288206056598140406666909672344490604876153408046511585445206409318765004745629651204234462615983449629711566255034131409744775086080;
B1[231]<=640'd4562440617622195218641171605700291324893202729297522748461966164030412649865353680449800222182154218859118552519947720498568998969385515998661026164880373955954067787644788478680331285923102720;
B1[232]<=640'd4562440617622195218641171605700291324893203138471348735479699915679124753315247707530055977565252904270539564536672271082888359378153484488857705986818057749332308590211945673885532314493059072;
B1[233]<=640'd4562440617622195218641171605700291324893217050381432294082647471735336270611644628258751660590608208258853973105306990949746613276045869581525597255225599879634097763552266279409914197187756040;
B1[234]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721369010246075625358620046339882630023950176211912738146676113408;
B1[235]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721369010246075625358620046339882630023950178508518860126569889792;
B1[236]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721369010246075625358620046339882630023950177401709712070009683968;
B1[237]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721349726989544517475313542794774536072719909780725127008223232000;
B1[238]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721349726989544517475313542794774536072719909739096103852624085504;
B1[239]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721349726989544517475313542794774536072719911509982426691887302664;
B1[240]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721349726989544517475313542794774536072719910336289247409391796224;
B1[241]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721349726989544517475313542794774536072720065840038127202767732740;
B1[242]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721369010246075625358620046339882630023950856454031433228984783360;
B1[243]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721369010442235054589453820209751049499189751641599366128342138880;
B1[244]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721373831452527260791114219965896492462236894343782117174558064640;
B1[245]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375432113469784394708998092199410417173307748731105261966852608;
B1[246]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375431721150925933041450357779493591038777418262918910835949568;
B1[247]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375431794710711894604115558980152161906178223834327997592109088;
B1[248]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375337564624895132829992820939444817910329027106008501562900480;
B1[249]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375337564624895132829992815631609292303131779362685557431076864;
B1[250]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375412889845743134014678563592031482791347871712638523814479872;
B1[251]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375431721156912243747955184021267406455856859465436987306016768;
B1[252]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375431721174871175867478553678459238854119992128369671977107584;
B1[253]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437973828513637172109997825448962730174457268843658115809280;
B1[254]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437973924294608476228054069001845283609904969866499319660544;
B1[255]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722209636976635814867597483968790678915516480;
B1[256]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722212146890435441423892139727125256694138880;
B1[257]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722190453930915355649653048740834245058035712;
B1[258]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721369010246075625358611635920986269330149181821092851243372515328;
B1[259]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721351434361216542652481304938593495769746085985368626581333873536;
B1[260]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704720861224101191519818229546844721392433205131228372900286510202880;
B1[261]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721169756205689245951133591608887150825755647823173378537647801344;
B1[262]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721373755734987577689277495660168649019273898697653419093853749256;
B1[263]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722091863585872859986449129249041156019396864;
B1[264]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721413913332049463501970196770344528387244032;
B1[265]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722068414875162995573502772267230413061242880;
B1[266]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721412412902800830447866511634718320992714800;
B1[267]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721377023373225991757952142994251783528776192;
B1[268]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722052861430887653055835642227685124196598784;
B1[269]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722073299659686971507591584060256904795469840;
B1[270]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721732977395157882883157339526808315456667656;
B1[271]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722153590778358448945436933183355354544751104;
B1[272]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722196793489465536994765492761694681628295728;
B1[273]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721797337807636216704318855856515460341469448;
B1[274]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721797321343267372668551946970494698394327302;
B1[275]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319717962836135743248312694503691310921691465984;
B1[276]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319714478712101575149515249745107569425873274912;
B1[277]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721146125378138133998989579162901993964581120;
B1[278]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319719226238242912209346154070112096978311911436;
B1[279]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319713741892756525228608247528325730683699920896;
B1[280]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720795221313215625497653646944557066633814016;
B1[281]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319720088134996188306355994046351416337036086785;
B1[282]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319709810687813596590208622738808719634230953984;
B1[283]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319721939767642160088171999855284216894366696448;
B1[284]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319690757910865643892001221987746979254951219744;
B1[285]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319654659428662546437368544833620256177212510596;
B1[286]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319688624771940454280747604617400916958064427264;
B1[287]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319331881936713922586563328711290302939418071056;
B1[288]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319531159949540157435911695929237296182135357552;
B1[289]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319437771857844478025605186063027167398666986496;
B1[290]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661316738420880166526274583982908816170689584236296;
B1[291]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319650585273083959274818769323629417774665760876;
B1[292]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661318617348908045447713449264576553609377056043556;
B1[293]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319416297667051014686559958070954309662497845776;
B1[294]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661318704922065903000412518292976730332118734881346;
B1[295]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319414338663143747287136539633439805657724754112;
B1[296]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319567535991832049396271877039595166187027701832;
B1[297]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661318205946097512041176566805151062907200153865004;
B1[298]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319683579889485405061004691633964455240406145300;
B1[299]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375262239404070492241295385728053645730349478630634246828464384;
B1[300]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721368817219066999353069650917783941209508512854702344707101950336;
B1[301]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721324224693666926654706236782539223179234707533121809085361570192;
B1[302]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704720964269688592477251328415117778739998112197671589133752332726308;
B1[303]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167191025172294363056130819572590027677199425114547971540671985148979541439869473292871784393092621222933287528590413926916;
B1[304]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167169589369856211060132125658996952977415586129277932639742716131930721296210306291682279182124449268998239311828922933320;
B1[305]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275166564356101823540532842225424770497044836558015184692855440903757549450232097112615752830404406523492167025537725730674690;
B1[306]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275162046659995200990160362390241040177706380400701749463883502404046517939482583351517322868870369208280768877478075026151434;
B1[307]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275146560725911869246362435632784721334034252741254714052172290288740141993334133783639778189684998321544597272357575561615364;
B1[308]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275084615768097110922103789780506332229844815897066393429026638002837419167257493736220538075837791420436448808729997787842562;
B1[309]<=640'd4562440617622195218641171605700291324893228507248559930579192517899258971650136356209455495462591960558218757265095525742199718536452927590181844680975772647544363859296258823473779090797387872;
B1[310]<=640'd4562440617622195218641171605700291324893228507248559930579192517899256079843124823261392036257804444862403539381907702468560071850007611891699771371370863820200010400224747856470986381662625841;
B1[311]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274999362435315665788989734895482824161798750153488128567657645492500086398677297896894626165921035750988001377030386647603248;
B1[312]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274831519975830206530143432167614869625177351406418683371645088922494159853931256434331607424732436005692156812179329083508736;
B1[313]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275164665514298866477673275029453287730956728745395043067638184056511247277253051407084066217116172716500322536083453250379910;
B1[314]<=640'd4562440617622195218641171605700291324893228507248559930579192517899105936880667082864654499515758239613992520898751534633452819506120404103375810988235557967582606238611162738252841164803408070;
B1[315]<=640'd4562440617622195218641171605700291324893228507248559930579192517888444426221065122830080439928733660744966757375171639427768380155850703059572455995181498617640683635928804284270494615416881216;
B1[316]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167203633929712779030541121271131995702994588457729675363597734467792955114791563142115931991844266635839462622254945559040;
B1[317]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275156798982565468062559301911209403971564652009235054277801030339124901006146899782570500285094026850967888879993684328988672;
B1[318]<=640'd4420769373468429848921707735192477408173292593975689760615681519761991458561939796321717350661851357999311259910150913615431887128292625879253121987289353276026027784132289873481618496998883392;
B1[319]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167199851337117920447973821031424318973475037550086774283902726507208719367956022906394107022124472380286288361377008714240;
B1[320]<=640'd4562440617622195218641171605700291324893228507248559930579192517899259301857230803250687913673824572932863829542079171922810341709063111905329479624112829197388109410988319150727217346683867696;
B1[321]<=640'd4562440617622195218641171605700291324893228507248559930579192517899254594383551013760071075895954314720492475927154637228379333464511504377644285854430783497521736864407575065173508879177756689;
B1[322]<=640'd4562440617622195218641171605700291324893228507248559930579192517899269881262481633913813892224078835488241435835866791392460179383235434091458005893267553560725817230469320181349476472309162057;
B1[323]<=640'd4562440617622195218641171605700291324893228507248559930579192517899273865714391176358875678020734973198110586926135312311483284315901027097693248492504620342178640951337427935881714917755328128;
B1[324]<=640'd4562440617622195218641171605700291324893228507248559930579192517899274588744357040693280781678103134041435399198244355378669603750544211690948383577429425075595329362272465379626724413438707728;
B1[325]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167203633929712774317978199682645823927006545127020780060484130861039699046960075098447522689188349638410673159419803738150;
B1[326]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167206155658109343564647785541212233118290069304053742027676545184811606734601782770261221955572529652843292534822427432450;
B1[327]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167207416522307628187982578470495437713931831856107009254041757031167243630553916070280769568659802865540502495996103116300;
B1[328]<=640'd4134711809720114416893561767665889013184488334694007437087393219346218120280381555130610633065994251523085545381349908051948686656090218937897347703113019802170018780445797087895748641921959944;
B1[329]<=640'd4562440617622195218611104446604873409104058449227416206776707752844395182247514861114685052301882630477340648171001698395766194825184447717197816957503708209812703438653399110150692552875452544;
B1[330]<=640'd4562440617622195218641171605656764333931023081480426793310236013230871946382859347833006640866105901307058289375933915898497297391591437026509583694269594167932347688606694998428846544237126352;
B1[331]<=640'd2281220308809022851536145306370889458514768673048773742173475040497058992447423149903218660901269342490994276141460964088544863101663409723420453785664842562935962924457545727096625066403713688;
B1[332]<=640'd4562440617622195155332316016593216506132599113563423689286923949253327384927489354309555479164062401286355623240958627141800902483602318124708630622653728142881845022998730963979586003421127200;
B1[333]<=640'd4553529600790901868604763067407907943399296420320340086964780032512753145397722938483118013043651415405590639622503460506382782359265747359302022845050761253898691953256558467898535201608066048;
B1[334]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386496811922121795797261631620908423813569955043579402401900104321663531238746901771678587976921176903598941151760;
B1[335]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912669110804870945741158080443046253140485847962279405209118252553297978217367604839232474313230730394363952;
B1[336]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912768638641632450122135255144700805370902237049677079382274467636217545875483673396066448909198568755316736;
B1[337]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317097993438044868240879704678705881642028395974590576766549456953051767685416155433337423157419968522;
B1[338]<=640'd4562440107729722114544756863695613034523346270839166912628546246432902494821259920087759781714670769813880093421458428484122061432752409379333800760581676874354840565225583513780119731154588241;
B1[339]<=640'd4562440566632947908231530131499823495856240283607620628784127890752637899969935639864097508357738625201731809613572271289437398789690679370932031753809573329424862747276977170988939714247008289;
B1[340]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811264877248363179068390145766086369881079252886524068570977803145591763397333577766259754731481952690724;
B1[341]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811186136347165613105384225701820685781826819870106894073289794005773768863421199402212794947056057985040;
B1[342]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811186136326045846903679602349569593669067636115368279764902928533793137349107173914302164192056387438604;
B1[343]<=640'd285152487612139890755431751155800378768838558062095693866134905222067430711800590014804247616500421291262828299110951174912218067428011422676382119983142710165475676025356865296467224562898944;
B1[344]<=640'd71288109155723145086447569238833137432962583605289098017767569518857540868264710843247236061423981381548847474122262816292593881038386495219203900655231110812174938294487246743085838971711552;
B1[345]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817676646512415206637446503220078003696802631854321632899726631467575249160773436961082856046790509765119982750924800;
B1[346]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243817640572898343660561433780278192642053162622839374912976184157748170131755399795007388750622866223995653798362087456;
B1[347]<=640'd35644067325173400145634153169533525975728347712879374457649941546088087243815638336882219333212146212060901666853213860586832521942418244590819420162146175180468606217556635739246544367386628;
B1[348]<=640'd35644067325173400145634153169533525975728347712879374457649941546087778362348727208599413836472037776802428760410515541355559844993325816122025864732387156774646021118789724922252704151373824;
B1[349]<=640'd71288134650346800291268306339067051951456695425758748915299883091501897400097500968819575951394024463948694313565426861648170182245131376080704648459346415433698329412231772764736096454049824;
B1[350]<=640'd142576269300693600582536612678134103902913390851517497830599766182998506351188740099496604587968700663074548550569395803626160070627279190126645560980279815990135308410931733876911660588863528;
B1[351]<=640'd285152538601387201165073225356268207805826781703034995661199532367350855326459907525966028156484597396596571557638802519823083312365789632001668078683364511299925690622857585298837925198565384;
B1[352]<=640'd285152538601387201165073225356268207804569799709602877183114467524446474356026524232061466489229595634311813878687054670209851463033121881786574481505460185695315991493167910687207939406563328;
B1[353]<=640'd285152538601387201165073225356268207805669658953855980525808052049886870784812207139014995244064284107420919654455433235470241662090837918744271880024525245252718903775867174305311164788115456;
B1[354]<=640'd285152538601387200423082020936954605624319216246590538180470011728691371811853366533589239072905095682027541998336803078547868392797367675109383241058665707350237010389974707523510830987476992;
B1[355]<=640'd285152538601387200179374621577716709302151808470104983719440308812666037527063803810514065919943135231749219879748782621879159923426444521601390903763094481894231221532292576294137308368601088;
B1[356]<=640'd285152538601387201161208452421288143218505559783349741308125200443910750895276153660214171118269933671448346148301503880340227826653347945078301791763926285860760572994294048447801946511769600;
B1[357]<=640'd285152538601387201165073166388103617496280934811639621521858835363099446985157907660303845511279060688793554493523484647022279038679072882432782588410732502857781270904818081013660376330404352;
B1[358]<=640'd285152538601387201165073225356265571723158620654091868025024392586170663779666938194136300642206796866385574208050945629614794078652435560758305677149111685657622081046962805143955115572461568;
B1[359]<=640'd285152538601387201165073131354051346257548530334968338681138938476285191130298818843776413862465819503113223704928671327483919363966535285805864310245466352809053194016231489832080911722610688;
B1[360]<=640'd285152538601387201165073225356268207805820439503269083334907930542244472904501170315777983410489055987749662356996093481666079447829137221521770564747814054471259519100248084662334033881989120;
B1[361]<=640'd285152538601387201165073225356268207805826781703028898496062196446377780768462749803997071474698963194726680616109631121368374291275662479117300301525511769437419246976994514832868487397900288;
B1[362]<=640'd282929135476001018612043555889760440255338843996239580327953264752763531588869521605105191648003436736139200219230308675717642071878306895416301463094674301325534093876730604318877602906374144;
B1[363]<=640'd280698117956349814885887072486723536303436534342790777582519837372208814484796489677758510942820689827713901986762609340822111778492027133260446011004776449801039099873955594703032195561291776;
B1[364]<=640'd276242065655398495498173745202208335613861681094635827816286202123178614942753178882714734695700371335000788745282571374956092749623694509770234613074003962789870647753215992762603934752702464;
B1[365]<=640'd267330521935216271228803306838324054071260780430592692858435617542718333646405646733565047091630518874805483947536172861734761146796031204986345948940437074483233518972261301184314815929122816;
B1[366]<=640'd213864408200144343407941708533906808062108142007753097768458037896250578171709012321121797291232318218080061729414431699490295564315366309437017009916439720535526818259895339406228414940577792;
B1[367]<=640'd142576269898223842501399598703920835848742694821612493483864703202352203821585902425778202708849770141161053080415316823112910475496826713267695197496661442907856310389404734861682830915665920;
B1[368]<=640'd16079372829413847714235580259739912318217088153851647772584721135948712027672873929342593518233982811402894834529967909702667894933721004623874235225974510319976730658587848241840128;
B1[369]<=640'd60783919466030170290708029036124087068484670655150575693857884451870158556074599284253250034562162338874881892656922736392506889547313816130732862603866769541751574022887134199808;
B1[370]<=640'd506532662216918085753981790584784407646247932992322617817011756452466093410462473124010247918581058032662169831964759197929843647441492261191888989002517276213306575420575973376;
B1[371]<=640'd33196330329941969291071601034574870093933763237140603082574504672215572600569495233287604791998215404540125312155073298513764874857214743751065187155990939860643910341628791772676096;
B1[372]<=640'd3215295219150358942357849545235981631400801812494859587598032132605260555330717611805762910138997173538206504064393560931893827919839145472806527020537106180554061301814525952;
B1[373]<=640'd2074757832747215516971931524441995033691617700613809786324259577332472193924938825896590929693654228625760280600262291974009248216541413943144803363613787156661369532971559807877120;
B1[374]<=640'd502480400934278590769093136823907772138518908671749223752934148495299654506536642045791831753748441373809660939977092541234026489125668397375055208845759797475173831382301904207872;
B1[375]<=640'd128659296210645118631589091789828621967601451111833762837156891208596675545571475779856906749851085788117723193416795016835455688005774132314593810842623493840444104082128833085440;
B1[376]<=640'd29315577825811505233429304055463543763200614263799905910299096566799527898284541047873561193124323802175544245048518381252330479279904157909255290953529000708100201488732425027584;
B1[377]<=640'd16082412025387609911467758821183943900204664431809973298926849141635646872843165171130885452396175295197993926482075102553313211667408458736137625584576587723225082893280999374848;
B1[378]<=640'd16193462892581406175669072224567958897889997953078025845932450936856456258505756464239056051608491222754072074772217317729271789609942731459148461593292630337579581116699826454528;
B1[379]<=640'd2026121583809927977890271874556737988534204953726117118415263390471411496882112730884293791555444770156402337488080515393038070656621056692198751513584628234191571370117253038080;
B1[380]<=640'd253264403070663249116191744802311470949573529059754294108026965477826764386954261676741031040973583812351377773623666525932670976967019389564759023037122697822745225803000184832;
B1[381]<=640'd62327140419051616905119852084117723916501322827875931061806090839553764093927321685489856203801043895428996315416334555572860768312696265374212300056151685128786370234693976064;
B1[382]<=640'd31411441238544875088780143511861920902406889162651492890151964106483112857442922646760476264289859187936746049256514854864118422134899694513984672124418067838013119611260633088;
B1[383]<=640'd7852766660822532526720738979383560799070561844199207302164278918229956662667443831093659570295574481224185764931587677059485922366805093412627944182454952322076836007604387840;
B1[384]<=640'd1978402142542335649336816276078601882315812479240849381420115458264235683330772683548002538686642286154873167239529665338048898244983054228460200612677185268394992609408319488;
B1[385]<=640'd989306510273049228737587287351971930309357475860196076862266066277480032974749120417307212413164182209186776550360540793773296680943917284490274266635606035619256180968259584;
B1[386]<=640'd494660801276213118821480403339373527529322450119920006619946917187554502901914114675276282221385448391691064201206109403391966958832902288866877583568274768249018487547101184;
B1[387]<=640'd61832600367418746030366543317883964367155334095568318680866816935542417578309340489052939564106282800559740738122918272809970609054708087488497476119630553152997034754572288;
B1[388]<=640'd15458150092068497877664413599186509937366448810542335028421177159767082644153382636402154944227318575409496089395401094783547607456893232118364751450849965454283578997211136;
B1[389]<=640'd966120513541436498881514731090623656485258552107877730675785991692322877439951031894294256688135784001636748785745045397676392748369552013689548003807894054738889556361216;
B1[390]<=640'd241533591702030197420808011953438039853280764537423643934488145266423705626629059686563553829503234989273230511230035131505615897493584327875469774917643813164180565917696;
B1[391]<=640'd784984184362798223694259455917321396751829131590668283695752078790084006387615992015189553663827843109916014082788157996089496585054556300869551922665477305140527212003328;
B1[392]<=640'd241533595188578417771938721041257086685391253934745512439781817299954637600103569574227691621578583139997708073571190297586139231842890029338497888541927764441772893143040;
B1[393]<=640'd60383391204403844223693808079194219715042613325616649428780475099529920365747734095442870100612724539791425831875153106664355466868218392635744027997455845555255954636800;
B1[394]<=640'd3773645728091004208056949784827764523180490349462953655457142638690932974360276145564313240626266342333073889282371199061341891919691603473263960709190036125467516338176;
B1[395]<=640'd471745302883153640582922563184931721166190595945259971617364522664516103500958100114356601310213807038459409897413760131052814533480253777976630272621424481416603762688;
B1[396]<=640'd58968162887823231466104543804922368292889527754174562775233216983663451250053683199685826048275154334138370112344195450013188521516050825650473627703393986589770121216;
B1[397]<=640'd457003262376013634324587295455236096757087760955207211307671103646545374286994844862237595329897168016102464400562591538496010415778811361764682240132580905972326727680;
B1[398]<=640'd235872651537630146900871530123519873553698641473472151894064566232839119432693767543874527371072091041679300922491792195639973290660067561322795567228757585483710595072;
B1[399]<=640'd29482281545498220938700669745608152637400297407047461852954003977418348663021537488364249297953915740916023728025428235797631244986686092185915135677425145518955167744;
B1[400]<=640'd3685510180489577798115940572444395083396047899115312951182040483968880252318112230612393919577768072571806764988899666195489324897844565968107523701047205513226354688;
B1[401]<=640'd1842755090244891601753755241170376335587708240984327448597851218061589974506197589896672054253509150409311175072421812379094871376589615547971985080669476476648685568;
B1[402]<=640'd1842755090244893232030829506286502699656123001358163252316796689805147418288323034743049871084643637143360003193338187687814649993594646451773898906272442923786174464;
B1[403]<=640'd449891379454319638277980831905278245597310273016628941479589117564257713086445405792031149802611993133039861637892265026001339380094179336227907864903564646774996992;
B1[404]<=640'd230317146562379342178275854556463282833835158254555781609006608366797137776794926202497525272142152827934094541356694795648215721091207106241537455722087962655064064;
B1[405]<=640'd57583459737011212996281467089024869103202430497929822821301095037397884012082281098357120772250556303634211533489019839042535127466091081900648785371017726297899008;
B1[406]<=640'd7198262071269107819253384835201429022560335725055719248228534841211926846078429070614454881237037526621997205692992655523377313535160084182159080377237679951052800;
B1[407]<=640'd899782758908639276540767437485807223954365305720449284497787012374305353954297873723628082356282172856324655620384606654568490243930588147460800655069881082839040;
B1[408]<=640'd337418534590739728710742614420778137765525257917398884720522671806532562508895408486116306398662696867539684412132752882603442155141935813332423276269041705025536;
B1[409]<=640'd217916133769172030523909576368966610509853666758105784612236444252593040302564126698059848194871781839133659344536714425340885713673690273258548819668829095329792;
B1[410]<=640'd56236419184585692705175068244103676972899477805896077674173850476109503091098269445044398043546907703676171473612373627996380017514562345596464411703352343134208;
B1[411]<=640'd28118211215894977212086204959341587437247727786923544799901070393784119828507134345338913061822771956334335798075026381944667252349004666612165974955803109490688;
B1[412]<=640'd7029552803973744348141326138385557602354509899703963649705360814268134132140002289601214688063379327126900839421216799985852747048779859735128864636732386050048;
B1[413]<=640'd878694100496718043517683296603990798251341319582166598904449514297364226528982440293636149227637598018294285205900058133136375981021545434368262424958171348992;
B1[414]<=640'd439347050229527268738344821335307258576521541636041144365118485341487774161371173866248048899836974545357775251521682016957480063979083128393445147283545915392;
B1[415]<=640'd219606851246595444108547176915098115199817279473055561211941085219434614103647933454500729761172613480157407335217337165708915741063983340333368065400172969984;
B1[416]<=640'd54906649244519264953884212067502499147337943185668288313519237007706209614780853209872495678247298481605410896976755862262161032496293439242166019582389649408;
B1[417]<=640'd13729595320261219429963801581180184558049470615461769858100723420424411434325511777414988831758372824046199367489690936845560274146735394221163278549617999872;
B1[418]<=640'd3432398830065304857490950399194112896869689671385969171327869289863404726552735478676101995466402017063077913544065185525439948486912329752938080094417584128;
B1[419]<=640'd214524926779280487115521306569308738744806242901587575900865259197299078858461262974468400027009657548608197026197210745335797069810451245551030424477630464;
B1[420]<=640'd214315682429633921077275074255328750195985036989507351119297805943245597954537659954723462565880118201434537313572307168241293146443842008487739086193295360;
B1[421]<=640'd107213362580422334668542001793610643267451031560179527276294360099076116401347714280042559145374667933501032572182199791706683382671753294088782755026436096;
B1[422]<=640'd53631231719770388398296099949500420539280034119815051694716958121037246964967674040233944092627153913807538044483600495277644083775616204910943778574958592;
B1[423]<=640'd6703903964971298549241883445050476903168332763741562834052227787882941180994027372272069407988288322112225293992334424221962188333231132804368168919236608;
B1[424]<=640'd837987995600072240742700831535969997489572349010469920885193435254654656786106125991394634993392880122482346856869254906567115988175192158321917447634944;
B1[425]<=640'd209496998905353079680844139243123721659438327624157031699709270586021335910774829105577852773304478554990416000873657089364012459660234775017844149059584;
B1[426]<=640'd104748499452676539840422070129252844860629195360968018362396195878598684523884988204030615995845018176413139354752598611174828787160782010619709116907520;
B1[427]<=640'd52374249726338269920211035148911058451071181316809237811381466822352293451711035528045681796055453520869632724054718135445826954096348069602587209367552;
B1[428]<=640'd13093562431584567480052758787310395348002369899548924365003882267788893423067041564638786994958227692740450048599500718780348869866241066401218420539392;
B1[429]<=640'd1636693938183080171759993618965011541290234084600513109970837182384525079250016080743664941435685946077036258299675711987537156398164933394237661118464;
B1[430]<=640'd409173137007357214792425770461873777481671383235688840260690366513737418462277457537962966439231765897678945257964198368389524625090256587086725382144;
B1[431]<=640'd204586912993508866870276647438889912179206371221606599555142886757231222589404629443399500339013031772890343556894444085780246027990626426363232387072;
B1[432]<=640'd51146728248377216718956088993241581432972353973296503649153462084738083898500210634717317598969814337604190330442080290757968668830697580166058606592;
B1[433]<=640'd12786682062094304179739022232574810163650989275108368457895011911987876299571971877367498945822882137735921552836118701138652256895139440832584613888;
B1[434]<=640'd3196670515523576044934752919084327136092168690427698327395617413037648803426562856408012351913850833222279476711478622983799336730743104060207923200;
B1[435]<=640'd399571620714902152385797083330363208460095123744138355585870530206696179694593382193112162688689843327734293780399638486568148883437879894896279552;
B1[436]<=640'd24964842654821933924239438094573438598164690667962997558010393687850687467253307981768794680758716585144758048131802329426332126421127557724241920;
B1[437]<=640'd24973988402527915669695224871826453818675311996650141715376652670470372546721480043991986379502951449483366615854628204033896114205731650657058816;
B1[438]<=640'd6243497100630564855879804602378228463434915026473782845935721501164256192094256554131015725807987475423728542778827381490883712729800135843774464;
B1[439]<=640'd3121748549589153507085990339243842497860593608311329790171838899343881539639126332006908179737300920446063365560644101289181797745753683677675520;
B1[440]<=640'd780436904990606283251194331664673052275698542501007367773009949829479196900369208742741061384736764385615753336344741718685055188749550169882624;
B1[441]<=640'd97507008094739320337495872945962698789480291718066344387950047246599364461731875982456460464034546889712001464927968705245697116325426025725952;
B1[442]<=640'd9145747706003883490375773134159666911372846121088782668532686405152456266073532090196209286318824134257305462269745965514007741247914898358272;
B1[443]<=640'd0;
B1[444]<=640'd0;
B1[445]<=640'd0;
B1[446]<=640'd65334214448820184984967924626899496599552;
B1[447]<=640'd0;
B1[448]<=640'd45593176660108404930896603017233554837679898624;
B1[449]<=640'd45490732611852654880840173311418576427011801088;
B1[450]<=640'd8647113950730249123130474760219402173943906304;
B1[451]<=640'd0;
B1[452]<=640'd452312848583266388373324160190187140051835877600158453279131187530910662656;
B1[453]<=640'd0;
B1[454]<=640'd6113897090266627063976058898204267089283694202907969615560704;
B1[455]<=640'd447576932013383009518794189701917600179649766436916944093130522624;
B1[456]<=640'd3242178505544068212720085574841554886571161569203786379808083950217609584050176;
B1[457]<=640'd59285436618827368806579137128181438006925363167447131384070811635761167627976704;
B1[458]<=640'd48140561100416735743598825635184697194664726310334043598498472463408329979330560;
B1[459]<=640'd837153302757004042579428498828134340502019406263988708846325465088;
B1[460]<=640'd421249012885236229817993396757840860687753187094488055648398344192;
B1[461]<=640'd210624529981749622609049562763130767372625653931076944564328595456;
B1[462]<=640'd1759945529056126297618065354769264561795253338643584044225287554911436800;
B1[463]<=640'd3174803530148166943021607615039634791368706239921136882480880557404192768;
B1[464]<=640'd52656070098325018513905604258913285218868469681193094514751832064;
B1[465]<=640'd3290933378700809870669543538898694655536005502682720013685620736;
B1[466]<=640'd411299618761458417299639902067337383738826041714418419289292800;
B1[467]<=640'd0;
B1[468]<=640'd1889284656273576792668776286210069668170201895132790795504250736975989342037378227832666711420114575889594950196641348373591943950455706624279299673374874603703834247168;
B1[469]<=640'd6607890421487510313463905142674537622518142308797478239563824853379612013111671844919897614091985004751303654356996095937188865014969672851218766654391397744708736253952;
B1[470]<=640'd7728636239978652124188309973180089028671267944634739301573744398175949638871102000334130780763501950016855727464506173842826009111444824557649120553612185503286226405294080;
B1[471]<=640'd3957286043040746409397586606880262768063309605959119899564975469922474742280399275969434786445282485660931345976293426902354547100658121557343360614913504383590008911585869824;
B1[472]<=640'd125620100229412392208694534642375853520471731674668148528263737710799950757684943947152768006138989708928940906381016159212817417163486173230207889623080594617001162623555018424320;
B1[473]<=640'd8299031137761602623966044789588735269137760843425640050179866114650298701656561098130023638021922065391122209598499241735539788854033065329669149558284753918891149595924311398416384;
B1[474]<=640'd4491152483519584473442193986591803340011211496723556952698835071856714311695476966527092543770629411658246438809360252610760438743492725507651512650978027339540738556535559941560770277903695872;
B1[475]<=640'd4544618584507344573660645334282429404647971275841456670268712825329634580574967041405628104824046380466852383305014701495803037729910793788987301059992361800802598221131437725086999127051468800;
B1[476]<=640'd4561953296405378072571232183501032740177114459709185459436624836938440244329111417174967485698712638276110245702994020716302009488174142603148514094696914845618541267581383245118581466285998080;
B1[477]<=640'd3734369503450600479135024397432758391954957406466611387305794092064044092817932515566679110038803699059138093371979732224941783291470854937336971279290627619044382984661180421045747712;
B1[478]<=640'd84733107916549849795086394825784045012792085144508325079462779757200131775607482630113940644027711647878792531757649422674726711056083053166851307276870829352201641346142991614719557632;
B1[479]<=640'd16880229334207818971829678044834007697445335460459978638442807354134721617526906409568469450305001628537654090960751044748825923796345605397023460665973934299876495717353814858843160576;
B2[0]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[1]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[2]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[3]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[4]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[5]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[6]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[7]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[8]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[9]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[10]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[11]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[12]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[13]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[14]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[15]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[16]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[17]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[18]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[19]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[20]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[21]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[22]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[23]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[24]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[25]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[26]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[27]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[28]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[29]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[30]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[31]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[32]<=640'd4130256301304467741875357498519697322437522291229897515280186976652957109377386657510723804776565710541798262670626968336922294215542022484746305706428215383310155335089810164772289429895118847;
B2[33]<=640'd4562440617622195218641171605700291324893228507248559930579192517899275167208677386505912811317371399778642309573594407310688704721375437998252661319722214188251994674360264950082874192246603775;
B2[34]<=640'd1140610154405548804660289127462648009681954885257558994375907212553598375361740970420177957205180457795808491266673424168904634711968828735718265559345923622270366107155814804824674898666323967;
B2[35]<=640'd4553529600790901868604750330284555461429937235209273856363234963583926626269340846915388843042246141351798677339874042109840667482057650733787030331291885432513349066182968652933813818236076031;
B2[36]<=640'd4553529600790901868604761652171995120544887342865198145630736808993968247281688624035661248283415158709520216915287852361336169129593716683759054238413580510410471931802428732438742159157362687;
B2[37]<=640'd4134711809720114416893456089346963104717846656952431262366107478959952975472388115955189847716712849715040755972352636815597641190618764189164348860166250589214230278243502609486442940673818623;
B2[38]<=640'd71288134650346800291152831933923017020745154127857782463629243465074975497693599798586508821342721126609273166025856443443081430623172515790804776113714126542416742293707004453302830733721599;
B2[39]<=640'd445550841564667501820307665330163141576785291711463616582243994239285344746196671250554413442536058063841798681886055658099809093218905038882602386178596274334664499946484504929218847613911039;
B2[40]<=640'd1069320931984592715629523790952906552546163565267606351655438166628321855049494310718417880982074209606035774337966454023762300683419161301391462169877677449194236327210966376563026552743264255;
B2[41]<=640'd1069322019755202004244878578719449173697711125808803400399983534504207369391855127599308935423185832876639858573885249142701436345336491576853013636383177950640336287693605424629846382789787647;
B2[42]<=640'd1069322019755201917184091950420014821883227179308801487374609265162040867420824320603843042235260453274310158259936013820558749110099679215330580862379465474910963379430685088904839379426476031;
B2[43]<=640'd1069322019755201941044712751919529492907328396786928086029423444990687253922395154124667828178676480481730330338833045960595653784943288311048024587948109063558275931436162849953515064979881983;
B2[44]<=640'd1069322019752089867688499313578416710393040226159502899500218519043183024161466005985888666354863784440125697880618112782538003027782045482314908674475218233961986874445107026085554887495516159;
B2[45]<=640'd1069322019489633001557102370131082497919271291015910102551804478797740706103041325110150742798660501758516189591522633525616969334441062948362363181775633632329731566292612061249803224610766847;
B2[46]<=640'd1069322019261393404549707279198668952493406910713075027458679986317887349060591415860231704551435747538928496192764311775075478319903900266602651540047217941298817935066711316658941093671337983;
B2[47]<=640'd4562440617606634434037901081094203584528799661529443406310750217824381413876086596699175341004717487314671400229991037719904700309186251515566504886794630024048303242242232289543236839597408255;
B2[48]<=640'd4562440617621238793208081109977060663597614844749510444694379054738579789268408305753994016590866544119852521192941668570160537278376518557494672989062151341496788746092852366970006195463520255;
B2[49]<=640'd4553529600789868512106822691272881919815143729842292279509177911125088979186833186565984090963271710099465812701311395474715207528642148957733091901560863442462050436592094225360975466449600511;
B2[50]<=640'd2272239674660566582753894284570342119444893314010740735962079151502798394429468289876818026871370609737833877633861609820981070952286739395026382203767760485791271276500986228322343734302736383;
B2[51]<=640'd1112206288255573895653345867592020210623164220973623738115348656695269213298120776909501364737590660395370326343851467607732043376175529687840611944605048341804629718659908518706603184632102911;
B2[52]<=640'd1121117305083755107281780850839391023435290434115040314177146400458785099190389082315158280548042831889231348875118912688049383947538337804395722168300210465469273530371293006632413427537018879;
B2[53]<=640'd1138939338745843414814613074872380683976925384876972422000004568053304297336760159433248512319491538201407745956038921999999335079417615565725828911320457858505487362211041407493249964464668671;
B2[54]<=640'd4553529600790117344921589832685408998362600250318891799354635570818975217127808644361613867244048280968928335245133279173982143032134970751518538817140532885777090819139890217908194311046955007;
B2[55]<=640'd4268307444869735576190904803957777642360099610863134299823349307242185168101893410138689432758075775863952929730304121294575268756930735770390566241308196176726484426423538973794288414670979071;
B2[56]<=640'd3483711557634742818438480147292515715571341681106500274689321854981926134973756421746764343259963109594949198182510921804679298033556712793872252041355627105199481346391736170208313026667347967;
B2[57]<=640'd1085194768485934039931208145348386699020705216273416448400469095566520697944302169983235678456170913310813037270136653523168485007581826168120369761805122911535675676436347871646487020686016511;
B2[58]<=640'd1085473237761914616632736652451698655617302377905694659195418254563306575542416751952201707818555990454162185130826423760857941836671147087589367019882882833459241435883824957739639126435561471;
B2[59]<=640'd1083767613446549873975995531232966125887263386893058211834341601768733804123662879935977831781322105954214182334059697714182267250288267768980284073734284656234022900650782739816289758271766527;
B2[60]<=640'd2192945548319513082766019660157158852429167473786564288906380645288469032755375681689939655196816994362016295802114464325202945196057463992531830913597467173230080703417974904643723305418751;
B2[61]<=640'd2303254190272850116944987996405993149695962261300433629919602342522599408111576437650208452414357112812541470739100137916227101441851449917779009657176605828952303594200730360854976350235131903;
B2[62]<=640'd4246656458662097691024507529444571887005222801881057486766632939682166701172502276668530791017702853454060400380791418082755394896408019565315436496553836749961354931580308858181781888696319;
B2[63]<=640'd516838976215012766931893277398393213108944209617180973318434387829183076840324842744980429299038168408341968143312837314048457872652089103478683504110309664956034785919003090987505755529150463;
B2[64]<=640'd3992065923100418216662124548319682086248335319561263057627346747882728424956654537976980097542124522223804038874550779691068499245623468053467992591654932469366277298576811986592697865226682367;
B2[65]<=640'd4562440617622195203043898162802636645702788275468911248840933760823774693236628075787821668363528574716843628528179506635707009866418882123066530842220273686183583863365010690017092929335590911;
B2[66]<=640'd4562440617622195211715920364453364371199157918701560358145830735296725246844704982210539106477144090160642236818414519340773670413043842599477932330293007240282108954402704224097172857389318143;
B2[67]<=640'd4562440617622195148893998390284812719831517579729904580524364016977207492051447732449135518274039655805431309020433322415883721925666287022612165443337161495253825295894527427354782443457478655;
B2[68]<=640'd4562440617622195184633241403148417891574131867169599931348534711564374870294388951233176836268839781531359074317971561989684684233878293382682028970567129864229608296496287406961508220072361983;
B2[69]<=640'd4544618583959604938708123607400498570191875095125611562707543390110879912558510547842327383842192756505594153487158356775012079300077251451839080317749108609724263209530925907170816656402284543;
B2[70]<=640'd4562440617622192145313602900903351089088902317221837753298108314339308298103903196866194572545663931707113216154405377428715361749038720825412964014625621720772703179576439567102213458231295999;
B2[71]<=640'd4562371000303188484122619171665219381825390639672655049780210030844935292434236692207331654132987769420278210513939988364240570909140654587027472103616508205650003518259772851392615248983752703;
B2[72]<=640'd4526761741637524518498339772240546865570976737618614836632102696658617571911264718762562730503494959215949670792862115293129012129007062148745962359702754953797820781675047261183313998126252031;
B2[73]<=640'd4562440617622195013047775381182147387102183885669002158439811303451544559713973012082788584184299658661606197277761254165593745803151546451613952433567975918010895661397130355524308048338223103;
B2[74]<=640'd4562440617622186908339682109387946892008522247163848846897024565693395200670959408121246895628601414589320212519977505735914220171439604802125602050498184435568612397211058477841451559428292607;
B2[75]<=640'd4562440617622194719033760630029132522678136048372890682696025313610573820547527318348153613215892214962892975365240180416531485400053559305003204521639772145374483321352539435152148631509794815;
B2[76]<=640'd4562440617622191172315803505710114095082040482592129520938423689906970226398085135790384273152869548311929708001031676773803704532721834989450104341106593473388561063895263341188014397143908351;
B2[77]<=640'd4562405808962694037535314009453731914141092865986324148766950317918458750728807110175130930154427257963755912627338190252622567896680351336093704203590834596310275945991743173575963332143218687;
B2[78]<=640'd4562440617622193239997959820864018840873060350120987626333455583906661410380919304220089529345073575661180330983240438350433546514185620836348258404269765345825259825542089228097309567554158591;
B2[79]<=640'd4562440617622194712108509388782205568990769363150757624034376073938053378769548949614031520280270179617930084919413420176708259602699525143476536187391170455546800913785892856025598994992332799;
B2[80]<=640'd4562405808962555928239131427881912529533355495166421795376558832933977271642649191177289253062544697141368307401622547728930372961865624689677117070209941493965515615207919431973580711535837183;
B2[81]<=640'd4562440617622194207554490383648956085558922578943419421475424063983376827987328900856223781616221787433537704123642733049170330614054207762132011316948977083056790071747583815296523328641040383;
B2[82]<=640'd4562440617622191172315803505710114095071984625820543150160595893918228007501258586263191898917519278445878991219251914101138939806789441155635791826784762193146590202008723178051079059393216511;
B2[83]<=640'd4562440617622191166379873870355605277626628025317103636417546520219628369857278089249703291192281218231005404724080979578015528351605854828111538903675803110473766043864708408705021637633769471;
B2[84]<=640'd4562440617622065324671604354768675293937229324858732908817295490749649408644984053481406123408232994416983448870001663663928033280159829982388667493919444740391459630940136522181844489568518143;
B2[85]<=640'd4562440617622053136229419760177236792372993476645184339120978947471938344776861947929565536148612641701826341720929175736398706130335270763482611667237394686406252035502184475437642804965146623;
B2[86]<=640'd4562440617622182808776445092312018705664110716195888412113847169370875240739293238072542910630774473135607902910919165702180849527913657728371508630308890878694048826189043386616300477182115839;
B2[87]<=640'd4562440617605564769933557139666133674996351465962858191272073533935900796206844933734885394050721754254566169097095464079431512653737059071212594911049621380540779390243499406735123448040783871;
B2[88]<=640'd4553529600790071123627766334662992426688077141415038967628851628483942553252693130102125256555136157277665873269774985413613267405786414961724068520368973481574019307972334598220806700773933055;
B2[89]<=640'd4562440617621623058340906208165049665749242832539375514036999183562700314604426051134789201762725114372489483077763612235775094939939949527713886100091789680756138587582690809862600129997963263;
B2[90]<=640'd4562440617622172044771875181697867992049019050385442446546409766191615758197058780155774393107784155823686913497951557958790073736772899885749928165184904138376151125775350567543391799578984447;
B2[91]<=640'd4562440617618021516137669754903184072367001792759539664050264046164816991905575444585592612007071368316785900652664335299732234353769166740537050194989972707512712914522303030646443633547411455;
B2[92]<=640'd4562440617617539073456556317199045656149500868950661781165714177446965576955655329714153242470112937222793456254492287874884034545033005156718859108656102281498674864355924462500403970821849087;
B2[93]<=640'd4562440617588492494154037543262002888363965263251293312741119061049669190304136461022833985010807055993996591901435093130287206644900172371013888298061327617120239723707865079251950072332550143;
B2[94]<=640'd4562440617621704372662337717796503669042073419906834130058841334223442716154320925793672603960945679653205608274339845841633217002166434175059155597773524581973182665675915750403181908301185023;
B2[95]<=640'd3421830463212297823284838816106211190599322849850615454123587480370909422975056924511039202897796102312774246552397149759939279216892284690835521519530022052620176181024482449201900567677370367;
B2[96]<=640'd4535707567023799180834851597673431051614055659864508049709766583967153563718880860492584034418125522894384801885291013742609617643558246699331677992465540197245438054892868397038050786678931455;
B2[97]<=640'd4562440617588739749119738198499180502431715999448884038544312525175338715847117601787910387126544894550238758315404073321892569878606998922584719136250379101331699636599560038934738606162444287;
B2[98]<=640'd4562440617622192176353568285777970113681968705078518401390976991646807322831275747829468336728364282961942040724763203303870581811466476764710188153231986841585560009292662219877509906363842559;
B2[99]<=640'd4562440617198943614334690670945495268191871200115376779104539996249190612348857459815316792412921970691001466530370053494632406651183855780010752352874539590436571799916316781398225977251725311;
B2[100]<=640'd4562440617223744468520798626045112365117059170066969145734404389624632162826050050670377899222223452837682428500126657237854444036419809180743854948817513627301368093267640738725769233081303039;
B2[101]<=640'd4562440617356528935808690216579442659192361199442688233637164734715167808810820637447000672054659378737193448644150357286910728274361153276655141229644557869683518538766533424706160206672822271;
B2[102]<=640'd4562440617555705618809073495580859380918881469583601571503835188143265032460163606923869597535038255676161188630062920917151537299038506369488128856156121589941665207006605098576302659617161215;
B2[103]<=640'd4562440617385600837045042208431787075286501317654147861884200449508009300520593206795349902839845575669465878355677680043385769538935499414305306848613327272069374966467473823155451277057458175;
B2[104]<=640'd4562440617622188724857815728604197299369287875982927425496271989047733831500730462758176081117029942423019207484341542231016929781825097219266099437262333743766358451080543257667174796143624191;
B2[105]<=640'd4562440613904221742288689486092545616843479706629110014698534679990981382970583299845066273886971117914514269648216139768970523039309446136138179992665627180220975876211905004508002865043734527;
B2[106]<=640'd4562440617091055587507825149166269501572060645875875973752215899676814549607951868696873555699826866664757687349986368494910306545381550214189358009062592484561695933376798757221154507408277503;
B2[107]<=640'd4562440617389820700552683795039817777821743576070114044544412309535617444418970242691225085367355091448885854332913868166994400847734428462330527587725456667875806136434020831363242102582411263;
B2[108]<=640'd4562440344517669292948653589492590322853540561904997944644189438742416506106149100567418444378171873139899443267253972355377345493099426226914268088024176509643798247016906606781820612649156607;
B2[109]<=640'd4562440293096866158350276690360281566105424237650060633320625122793591112565583798718916069509283796699312227479088501716912974036532550035324258583210069492206015497220145190138284598829776895;
B2[110]<=640'd4562440616688546142778644107903007820760431167011450770039937489696850250848435560212504157236958532793324130800001292697748921413948826095501242166508419307351160576437328824819062203962359807;
B2[111]<=640'd4562440613389681233859963317328263209381635361541599450190224548804744441731527737166520224355123475940981673956955897327100974555638532011665900274485415687107169741425325827590358993974853631;
B2[112]<=640'd4562440465293474632774080513457181634896179675258238986964121891980338564979228917585504026680842497213561777727759273291926792779081697296212407187867474850614241915288124099669519043510927359;
B2[113]<=640'd4562440613447778504093324029138157483436006707216999694204799821566036338638111772054730228522776751146162962713660295089776818250150601393130542379234590561566069197917307945362490470774603775;
B2[114]<=640'd4562440564724154537504946966728388947809783962439227246763461119878312248020297267552620987639297081549431010615037922608819791799700832544458760088234964996927272862293014476438258437656150015;
B2[115]<=640'd4562440562798779313546098502740140506714172027707649029654224645830022516324046290945659062567232708177126089805527892498671649751624324743674494611374009150038451175493282519789538976171294719;
B2[116]<=640'd570305069268892530110956980870457949976169826681729780135192505925384303610793427953168296562847166383901328930040837560736475335400862379651696876393546230092546210965531217450346767009710079;
B2[117]<=640'd2263398054257340526483275095084999776195094180948726195603878380654065837630401190953972634462335670766887390741767543910751479095705400611858842175282255944202426110090837243019786392241700863;
B2[118]<=640'd4508974244720821300697537326897059842612942354816595582395188988871317813086564713598076192214575046480659744031076037282516405364167148203864288073248414965826682835217338700846807338463526911;
B2[119]<=640'd3700288861521650630734321365435170153109718325279572838720264841524325928487510789243450792605958231377832156840871053194815362805497251623148882454759096796307824605998538370563248420483497983;
B2[120]<=640'd4508903811555197034786149829670942545643442198278254058875656251216313187890222301643398374007534631064216470357866227086232100566926380760891998904004993695900591398318438237521400932457250815;
B2[121]<=640'd516786219344605209315602103810024896985175702521944513642767070203403231869505103934076484092726131616176934082896842596313080260403365845278809282032369624297322661275979547310692477377183743;
B2[122]<=640'd535721586225799950807669433480307839184934613320045521453132989988635290705312790898608694924845073212937715132348339399161372184801645059261983840445775400578086191133264342201077885717970943;
B2[123]<=640'd3528814878189708465844153808838032350102809656170763325364729343976352408393012447888990165330411042183766792050171089145627582272045517921917642924725939193544851544780994547574843235945676799;
B2[124]<=640'd2281221124647350156373925685477879573183122097622990600385835734775211874168110600318216133074927917911758783720695281047281138190567204668406870357013942708057477561614508912374724532499382271;
B2[125]<=640'd4149484022419776909770176489211097571683313132437395013089007819989808952980248852719622740693398071542760470993820745595850667762114027533975511707841830493020185360974087578451967;
B2[126]<=640'd4149274297844557014265536118697570381187987042890149255111643920744304012955273793956153601825246139183389520693252822179297829460923615579235534120484076334978558221164490661036031;
B2[127]<=640'd271950951258161129352376002374797560993255415212372770156153216866122404296865767623830444976169361877038863244670101363895069386535177705475371404178048861907941114074804608145716936703;
B2[128]<=640'd4668038561510149668392577980101729724807804427975754272245367402571454711270970223152905468321798490486330752499906119048761396806095965998636791734819736013295652499851984190308351;
B2[129]<=640'd1037252259052777545712563599245007398026947966124741111481578661192517286569857922243512485655122368547313856451369075891972764418953254654127314820665987255939683285628634152304639;
B2[130]<=640'd5835128646222480653803919138116051217993300107921319643843726680325740967884463626062817482312960113911514982360141842675952373048157884407015924589862122840801648876667414446604287;
B2[131]<=640'd5964927146254586310696226213630479825114556142721297969041431883389122668562965473596411914038091041864129929943773792009980721783950106324179260013344795184894821947030120593096703;
B2[132]<=640'd2074733283083957740042620158099739148342306105411224603029668956471573464553407982469484334690537529315982810684817789043011640768041860339287791554436666156657350693738812008300543;
B2[133]<=640'd2074733237679373445242339271378467466200793780744337835093327141752559324428043382004458541822575606158180340468842750110280497104728968668924873849542693302775192306469470314954751;
B2[134]<=640'd2593282014625977929729817311028183207246045268771077679625606479061999442088603644911725912285060244693131264059671546331045421760134456239957492315429220989184660536361712793681919;
B2[135]<=640'd2334064419096076569032807052647243371156053818933344879772750540719563077890366309546019264306179820012041257546576420968691770039937712280571552067429910766697378658445063847149567;
B2[136]<=640'd631907427209020445718478518307561420183064699560753301715609692522010147355422602897364200514560301677109381807064821450783682558071791214445433926489076068943997500946371624042495;
B2[137]<=640'd129656533438660567407308174288214960651652402501300194864411817720835863819167101316876012546421477135218845201628842473967815554006868456672659680137811186795228005121311991922687;
B2[138]<=640'd109506153578405212522083473145852673503803848398264572580582546868714824431012155926600740684943428986266161388540439129218680971461201962652421968170621915723775646566201151193087;
B2[139]<=640'd1887015853978340682131618835634043082778445411000288253887530781808464104474223549965350512181848007942947091088331941092078673403332340776320359457045197682537211625471;
B2[140]<=640'd40522612979240462713661621995075594333714944927869123940619738078773229640252947695191266355803285882816731332629889892392949329077771516802345218368833036720050707394984792817663;
B2[141]<=640'd6298410664383873629837794628162925536058119302080100224746790639518191320535896729547537452345577273117631473622348169333951491589838452450824225215207372989923327;
B2[142]<=640'd14742828004414000326038125881872597165413370156181765795142782735689949391502504424281097491016193728374768693837093510662757412925851503837123525739140309750837673983;
B2[143]<=640'd16209045190941378799632631519588467609509219310759305958354763572231016692493367018205189743298010424132951756287594328164176946245525950194866474105349621016524709947749068439551;
B2[144]<=640'd6864797660130622107014852414866155905156525644977751613238302661676383590599030490328638704986603754614022561375436370944929475750374305273682852953173524479;
B2[145]<=640'd1716199415032658525910975955054823024942201198321142023176956355419135206297048818142803993129513047890139052949418996249339674131488890661519113011932954623;
B2[146]<=640'd880410299911750695946428913764449485541094533513196328509020544089734632998226219774234808198178405010935463616314523697080008563232720748898921397506631794687;
B2[147]<=640'd878694100496718043517683597560650076900781960624647521861589692998418017196127798358680517610227530008188545309111461284073873119924474633239187499322848575487;
B2[148]<=640'd27459190640522438859929034160064029845113249441434588457130905908299558869929005136832527460460271105278555147178588589747041338359819458390241655719796408319;
B2[149]<=640'd1453677448591213589447290002027187059253273064461255371616779371270862768234552152816316722181181779056497505927956050959241672547893247;
B2[150]<=640'd3432398830065304857491858947945896886405461565747505025876962604658662264779552252385864850481764049204769241449519464152112715292881444582474379906175205375;
B2[151]<=640'd3432398830065304857503953998592463084947249111100473454835218960765708682770417969842291309540610407956712712570431824905933493732072710302567424060318285823;
B2[152]<=640'd3958252557950426859554214174287088037494752173728828032606522922058651829456560540415132322708144585746494280522657579395684734240251433865168557991180127181160693799032193023;
B2[153]<=640'd3957286423569672544968040336314355040573728165994352369078922973755795136740597660912839224063726826652349429249196100022686328237219468815885270101927369231774241569781055487;
B2[154]<=640'd17822033662586704030194075252635024948358307480738446250114754654787992758272948042816662230648885295748210769426450972743056505223606620602133899743721353206856595616767705297155306989551615;
B2[155]<=640'd151487286131986951113605953916726553517850519819031721518182304670480478136437936217808059290438125565522140111091687719128223413209136557904857410214006803794863196474885973649335982214873087;
B2[156]<=640'd441095333149020827299781851561449395829164858904375629492983821563919877197474115809986446000749030793632590786193857698895316846435165445756000138033500537529456094649921243309238005375434751;
B2[157]<=640'd169378937113568130858201078401974139032694625731792542359047416412454647910820435332660760263308126658167660961155986712142687009878984506961226308859494780652835814439417076598567443512688639;
B2[158]<=640'd2765130293141723204865171607250113771314633412044333204037168032012367205278531748758748992562673491775512953074483582852042852928309644991047578962243644149283447132868222133488081533979852799;
B2[159]<=640'd444471773120253073703762079639128936328898171088318269035705366331103943567886703760494987441268872584283865959467298020994392046076584339264827457588067510811961807158579476231845621499166719;
B2[160]<=640'd231146937384251427656044696486372454153005170780940454726770860572797331484076466267362025348199129198581748289852559376621072910412324177491587267800410165078536945828093672308153851475656703;
B2[161]<=640'd2423257043893733511908337454181076249633162349602376114514678438633968725135227125829253013497775853454426310641700079266097320265841694680767553172496854060969841259634480229361543630278361087;
B2[162]<=640'd3559414953195463507767481378780504653862087806359166737303633450851267213521106836402292537758342595714769438224703773265425315838605924872842811749750125893407104346144593572345567576110137343;
B2[163]<=640'd1962332740370230994583428723140603072924500081068058865465246881861839491259811423962439932406699402041598642649173038447465615826602213574933638835442255008497620881447420598615286097939267583;
B2[164]<=640'd2254764911765238510093064297336543451626332625763913627176689070450163253420998143425508161540812861757129199647330898321565508743460297413172092288912141696751042365899252142780593308010807295;
B2[165]<=640'd1844705986147057654310094351153927636646193149898989745595057345627487739619331166542151053354558487337916649656371255571746272045420319461438364696544399756183551750562458589029863245614153727;
B2[166]<=640'd4055765090127893613791298721641192853797824548394908622195726446280244941207838205546528359159899773011999554461494259509987222455998715794240995323504233122345986410522839332251700871609450495;
B2[167]<=640'd1759925038197870396791605963444704634446908137388947257275879471945397664915722256191539088226626249992189883045350508474397470663935771860435732654240849085606356757985830747927180322468265983;
B2[168]<=640'd2788034323106867757788843427959343884661918710164325716516653047255405504579949100748256151711511629536990371369214618891976154569727069282797365379883808745758560135869053034718688984357142527;
B2[169]<=640'd2352369140841909978192463885775481748097332209130213499114285268390270220506164472171694793695269458856129508974310163438539911611688718402975314584784944759773842938069668160445313305347620863;
B2[170]<=640'd2919332599604657950523467283386592070993381745876617899141953221726533849902705527399385270518772041569157532062879566239278821386244685914198031365214085345590289880247051679435746223046262783;
B2[171]<=640'd2121935863959291809606478946651085778781968705662643798530394510255553813135150368423407973099453275986470257639930285847003735959149080887658396469729043195926188830198859671714287852841861119;
B2[172]<=640'd2108569342849523215771215581857322476712829631960820598155652714210030913077965653843323864294974166561097842593056605923589010195783252383505316616681914169333110425156526629450718272641040383;
B2[173]<=640'd4330614778609847445252594321331801878193768292602042885418422779499919644122116777031510449368776082032246730355794457250805164534312982002017553556319594536864593862875640417860189758102175743;
B2[174]<=640'd2325357536102453583107980004664894607617359977200799663085476999558950707989293269104677869936619524802845956968975285561861426269105921887484466931208683181215954873957394240880302389330968575;
B2[175]<=640'd2751415543419707459557821055525936755434307869570369033500654186755307765991593365537015771034462594270728691859086396353384349689249790473775918566536640835992266319279781941754072302144716799;
B2[176]<=640'd4445761854182069126164490458207128826606447629909245721105354971922571501531619179767099867901419198093938513121203028171187035282094267428158841094647007857043502540580290278602164930659483647;
B2[177]<=640'd3412500790041376694044961734282889415208596353330744315922979154267723916649188641305560353685300947053588900769108490505317624932433073284418588521235605855213726001811340203068225938356436991;
B2[178]<=640'd520754116422216666599425043224272673039822252147651542377991159553516556137421468708899853785877464141813453726813237084233459733594812256232503152700453015152746524632424363318167028688224255;
B2[179]<=640'd2717860624481957746552643086696880933379647828167009902211630700994266736749120080812565869550186405633519302724424127011449396895638717161684778938681175813240027194495658702319032910491942911;
B2[180]<=640'd2307988320301490463837404631487292048475818231382886942294583752368566398030056414437768637544771725413286359927240636002408533503757497729370755162586437831183159697692216463521814894734213119;
B2[181]<=640'd2299075145439934237000750145563975078528263952617628136515434504028516182297419883266667223937100559688985795021158653625512434851400949018552672873616763585983543127368311855201461832813379583;
B2[182]<=640'd3439657011452583682920890811355441940047822143049805215554526445359204301823503476419551014975177371386198357040575677276362943742831447467729290774478849450630684170737914022792376717739556863;
B2[183]<=640'd4423206992235371382782118867706178665102683425553035223033876783482464427753035902073367978196041404564547434454484760707178391169961612137414522798397288299824914160022297957696583645888774143;
B2[184]<=640'd3992205300909150968709084644246767375708204629103639243998679147251076998899634563895774314518529346424515629880205244881879287013917653242238243861430913721914309637030814315968769102790524927;
B2[185]<=640'd29772774206721124477326526366958437514029956046945045914462893687779571449075551547069454782096866843891113057064232433308863099588887110288942250739055529215608716477356727669853519871;
B2[186]<=640'd29747877113307838519575451974533778133009570200935929940412762022656854777277536281770517504471854517462803260771097979622216165982453588108311951365687042287834639741906088921017614335;
B2[187]<=640'd137037751662294792454872269697730206615689102074107085493046701450375336117256504394090769290285643045624013523657966587411620954316207181795787659212614908919759296473439149901066797055;
B2[188]<=640'd137037751662294792454872269698373781396327127172028987570146616721668768532245775172355466764767225025444020745009705014971650348099204511793688860699225662633360293303532852907876548607;
B2[189]<=640'd1037378892220248239628101939107174428843463775481863395807633364404599589850443254201030114079480855062461893005909044567103768988831664330152304730935900010206998000667320366661631;
B2[190]<=640'd1037378892220248239628101952514982360535947274559169171908454762796298728521205515368356959665281283304583874008387854982984537610522319469269801897800730223132976545362973837754367;
B2[191]<=640'd1037378892220248239628101957542910334660736912106660935822018350865446182592413866869985770066640898273980520678871621637515069200383821551894795037745709623196186459343154598379519;
B2[192]<=640'd129672361527531029953512739088819076967675765148687192250940118858803689118203030914723794054627472233363713271587422264220903821952774890705950936131206568471028332912048104013823;
B2[193]<=640'd259344723055062059907025484868448550231568412652352449920446148797265023503101964766298671730825206915849843326807073732095292757561654062718000258204986662773049673443522631434239;
B2[194]<=640'd64836180763765514976756364686697885731185181490323887007234655183514719842759641457418577299793155776136407592340359487887149984711550191621790466875552367339446664235047991640063;
B2[195]<=640'd32386432090494200108018434884839738678707851780813329939986161812512691199256201760492669437723284297298823780576638962468727345411784705543537408800411178099135115680388103536639;
B2[196]<=640'd32417162892877233346375452349330584890111050725523479735157302605993302227618534535046634339795618837665348179302218093903338201760366887909978691450466479427646493356073785753599;
B2[197]<=640'd2527747619355312476165093262532130435090206601086157711980497579844457211984777117025611494517642810453548327522601108598443034221242658865338651519711096232407858112564209647615;
B2[198]<=640'd15844603844370759213250785629672385282375394413074043707634080921785138042940799860208327176677498109997589121453217189314929325175682796738820481735923440913614396401226088447;
B2[199]<=640'd2026146107017764412057013711797053755346549580608622236420080462246426785539777901270568510439691615088625561455209868413937825801481705279326318996040263866687184710484692566015;
B2[200]<=640'd7729075046034516688893046116007264369922411912806375581063932533225267834041371437439511710245552312505535518670060282221318197894377655250188962439671503745318000057647103;
B2[201]<=640'd3864537523017258344642977641205649074378716294387963084211465269316401174121097295923700850667703656550784354811559319321424588650543715863703190009297271867008383243517951;
B2[202]<=640'd3864537523017258344512042016889803399578188706684089446133102627547645417999986440877735985395700321451715234923825394426879305394551747120852481150900546944926928974381055;
B2[203]<=640'd1932268761508629171679904261455180730666772966700387272276421672522705206026442822382938207783935142864446304803763987236079350341044017700085503011310705190795587419635711;
B2[204]<=640'd966134380754314585401317789269507354751619063974964821756785842781773004810147981982965544055231001212528762771449583428685161836059984989406297638520214604116639283675135;
B2[205]<=640'd724600785565735939433975043075979114855257492510300613115079104699198672629652580774597965769297344671962390147864776690085272193060352891514074587385102159731799835541503;
B2[206]<=640'd966134380754314585977434536259228317695811294104294230861997800371195943796192937148911759056940814046576522854454741898328313357489782749309823728526962348504936213381119;
B2[207]<=640'd208851956983437891961392306604892796654548837272882490185947798502454866618601775473308939533497875446120407331896078033720755891815836116417374148394777804650964951906291666443313432494079;
B2[208]<=640'd452512573464115432502505465914408177636389637193491541623653628548627386220043174027520367003398058155770967471254707745557227385279532853475020732880239222777003453272438213725914346291199;
B2[209]<=640'd417703913966875783017033631252615668758031012676995879798620469613260524249362462426192736618072851671735481440058127025256344495426325044280390963284768844950703877595415841087139549806591;
B2[210]<=640'd7261652245662504474990904403186336008759245241229302706294334805843026647546240948978008968965398086928476532904341079332598796599053098154740919923987932801427654750516861382688767;
B2[211]<=640'd3263459135668912344694706829945001109856623401401313801893854319648354702928349446564833810006744186798848354689299279878216206819702657650831761038560721650594831405156860629379174105087;
B2[212]<=640'd3267552632777613436700354470659451202327980355104464935648743528583684033646023065598019048183570127446038950395240682996639796915290495953597418444955069358262479838889147764997445648383;
B2[213]<=640'd69672553068823707514818509138182533273494968518467818365004837128496940572092763739710580929531296422649392759055067167800103680804677924349345161286421659195290028318961597796038767280127;
B2[214]<=640'd407913903516443123859253341886857147763981984599055268421923384033825447998453130167669322281980903579173734323381231985686418172008132332690959177649474676167730150825352730594909356031;
B2[215]<=640'd9110078593385149638888140606409598565932634226861540222720838579126984615300522179038069734027591778428551122666553634322014061695680222952198575056614548919863256497417897500073611231231;
B2[216]<=640'd271942652282611890293624375477677979014170379192556327839065879213862043453046049260089855909536584623293588522937807235352563575744479731187600864827146017627547270078595698578635620351;
B2[217]<=640'd543885304640412222634568650964759847142751429060760493686006292284398999656450272150961119743866144387192919065320423789471596563070276224490184386754765593846354733094897902947913433087;
B2[218]<=640'd71289222420956081115713575476368981471137887366185309685854261243769851566141514968810086857157365859464195358668874005995611389088872090636994255075230111580085493978741235725736872891121647;
B2[219]<=640'd142593673630442212492253625965141325258865428579815267639017691140558832417401197196590047632254210737138226482122409544049336790650755290040761895432132773757985643806341206992077827663200247;
B2[220]<=640'd1087770609287749696510384228883213764874052979347236457370172493664076868083391634644084611041070677948489117358882349771106728790353192411547217477825685493910672848547822616637127786495;
B2[221]<=640'd2308215512021816237371274191786777871767287680107776906489064850091048724010845145327782460280156230206817385318006910974762204355332480600869232246715795101061738688756497397357193196973588475;
B2[222]<=640'd3170651176284565101911175646496299579528947749140058548181927210251302016780967008665031647436780765358606153990743607590079100024031918481063210459038461991256141486173958866177727397455986683;
B2[223]<=640'd1024766935598735254185049634862580242629894694640587202998674259677836913512877016175094067422918445970423619745384911086951576447642037832584958845902617847265340746269172342793393216193298409;
B2[224]<=640'd2120822005847817308664749046396867638262854518379753645473510826715973944180875891705122138550129262638339971441287843554078654997278092043243617461210151179244197055952455326786330351726231545;
B2[225]<=640'd1853491500909016807572492897625366193444839536133295404429456302707099701263819485057648454279269800293237256936516620681190628398613777517114971042823060782908898309647044787014326115938205693;
B2[226]<=640'd4562440617622195218641141414000892752562462948262470733817091382330972342347971658353715954922132488685586621759933911743013705726090404393722164569514050372284588585171756831647092460439273468;
B2[227]<=640'd4455508415646675018204265372229265925424795967858122979953616153475333409869807973794887862528416777042900734688115629380144771664826352993366776445143537235296165572716545501058899316726054392;
B2[228]<=640'd4526796550297021818495533678568332977376252653693870182298187901763242893464492962416750507572333674973691750059287830724802692377558147914366199058022562210843140277807310319995020956223700984;
B2[229]<=640'd4562440617622195218641169718719078914122657109397357988795979122030918935695715754255720081867110001189781529540671483655541238604607610757586883989224097098303647887162967041162691305506140120;
B2[230]<=640'd4562440617622195218641171133954988222200585459592187482671674382977341184221894559076365747441117624385270061869762722207622147994199251521373505933658733652455280566974993096979604447275843544;
B2[231]<=640'd4562440617622195218641171133954988222200585255005274489162807507152985132496947545536237869749568281679559555861400446915462467789818481152363684003240975679950842490896459763723636897537965916;
B2[232]<=640'd4562440617622195218641171133954988222200584845831448502145073755504273029047053518455982114366469596268138543844675896331143107381050512662167004181303291886572601688329302677757748430462557912;
B2[233]<=640'd4562440617622195218641171369827639773546905449018526255308931881755637787778183371240180196692624441789127390658961500067957824824931566992239419148557289126570352050078619002739872262466334276;
B2[234]<=640'd4562440617622195218641171517248046993138353064087124438666640387033934063698354846438577649310555093712653588804999285959311340468216825966902082442451304772759031999111736875735660729958715180;
B2[235]<=640'd4562440617622195218641171576216209880974936692861414766608341807610828132705236539816801090648432631089979402650729366860229583303660185822587159001366689615333916882884145039987988354685832998;
B2[236]<=640'd4562440617622195218641171487763965549220061249699979274695789676745487029194913999749465928641616325023990681882134245508852219050495146039059544162993612351471589557225531377031512537354675714;
B2[237]<=640'd4562440617622195218641111104365168404558425384826683462393535006005960366148059980448661998655018050642357303854531402968571555556513937074072255716946037099897562525507700660275178604362583299;
B2[238]<=640'd4562440617622195218641050720966371259896789519953387650091280335266433703101205961147858068668419776260723925826928560428290892062513444852553859387591958303215441542559677934249776924435893516;
B2[239]<=640'd4562440617622195218641164293648093233156858539236559265808216366364410610355347407606206085420556764990241392703064375596826593126424526902011311858623165102443727688221680438095922318058833220;
B2[240]<=640'd4562440617622195218641141414000892752562410574811912024428065182529511835685250376855510846324072262587825620559792986040548372974400902896201606999453846183388392784526227701505215291975916846;
B2[241]<=640'd4562440617622195218640265854718334154968690534149122746045372456806375221505867096993853861518397284054141639159551769206478752311393765684184860223819703631497638531779776518964865670392502304;
B2[242]<=640'd4562440617622195218579339005332015191378102876993648133070409680623972207230161622482688505040738432986063209308283646063289286864877830915591856022247694234129472785990212637681050018497085445;
B2[243]<=640'd4562440617622195170844571521022840117701116320201740456290059304090087103815991796553524059480088069114997804488375963070938701643762938224618975170210936840524645376089771337608065107585918726;
B2[244]<=640'd4562440617622195171122818222680082718519181656348843545079582071828950423719312734658033437724936419681603755682274388684236081998026273971097054632145632195592691837532145667101841575215834659;
B2[245]<=640'd4562440617622195203793618442267984764573686542287864553782713717167151902367579550429176266640880248710585858365847862778903491928344079167598906029008271710940318737482460943715202513793855666;
B2[246]<=640'd4562440617622195203090272613078843745839132498138242857120308943160580732611962734664999782744180251444998592847937953589735113810610683313637320174365995689356570193476039376975026554491007291;
B2[247]<=640'd4562440617622195216662528393915455052409208339091382410298141725089580447896172937762735010465116462416111101083650047393907333313246329486983690470386303135125006883824761689501003097440213389;
B2[248]<=640'd4546845471346074262571060770651675463983613362139178167607056582656476629330160721103175433996725900676462328637254716223410566336830658375713363637822204265634303583365262634261092751048054833;
B2[249]<=640'd887758012247691621255395402870607363746778858792451261327563967769159758705783455899487542928239046481384179877028119266471202411936443265505129561374140161825460734904796975951259040605721106;
B2[250]<=640'd13401366836984904769905507700658564997241068331585299058545526437483452771356451504994836001480505908636339166124861537656005503065961810525816999070507465168923279039235635301111360043750482;
B2[251]<=640'd16996415706819964380952061890190350693517299118271396172471981404412771555765582140381042076886338469726239026222884147430958874208032931954550588570411184874764170854045406633746605185;
B2[252]<=640'd531137771208727378787925688342209793725710846249343128513635575199905300624938547286609517661733934795121018806732903304885737555907426644415171470393053309757613601647680297226645608;
B2[253]<=640'd136054316456640851429426138854833630474138666900516614734580054771397088790661009897335555221977389539201877426877079304447339295766538074281912878806744522477504841687776590226861502700;
B2[254]<=640'd259281406472284945146306002835316542257628895889782396018710582963306019023679486991986089560522308923495030909321239192228847321131164674419284161062209078811388926570514191849828;
B2[255]<=640'd4517951093198658128463245936927492457616;
B2[256]<=640'd2039283887267322535674134719698536285312;
B2[257]<=640'd23717608908436910108460621696125895451682;
B2[258]<=640'd6427752177035961110578263940048114321729239897176631530455104;
B2[259]<=640'd24003637036118667240909207045150939705097248890084020489519120;
B2[260]<=640'd15216616496880454732237948070544700168177026360719087807214710771630812613978219751615957187813433263505503556450813795950340516928563038777624248985815863119413440085148448;
B2[261]<=640'd7619630135714691990175698699015314890761263944020793224895254458276827166295899692371278321927919277222830785017914147922700215372518417745166060516385237366735815193281112;
B2[262]<=640'd132784498204191774672397051638117156832398279431757980799861034550100889965213060684790625566307321417222332371561625253838327097678260440297098431390369464786260274479610447109628932;
B2[263]<=640'd398353494612575324017192029747003283391770391301257025334631229423963808865165647453893281405787909919619273382411262365918553610923070898808094773733774502662295059421472936621654716;
B2[264]<=640'd7029532692261849434245817057221849345714710528298013850630283949023848223840299345004031336377342054841508420956022054907701847406459606715400780329777122928533;
B2[265]<=640'd7029551127997753105316828971506221878753135812426017165172994281944715050877647878048071245249183569797957915053180716083510708902449743377128088150622932315153;
B2[266]<=640'd7198262071262567431281069328920963956945663637356551406312206307636482129168086217973567882337998899242327426426877196304040916462741214287899583132823205010439552;
B2[267]<=640'd526988477247886105745472322831314057908270446649721589420500409910666276011613824093740400035991038751211965084649071868838785746261994358909422097426618314380850103834886153239401913;
B2[268]<=640'd1061757296187424073288155410407052214871008258263585786360912768068594151206075953581443319297548682787120748041384750899013545364763583399942612815432353021764508479807281444901036673;
B2[269]<=640'd1062017527342638015386608233015715200303408557824883017727103405627166728304720261125750362633021992909847746672020795858108135150956089877678433262754097620497105061611217149157722152;
B2[270]<=640'd1049600496465072356900438448928462865164938715854335547515276510206787653225409720065218879096663145117004355182750390990149468086005736496868508508357776102983375610137257186586835286;
B2[271]<=640'd1847800482797549253916055083633270955820422253191450353840710660128885136589531119340039701690884943513115569342951946198377020957582728005528539469242100355337849385101860917478628;
B2[272]<=640'd129669146247407729293856124616541745757875990338273165139886771881896991220381838313273119636462457343134102499383395292687682200329411344318780994809933331955786746170090786918464;
B2[273]<=640'd3241808980220212903578943473078441283687792156247202800566205662709710438299345561878167899135307082106671886004436255719559531101490349900513677246262337920173031214561663869595188;
B2[274]<=640'd8299031114574760778921265659210210956042751313379647080163668626125880819108741023900428881180292032141491319073644256466603296210776332453133245309715428324238249275441064918189592;
B2[275]<=640'd32288418020355226458424673689346847706120523866074692816610259653140140621454103811513429922813847328723437433924233966836546624127925667210522387227566707448815028796839278453278246;
B2[276]<=640'd129672361527531029953512745740348785920403303498694781791061077511632293469939309083757763304932784426705789963328072528978319136450295563033495959053191990358581478090540431709952;
B2[277]<=640'd259344723055062059907025491480697571914121445216156371796307677112641211742317561064504158560360893355686013618986949278578320107942408163036754732752065555462501944837774745340058;
B2[278]<=640'd55209304643961611313007586626410899114220591725423499491214068245199201053857713150828908385673259757419711422944524143346851351276717982934911453593981647597661523120845666570255641061;
B2[279]<=640'd543885304644369509058138323509727874385503351022235142192820604140537662303349678217546690702432634215480915383685666566045131761643491901488326240696617179246341257825318646192841717804;
B2[280]<=640'd543885304644369509058138323509727874385503331209425577265787847483385901941180636788882337914989800212087725162700480154237125281530924832507652164512861087051680977787530138590130750610;
B2[281]<=640'd284596687820040655526815807989641265918204797276714164577837085291585359804654240570215103634479544475979750335240957479821493669149904790234216231305357170607108570043843293102098367868137584;
B2[282]<=640'd4562372088073810028083030280271529099181055933826138316523767925461385086494754741351512347258421625190622764050736199770791878323039363626150773442964990965895828027420525906999479934491178776;
B2[283]<=640'd4562424165091729726463522597016005155625028345772145217852268778497974907527380241927512562225169069717359029886380941255204302881335636117863473380930631670617752181448162094808137830703905310;
B2[284]<=640'd4562440481650869057548794341165710447461259910872721792272949465421900423924739167308409509297238690927679968356314738295919049939661992996245543167539568767572616875850043955838792662748654661;
B2[285]<=640'd4562440617622195218641171605700291324893228507248559930393121804479599803228050491686583650522839337575963515682735303019915616930420166414115016865600367544004233827627404758062465451533959688;
B2[286]<=640'd4562440617622195218641171605700291324893228507248559882945089882462381988168192312757647647917131445407026294593529783959178913121743663072652750586084180471945193618416778302863587445715286150;
B2[287]<=640'd4562440617622195218641171605700291324893228507248559882945089882462381988168192312757647647917131269537486252486393400740083337079855410971056510198632509871724891655915682580168216659358706464;
B2[288]<=640'd4562440617622195218641171605700291324893228507248559909088025117926770627446271034873394739548903646976021903170492197937546233784425641089435673815441746335054967186364534910892148864186343434;
B2[289]<=640'd4562440617622195218641171605700291324893228507248559909460166544766121355407524824512053061137968023647928750034615179918033549298485377832445491780758881978018385629263773469622789184762725194;
B2[290]<=640'd4562440617622195218641171605700291324893228507247974578908956951637444528207848630949452367465501610685818018339793803358471805767779729051299906789419824971836687440854525114922851267480092804;
B2[291]<=640'd4562440617622195218641171605700291324893228507247096540239360797064176730868991808455012054015765626889376175565403438015526991915594063340576236023682912264639893064041179417323276643638441730;
B2[292]<=640'd4562440617622195218641171605700291324893228507247035639294858537317545871686317442020684003630523269333886861839402331266343116039676069783866190631872423402404261213637654991153387674746307866;
B2[293]<=640'd4562440617622195218641171605700291324893228507246999056304034521783584368593780803353038512246038914203212731093781721441278821911315284946720915334436470321655419375419093740034615190972547434;
B2[294]<=640'd4562440617622195218641171605700291324893228507246999056304034521783584368593780803353038512246038914203212731093781721441278821911315284946720915335058837777512521905024666099780258792721129745;
B2[295]<=640'd4562440617622195218641171605700291324893228507248169712010403018870352467554953240717694236549538278384784914953641235843336234018860399735369724823620112032313317142060881537325881561002803488;
B2[296]<=640'd4562440617622195218641171605700291324893228507246999056304034521783584368593780803353038512246038914203212731093781721441278821911315284946720915334290988156915447699342113537769360715954577060;
B2[297]<=640'd4562440617622195218641171605700291324893228507245438182028876525667893569978884220200164213174706428627783152613969035571868939101255131895189169350075975828425873157762236316568715394948314180;
B2[298]<=640'd4562440617622195218641171605700291324893228507246999056304034521783584368593780803353038512246038914203212731093781721441278821911315284946720915334157065012579564698526428616984044684916091426;
B2[299]<=640'd4562440617622195218641171605700291324893228507244657744891297527610048170671435928623727063639040185840068363374062692637163997696225231128271887183255091258459883664208696916253647835479245832;
B2[300]<=640'd4562440617622195218641171605700291324893228507243877307753718529552202771363987637047289914103373943052353574134156349702459056291201599622843085329630831089585258408592455490484785790265347132;
B2[301]<=640'd4562440617622195218641171605700291324893228507246999056304034521783584368608911289168019020763004882825418172184425910890686197373596927923302839910550159309144096107237209053570151569244087296;
B2[302]<=640'd4562440617622195218641171605700291324893228507245438182028876525667893569978884835856511031838444120487784717357934739942795040124270486896933794756339173500710488273746403133977134628799631122;
B2[303]<=640'd4562440617622195218641171605700291324893228507245438182028876525667893570117598482793789187077247914664087473660280122872165087015312328043750517282247708585024603272801980080555804223585230955;
B2[304]<=640'd4562440617290233973130692169019298695797935615166003357724639569783931784194304003654889053961247470071392665456013513167048458378377483779501584158196483456987727118539220575068418612329469968;
B2[305]<=640'd4562440617124253350375452450678802381250289169125505508434942093784105497421973384926587582120977559346741163505351745661589114981877127274481437408956745012022965649379996091884171306937910352;
B2[306]<=640'd4562440617122178592591011954199546177318443588551169941025189372420875826463244042333167607605414865797408494848046123969263618077177732486255589147557913306542761343571768914090117776609140804;
B2[307]<=640'd4562440616589484531435914483150515817817090775789947155961066535383933352908139595695048039485463305731762712021604509944737693123277223963094825993694140851760093392350864755510864751503631499;
B2[308]<=640'd4553668834366618134027852163407107434039761668062605924951315867015580934032162394815117259566649386488220660195631149755070595364291125955435552057766191354591343392376290310663838371772647637;
B2[309]<=640'd4553668833304358357439508907406675210028041957001470722580951968121388039135568559560949035327719928902551926041697055290019292800235560041086728511294903206857533568801090766251663859474761889;
B2[310]<=640'd1903598812683433450234132852533848731787060453108042169643731597175458877991931679989661998933373998278287485388734366355458244055155681144902498832298278714047269085999216903659287752705;
B2[311]<=640'd1903599590717602615420312573610316469975808174894610612095919842921395351647713378161630831088611197561906006494950874234918353913823327176860461349478611875762201464731763142127703293952;
B2[312]<=640'd389017087481010974164203941480685100613522215692644655190543483039750432526326478175533898644943371741719817315222693115429091797466787151037302659056824827846749253328045191514708;
B2[313]<=640'd55649340316706700862229826580389869882266140403410852018690299497728219254817955134363426309763951802058199545946279955189786175996987795212885910941429640615243925276072132696;
B2[314]<=640'd2090966829631452553040653094182306584683394419768485648432238284924437543209278241855895439755642080504021208470927827772674348766546540537372478366776917509499595146825499341521032;
B2[315]<=640'd63331984303028417586482097754799006183741763518715189698877630482140897137024939279938979161916278486204053444798582403332529454894127306585613004300273490276037127638261338694;
B2[316]<=640'd1013065324433836171509127325413703691375625100805323790146832664162307651449652674503743892465566210110909599795163940189389723347460369464598370104538234917714547429090395759214690;
B2[317]<=640'd4562440549636532138094982973433000886177244209060642385809663843626711610371689581491273216993364506973721926264798107204411184748617897319883034798586630027679771078621201403738376252260261952;
B2[318]<=640'd141671244153765369719463870507813917148985767027911528599563805848489187496284130137403450600009036827568341666171625214097029514303402852329299528794434450752176588530723181864039843468314243;
B2[319]<=640'd52679396866785518494232358655023498740733269067989600152464930700220719008209400501704111129823700457439796196251712504120796355433429120944165974969016546471791922348036932650498;
B2[320]<=640'd4491152482971848418349903299361224272941771811822801181663892634807114858072488385596982821284084298502879503518022230084337556722416107147568224497318032777091301175467463910391717505146591618;
B2[321]<=640'd20572825126372745841735421417085058149833646439770082309364516825788063661902527801796976215375559269528884501197891351347592;
B2[322]<=640'd5285946195752592098919093292564290400873737727615918228513541517424037715660072531175617776731422585256539857841554914046464;
B2[323]<=640'd1301494286210147037133296636426580531722647459094999205199557936470450078629178422235546173647536708674897123223290687531104;
B2[324]<=640'd578464320345812632029639268265737206910375350051932016297004735234540549012542749347822052519076072550517582314261215707172;
B2[325]<=640'd5043456793138493339171717132818382567049280289905719559700125911468352362710376798742557882238666632166805764410726482;
B2[326]<=640'd2521728396569246669585858566409191279730828076815375300219825988645205964130571799953497227095939496344337380295188709;
B2[327]<=640'd4545593226425531228728586712991253994256263155399894288745693912715381969723602497415403017837912560892497812781118798566859318968932410327986466166252668944499206442324795204617196317547301095;
B2[328]<=640'd427728807902080801747609838034402311708740172554552493491799298553057046928295831375302178251370861278089210626912741503528058775802981287351944799729975736547336281481541873772348908888152070;
B2[329]<=640'd30067159095417915789170058021143723802484765054879984961162525391227759015488769301238315830470764920375326775722864210204733089948779346283421898691600766171929256175603798;
B2[330]<=640'd499051743775992878936135706500705365983156802319023441268102190382228591081173970800949512322418421553212892851538705003660476685205098908305804565490838742971896054414720317491302199282377737;
B2[331]<=640'd2281220308813172367105026299329401866378459834199786188405717477402216174761254236602694150416102057287648033432133385326092643686209674956399338366358019512581118011245514144139469362190615554;
B2[332]<=640'd63308855589107074818760629393685136241292268568645947782281188032196357332153308998492286686332635780168875829393190004581756218055281836168219069445942600702432742649046779141;
B2[333]<=640'd8911016831293350036408538292383381493932086928219843614412485386522021810954448022794798273719984373051669951090946804294381733388957207705678593770528871788173384534541403868658055069696075;
B2[334]<=640'd9100889195575602517010688665170593740723707560193648404254780806407092258132918171154032465048188204414815266;
B2[335]<=640'd142206566528832901151493151361057498340577673345662461432984833869233366399069741070897661013326367424709;
B2[336]<=640'd42678729767328520174318449706505070388089970646301995802403834394064269574273626619739546354680263766134;
B2[337]<=640'd273406340597441332714702631970096383914704457616587160711524330917192072481562783547455015941596752;
B2[338]<=640'd509892473104096414742004678290369882236409393017950646271466372672387417466418153029602700629964762216152135978825680952226974375949389754235030691768205330314112674841876556903247775912;
B2[339]<=640'd50989247310409641474200467829036988223640939301795064627146637267238741746641815302959632774576910499960022136021016751555828168758081709032996205506284983937212172604354273122185777746;
B2[340]<=640'd52494151415463241183448641223644459085696589679357695826836451056861175922785606577434394944317555481;
B2[341]<=640'd2281220308811097609320585802850145662446614253624279965289596258949637583604338693252956405789920752502350250186707944503961887611145794129039596088627496814159989648295110331555922643458850860;
B2[342]<=640'd855457615804161603495219676068804623417480345109104986983598597106114093851627009969858652253242211191290807856338733500072127745550394789868114032131978708204723950005947792636951590629020672;
B2[343]<=640'd499016993541674912448519618573937192697185091621250544202163808791870488652190835790899516723684753256106746288851907882375218384530258380202537528047117210392942468671742279722249918079894382;
B2[344]<=640'd106932227470143855641723196608834492445679154959107774270482138211582895350824249567139983095664827325776176953621411514226026849992843864698163098486966676225726006214927564617228078130661946;
B2[345]<=640'd53466100987760100218451229754300288963592521569319061686474912319132130865726803558681194354408952052051024006186697741136647979622709479372771555072689946890048925863676957694752636372794217;
B2[346]<=640'd53466100987760100218451229754300288963592521569319061686474912319132130865726839632295265882986958976658699213339830381360694378838681733812817796268480844326707066396805490382957351139019078;
B2[347]<=640'd53466100987760100218451229754300288963592521569319061686474912319132130865728841868311390245331782550674485428707051672799731240734671739881049143807824932531967721798974726900900054520039746;
B2[348]<=640'd53466100987760100218451229754300288963592521569319061686474912319132439747195714254980706014319542979989495321909458086118238916755964305266026882687870603445682363985157458714081619620139297;
B2[349]<=640'd17822033662586700072817076584766762987864173856439687228824970773718320709446909202834214286716331060235919172019172961368792521943701400263753860232637545526501313019118404762827841755814153;
B2[350]<=640'd178220336625867000728170765847667629878641738564396872288249707731794278843168245179533678977873861078992164235388364019970820547678702177151404099703517521275625596326518982075733684176290049;
B2[351]<=640'd213864403951040400873804919017201155854370086277276246745899649277882366086985747847190206267683346518566616718218056793406328449484924975136254866264050520413243953314487668612453956172515619;
B2[352]<=640'd1256981993432118478085064844258223594491869287656483036041915591253838672066171929806174534964502296322702325221081184112149483327682393794862282376106240;
B2[353]<=640'd157122749179015135391480318817827165701874356792181004940119478255338898576248547562985910732008924285888828702855297686327381483604517320961076585038080;
B2[354]<=640'd71288134650346801033259510758380654132964260882203206396029403732189500626088063235552967715976039247728731988166873234699435176398771827500386920759293686645206178771226788252290921204287753;
B2[355]<=640'd71288134650346801276966910117618550455131668658688760857059106648214834910936777748840144604453906919819885674602069461434861420230866790594522880155376254816972195281753023887627434880926093;
B2[356]<=640'd3864772934980064587321221919685254353074331924793947055165797431356850860809960724543641962998974493640887638288148151922000375161803289619590226561281781829957116535767076;
B2[357]<=640'd71288134650346800291268365307231642261002542317154123054640580097781425452889730324244242217607939247147451787603210832867273782400358421952462509502519575551813814582183933325920553467642112;
B2[358]<=640'd71288134650346800291268306339069688034124856474701876551475022874710208658422563445001169385600935836394706530830250767474835800752321992235849288303028977844147363918735330964876752687729024;
B2[359]<=640'd71288134650346800291268400341283913499734946793825405895360476984595681307783602154330213762184149906367324799459486643655634441248660393825362668665640308273135575161407832594520067377469440;
B2[360]<=640'd548236387081524465130603430097805697386929579138812861162682470357575997173236268530934905852797304223399116702803979272721460116983917474781286192829925688383102426375911685101838874580992;
B2[361]<=640'd217779358359533653146194030937114615810181237596874168973109304008234031236250221671861766948013448742747317715997394320922462993615943544331223034262345573214061232862553550991321628577786880;
B2[362]<=640'd150377760110512436820466548790557640747623977821172708707067936830923592420358530537602708320923310324916366498098265133763630904442552112264534887422204135942102776837408969658919745491173376;
B2[363]<=640'd155942896526128246456432368517644834221139920514455013031802525850049208179999947896516309948404577998293517359209659979375463717124317674520678813514894445703871593773824524286799355316535808;
B2[364]<=640'd169310161117154272450846551863003427495224839119529927092118477660199287709975558661055959836508142438908530592786120648013309008661811785882905176566310639868369789319193546207234677060927488;
B2[365]<=640'd35644071574277342679770942686239178827879172277577997662652826075898859004952588954498244464497306606844073998620887639818117289616759173106989460303635893162513681235713455580372137121153024;
B2[366]<=640'd249508479757823623812188679386096355220697742642996380294836977042156359277965051271606509268446091174989177771146060123733907294576385764857909099236412740762177866237400698054399423913394688;
B2[367]<=640'd285152540161345710341271515697026539280099555773363507841089243557821727367455968720094970883605353549534022392048579896836309878917922467039134917492032738957629496253765474303959057226401792;
B2[368]<=640'd17349756746253878273311400656970543200560523202051729604130314328789749293963100636470655720915200652998109989799810107011665383307867403625414570084274705559370962064336459388688448;
B2[369]<=640'd86617085239092992664261331265866086614942083255366027072409124409606548509841216139431606036226384386998466250366768998689137158007729405009517469206646311799225182865854134630400;
B2[370]<=640'd497942612299331655249712162043223287950789080020242157831867364059930386449498910704280771932321577099251543231814913807901079623215261167427434184453181775549736292238229428435427328;
B2[371]<=640'd489643145672633006802370368870308101906332432797633895833785733040328151084303643620111686731919700698777164339709209207578010160949187491791915726606632487766393644178456840585478144;
B2[372]<=640'd62242738355251972121267365000028764233272732074375723872320555296280807584036561296138698856157433496518092488618230488371047144993713422538147294775087818142407109846900748662865920;
B2[373]<=640'd14393632138024716006139453571714329867029469812758168536412101022389951407891277005467401624730757237480602262875483180454274713244079373711866307351577504626951422001666788136321024;
B2[374]<=640'd3638930645635322803083345462751835450693193628433982036097197441966494297159878093468814639947187321861370381081854744977475177935275304222145543131782261669865179507040444108242944;
B2[375]<=640'd908687937734143338616175068634087010968639276946139815105203605241129730147188767382291645437911401798698808686220663743305634129772549033303580738178767505449353578905553040572429;
B2[376]<=640'd230028650569170429148676625845328323462695947795808801249582735614945493931043548161877039908034571891325945415952420624029672069392802221433856287478138719241694918138233580683264;
B2[377]<=640'd16335677390361430862244456929959359708383582370989812475649056327332112257927830687856464967487968011182423823215313342140765342401055303320376720025582964179239009693441005191168;
B2[378]<=640'd15582283264354000943780097915097766836440347917297602059458633033423653603820580569394419556878635448039544952044785355545781024919968758985126773873037012648017907879803617280;
B2[379]<=640'd6078401011601794131112926811668573804761512491624499416554746922659848248047806728213092673865857714581202889017054472063338933458131486763573661364289072218434018851274836934656;
B2[380]<=640'd3798996894664566320988093385614903598038456721571705055497102000488981117684604294102541597685030401887281313598330903755956147532819729814833336632487400197385346145940123156480;
B2[381]<=640'd190939190689393030478411944979666914880073543788762044086028104524885831287719913518746340475087431204342360595475924762408137837342396645054026755700692584676768341567867977728;
B2[382]<=640'd31905141538569773157863743037757642159663884472025379846347114487180265805893095956959358327492505501499646083193376708774129066534185792652302527562570474858971848360188706816;
B2[383]<=640'd23805524727734844318247338847008284469502802341716076005443164393613889247342239031587961863462825100915218004782532840173670920449426366087581709677291160131786030217231859712;
B2[384]<=640'd5936170704597009437166999161738988102607510205101144331379332938334408142264653189329030171443231431203779548345856006325295274374951507395808515744450340220900395683218980864;
B2[385]<=640'd2967979913296623316123190611096206457644760224727920022840312632246040429797792891032631593340284196659041483125964328355090924483797578428931540904485278920338826587323498496;
B2[386]<=640'd1483982410508623153649131963281202426699306362853223651255109223978324898070437625142148912921228462401469015769175394790565833905817133124744859224420818342307115867599536128;
B2[387]<=640'd927489005524999390211643440065583556780724646394854102254475845350069739220592663913058048009868397544563966980311274683158895361728965723705467166704632081512416555747508224;
B2[388]<=640'd108207050644483769152586844213446337607181762789483936944838365536471685473652689173603760466175354874021074585152139391186199338516891876463086019640370620908821451930337280;
B2[389]<=640'd29950179670596630258681299697093599827122480718239076624447283875103043034352330002269887925567182154542032136977185735083998259589464432946174758400070879490463804860399616;
B2[390]<=640'd15216616500367003181360599183408182399964490410722892825164251296701600538537147822178764177313942871033535610321751534449276961682987749061050422469526577198794259516358656;
B2[391]<=640'd3079553338654460121001092397553683159865085672847962777420384809936558670106350849016780165079429119022176709666815629314095006748166661511679905028234344903369568366362624;
B2[392]<=640'd724600785565736168401899240765619637390107982074335225016291569659376165132636623613815647610953317722382506020872695594879322592971458441828942234704725009292792564809728;
B2[393]<=640'd422683799172753448863225175945992600966876324053643867159613852954383733275855187876110960271677102227083600410623331088903329741929252889254588297409281625514030879735808;
B2[394]<=640'd116993151866198319063672796076661129446309594675773494769349850597453555581520784163725599925290706366010722496618467450535123351536565396778814857890433590124803111518208;
B2[395]<=640'd29719954095689177177349514035943898307481800559981478365357684342984129395527296901063512601207443731303538382266616016680042723890723987283741905296120725266404086906880;
B2[396]<=640'd7488956686755259473017004605977285499457574657290876488802929906806577346324222675672898724715908098230893019834873231089179073901794826784470473044022246664322357919744;
B2[397]<=640'd3316959162445527717916967279447406584290327198774594322155821975032426779971261870961416787653430178322157585478748687021324820356160579413267000108353488293934428848128;
B2[398]<=640'd707617954667755191159517114385035594859603218718701494833266965854408367138336330437311141286905140309518193480892552475194595901426029347385243240032760480631355342848;
B2[399]<=640'd88454044230174946318847910886275035520580898247468281468688101763076653465109011649776830761242632834716477294712591382735758845961676112144194008158269877487935684608;
B2[400]<=640'd25798571263428714016271204579620108004053021311593412653372206389013764587102889439598965061618095541999158661504965792764187616402490070234594479704610360186101563392;
B2[401]<=640'd5528265270734681351843031043868788994424028340065294770906944671966307455670021796862390006212631354967501643186585082751821460390504496243254595848320132152532402176;
B2[402]<=640'd5528265270734679721565956781729121151407692608451108449201754853726063015859156922068448114919496574140381694062889676072909023249298461967799475773844544916035731456;
B2[403]<=640'd1392863710790573600121215740098627717168641634651433385721116143243752811523971722609066516903702309269371811721798624913444637760172187102359007317785333647674441728;
B2[404]<=640'd691060398560067277021322431445488633843978253184047883311903473755348992300168284772944191489009304283242947346419997300228347202271375348469392644042598468894588928;
B2[405]<=640'd57588733403294614403668318614700909774024133740285795576413667224199063885131096665779575296887220760888829592976660584749860091776960224535898427766701459930873856;
B2[406]<=640'd50387834498883805880721508039920299593512366891630759631218400720771916574523220112444431712575358736570350250020181848914594215988667934391748508468172967060176896;
B2[407]<=640'd13496741383629589148452955784201979827246237910649312194392840678175547251447538186119897872842762951476110603228780063991450757914122434190342566183972687270903808;
B2[408]<=640'd3261712501043817377537688191001168625034625546175426270218895915666988001342541571453330414229911723343185812852934251939724163416998428900490347542789156165910528;
B2[409]<=640'd681866625139467246038198124986520080190266666261045371110782526094868232039882482880746274383157148661910342674524240839088024758539503673582558634623681188331520;
B2[410]<=640'd168709270542574126435351857094767995702109947449867015987863644757379790899518745303314498812857679646732503850176730458553810437712495038462325226493993247834112;
B2[411]<=640'd84354633647684932358177257721451103967380361443077838619399645930787178698320794705876270869724464249515790549129790300997810138383199160013398503910365468819456;
B2[412]<=640'd21088658411921233044424539529594479493507272707736732734137558991062250036456907673461520747173035278900885117739159191599817188200186207647851777815850692640768;
B2[413]<=640'd6150858703477026304623783121034277844750133409251704235073335265441765292215144849721403425133143197860777401813759330602349448510514423518109257457480595668992;
B2[414]<=640'd1318041150763908818297021782874627684197069031928694383870287564558009235618963054540271573838464677196057551180047850793315904651687522302535363276386611494912;
B2[415]<=640'd659087249250122599409136125189869356186978005154514989040438857808803885309915300783460840254399097737127960335879519860674071305051633561112212039822437515264;
B2[416]<=640'd54930113317570490485826200700825313508232489829271478198601644505304333764988472235939919551747912271053519898927803289611143210381221041428426180309268037632;
B2[417]<=640'd41188785960783658289891404811297669324224830076676347238698668218238636706224474624556981994016560987230117061033717055138653551972268056412859254862654734336;
B2[418]<=640'd10297196490195914572472851198622089825904412760800676997329608991737217293718432996763702487654327937932264987502537513525132754045525457622300852582445219840;
B2[419]<=640'd3217873903286024370375429092624804158124851107428013967365927167525584047803180154740275390533467388531971512667159972306300006354064213738693231630157348864;
B2[420]<=640'd643784025086692293295462525456553546080155375409511319426654496301322126513922079865211171519075812111228539932898728618595067256128831777723833269482422272;
B2[421]<=640'd321836491177740772517826798062330504870616192488140712776535015695419709894196838316732344699431311553242346110419735873285287935190822600335117908162117632;
B2[422]<=640'd160893695159311165194888300000131635515071633524498826809337792689001281817916707040503664036681783064217780569143645459106134923835692986181399152332636160;
B2[423]<=640'd20111711894913895649906166545945844855460835969476659080261121150377910811660629935283836527297849449301487341874706874429772259175130648323220042183344128;
B2[424]<=640'd5865915969371226309044311666213110442167719834000517734846414645824373266778891072475621530214601578892534440668364941617040440455952878325479047449018368;
B2[425]<=640'd1466478992337471557765908985363376716265188368854450532184915047437729630976678572150776475752221501584423371540519430372538763427151126663413188928733184;
B2[426]<=640'd314245498358029619521266210980064682617950365971958912692049857664255601347706347726375402178200704086338956906762705106636033540409047777810601870360576;
B2[427]<=640'd157122749179014809760633105448055246943139862786908207618632060152775525362337599739549927490373546415121405637511649876207752352459495765448661537914880;
B2[428]<=640'd39280687294753702440158276361931191013277345925087290708524839885925954502749437977875995394238032548565940325470720167581912543628397379257651204980736;
B2[429]<=640'd11456868493401487308292765168345386249482605904701456481910566293917238267334767521227559815270059788787828772456971935526482538774701661296015267856384;
B2[430]<=640'd2864217470888784655220763926365725374196271359341045178742223500213245407951072537006912347223316817367035761524907446312898310467290430439588685152256;
B2[431]<=640'd613760738980526600633020776768009866024452591190539794745919930230898775241829191661056355755389656453400884600692920812957504387251811635311901933568;
B2[432]<=640'd153440184745131650156868267058480843852171204657725459834985839229986753273478639256900314480621323758132851606051293634277797230686127861475594731520;
B2[433]<=640'd89506774434660129258173155788113076673358980497747224435186182827222792839162421782726377963168840624422101650974320759177860808887926251372918341632;
B2[434]<=640'd9590011546570728134804269316032385251300621227623215565439859312743531635961675916402166898003731308897971764419100140993673430700396541338982547456;
B2[435]<=640'd2797098894808673892548958149449854693502169898387138086508386282247342998716236970485683649645430316984255571093315523500728154416547311747065708544;
B2[436]<=640'd774202786226072077309280222404466832032144743535413227675737716377405621678469820677440926758982991317515229843168067181489888500192050293795454976;
B2[437]<=640'd174817918817695587117065515849617323658778608320290170506512228094179851744224147920161499532483990990710153795549999276497733204110992978955206656;
B2[438]<=640'd43704479704425305300886362832682713271714286969998348694936639101208541288062832138551266311956637983184690146884522390053861975331668771108552704;
B2[439]<=640'd9365245651674726693010186713853316218226155467827888003656246688921234900728242464511618042080283067705071128697003232429488319888759507719815168;
B2[440]<=640'd2341311645143676267056501175491162303844813736712047327304786415763202613621319818660248645615395038145388117503621481725738481490824647459995648;
B2[441]<=640'd682930120762194045960620747910443185340152934988828987360081951186637070562664377304170386795767008889089042117139510885230398230863585575174144;
B2[442]<=640'd185939719637427912524384533485376354239595170083312814949863388326132766132697707216342366282305521268416240056329674923400940359292701575741440;
B2[443]<=640'd48682052893416504828979375745370728171257377906660068807275180636305668577016026393944569102473793441007772923359503050335246055095478765223936;
B2[444]<=640'd1173124542078921578188934887947017470217442991959575794791776691346443718226484389420306973878142738420989952;
B2[445]<=640'd165131900351285148835979104461750259737352679220116240909106396435934670328561196396857131735993765511299072;
B2[446]<=640'd103445839543965292892865880659257536282624;
B2[447]<=640'd11062560692787161874640354538628768375414718464;
B2[448]<=640'd45750505531889566987601967340230418006710157312;
B2[449]<=640'd46624053413417497702067092191516630795516062580255940630506555180332598756865027866624;
B2[450]<=640'd338460656020607282663380637712778772392166509704418693022591216728198461472648125794609806981971642186780456161984468169523200;
B2[451]<=640'd338460656020607282663380637712778772392154853691065338648165699954347113292828528717441200077287975339800415349041239257251840;
B2[452]<=640'd237142424914447859860667563959872930377066954513170675232035771613799854957920256;
B2[453]<=640'd1867495154454072037241144126213238720497893351564359216947211874228013603015884800;
B2[454]<=640'd377083078400430820902664329043459383667355442251116975367460462364558082642552371765415513603754534984634091062661190234220835897344;
B2[455]<=640'd354901720847464302026037015570314714039863945648105114021429337765419895889729043284976596007453037606821165083472028841675598069760;
B2[456]<=640'd66544072658899556629881940419434008882474497766191406761049734052517842533987235658639398733298823472525500965261707189128242659328;
B2[457]<=640'd1077405652560409863528432196849057691399697193413836201702540839224929540660772358336728342807722981690402486091776;
B2[458]<=640'd2309331058939438568493808861038672275223475107039603791155926187470475963518788883497541479067244974423627633000448;
B2[459]<=640'd2292378743618982609505542648445295609345320956757751606019527741643410850643685806239909917467168450019328;
B2[460]<=640'd251978400088770166235404647302246471769131706598612972440098103832947462544293888;
B2[461]<=640'd101897040292261192899818270414085215408297289923123166692120726224361680768335872;
B2[462]<=640'd25937539305713487921939549399952946841120696043675477271297313119420064978698240;
B2[463]<=640'd1861227880749755298973234548121540320848548053739585951686610082297245559416555668361772906061126181060608;
B2[464]<=640'd383324879907010965671607409054253405878640290416133917473700731476659632513964094323473662730633562549261553660541796352;
B2[465]<=640'd40347654345107946713373737062547060536460826332520569396270782549134075312320861472599501738964004976469935384361435136;
B2[466]<=640'd3067035503326344183660662795767749040683520877065729022450511895005522810196012082856858968856233306263104162248781321079546457439887959464737033629794252422216631189504;
B2[467]<=640'd7728853800265553267504215967021742043292910602304832796473748749409516295275692712868040729376499756578940574448546883293733470685455285406452598969971004743287644234973184;
B2[468]<=640'd142462309226433608755982871029760292515840130106351490030008406732201877300244105879018324724949884662719260705293389333060409795135335962480581536514201611204968064527535964160;
B2[469]<=640'd4052261291009492730807734773817213402906595120297855708944851142350001800544632678710730482288595252019829939132894718262957224605909548107211016192859110224916022249238883729408;
B2[470]<=640'd15449238468854400191328073162513620234592984879539572925648245957896542344863638711308240390335761984271720457783803470222156153522328102159395255969111826343636767928171867668480;
B2[471]<=640'd518685488824073592875087465496007266877710926246885494203552746846584499889701017925685772088415140111008276865872043392007284148691114649218725363679954183114397283106256419030016;
B2[472]<=640'd2263398275164983351423063277443614978561929232571972460340454889256188238666521137127948072208292317993136262356146350834434916690739149696505035378188368491165318810196255464040705593337970688;
B2[473]<=640'd4553529601612505951243200041787572321816408693335100160258201843162630320305181178700069970341521772226445285819091246410797571998069247744614327739381795977207506163567594634235604681149644800;
B2[474]<=640'd66904418314804255098633403816660540031157150278154135757739546218974819820271620387327610100745767323332071315075936062428545205535803057551786588871069924175012583781140116951635736039260160;
B2[475]<=640'd17822032882477773123190650999126357919406299756833689319477871025660258919313364466876019280141525667161645387437750915159391026855054778634064804150280100468780968714589389685699904612073472;
B2[476]<=640'd487320984444274212603565907871471043928600791943588384760177109278319137642215184643876460669063574703628741428467668266182396355832536442607875174815734162821253069057462149277981077405696;
B2[477]<=640'd4562440613788237341537427000720154699548964103797852174830255542109114954197663935149845390309439846514280130652583181627043046469948612874582601475685332696543182010475055451209846690213265408;
B2[478]<=640'd570304992370078112127151881131237595713682622601040890173032770444428758678284911950796610673132688096821277023622290761113590138262107797220111936686114631494020456008332843616813760031621135;
B2[479]<=640'd4562440600644452268564648378659059731657694287555844324352998729314985514964878288971112394669430806350460283647408358430983934118916834429343684001402733056537435312016795169740076685266584576;
B3[0]<=640'd4562440617389773717545894380773383588512318796980833768016781232222516145636708937274859881298668050813685708337533492782831266549979452005432190255170743309862982142262454467554132230387269632;
B3[1]<=640'd4562440617386710210107167722064317162222193184386696269888697588394222294070401670535006860689579667540122376959660943495206528355696712807915314373887269959057256734889347058191595776780533760;
B3[2]<=640'd4562440617352995396109828504080181125328289690311840531284477200453233507085398205449432822582891986942075238032971642566488757651492192742179643661636468720004303918804830882554111950824931328;
B3[3]<=640'd4562440616825374766076066951643304850295412187721715190037290685717685955383755449330257308693542311266277467181198239063169293992960672209079964460104380960492628163333212912784581124281073664;
B3[4]<=640'd4562440616825366661561442096994856796179348953282839971019504755069649074991230827975309213440652613213686759560266590520532699240597759297145341396231582040014541373246392863276896841480798208;
B3[5]<=640'd4562440617619083081964503349883540993715371909834236390791425829396777960805845835134978255675466406514232315807652926000260043831903402527740859127205875467870652320319052201749988137257402368;
B3[6]<=640'd4562440617622195218641167846429475481514919384914070646678370577709224544691804536231232932402217040040980925449105750365456473579875756267144088992933221225199586253540182778406565710770733056;
B3[7]<=640'd4562440617423018408017572799172957072983411118629615891178007025424857486400924892504956179067933209319032332514885138264172726901950208893264666866188370688675172999495199308831013232911056896;
B3[8]<=640'd4562440617622097964370018778026095862940087652285257941972756865729903744140428951392199701712869885469340729107450756252760491356366740292237494816504025730145568666858246802838760385828356096;
B3[9]<=640'd4562440617622195218641164101955590569118744120910483403404330575778168410413037486214909384350030112536053710143425387276380260803394889407147114497479389156134342029187562777375680505162235904;
B3[10]<=640'd4562440617622195218641167890677010954422553951234224252407352140508683408105928810659405235818755430994138705768621877439495163644762962524166585789413966182067683697502180374633955060579565568;
B3[11]<=640'd4562440617489410720435043847241305708094245640366300358709025085809616070758331571622430693657865052057873893714728404504620180357648194108665491296893362338269599663737149707314850957294043136;
B3[12]<=640'd4562440617622130382458473743408956850889722789454823982453188583713716412587829692527359936591661921445003835918213157718917457883222936181907546491203786307801154521049859219645087360330235904;
B3[13]<=640'd4562440617620120460856729281207985556832021679828058229950233030491772366804340497786941677833741283066924095121409179367536206409391211493117661171901377105768459409830656143073495530283728896;
B3[14]<=640'd4562440617622195218641169777687241788226240458696872094406900431070763568034055554504954837890356257086649122392494157390313009755847147880404626885948755909633703890316644152424626097336877056;
B3[15]<=640'd4562440617622195218641170898080986982932004351578271018574919206267035804687695272957173488284607587967638624121253714225620080982295146617517569870524123527997159503101719806353153095947517952;
B3[16]<=640'd4562440617622195218641111222301494180217981477465368925045916484374669305583935131076171218117373785615266846105403535177062522218569422752733515187648754839288919783425893842179132177705336832;
B3[17]<=640'd4562440617622195218641171605700291322841833692177519142941918397595732341993199154371357165856516236586485559999648987140393119977088395841870866981136384770286434164359356706585602868841021440;
B3[18]<=640'd4562440617622195218641171605700291324139248654736296627750871353488586392964452775381331267519826327180060145746659124309283084832966062943669841482981494633685292328969741553785091070858625024;
B3[19]<=640'd4562440617622195218641171605700291324569869735988594597308790497682243392263853800445154001762471257901046384122324877723340292145994387392181332128296150468846989498403138524605512075821711360;
B3[20]<=640'd4562440617622195218641171605700291324893045095071583575838345074742804173799404934523485600168954838335400701352669008194841854539134839093600326747107721694672080306017481007645994581156167680;
B3[21]<=640'd4562440617622195218641171605700291324893043969849616156649785304466914200925030706652236435310827432839662371123085046520235479539784799589333059561711527449439485274855122571490886480725803008;
B3[22]<=640'd4562440617622195218641171605700291324464177835142744798746122164507564881499034235230087247642378345636460275030573045322852437555518737587464223287529811136033383819412165188656972214246047744;
B3[23]<=640'd4562440617622195218641171605700291324893227688899054272555570929898820458132527548911662672773302240450712438568790484278450841046784690373616546544449355317767288513264884347145779399503118336;
B3[24]<=640'd4562440617622195218641171605700291324891500156608006950533716622899360775168966399405188496093930390956427598379365412444285511580747395882985000021465136623472672665761794282109995705323028480;
B3[25]<=640'd4562440617622195218641171605700291324893228507248559930207051091059924439247423596883689700810491796267313669353854620859288370645080810860084828524229127000666580493368261312601621089700806656;
B3[26]<=640'd4562440617622195218641171605700291324893176132998833592007634236281449066044272539976094038603395255761153094086755392977546415675305720684618479049976155760416107243009132695742986094639054848;
B3[27]<=640'd4562440617622195218641171605700291324893176132998833592006907397557153459153723216170554576651815526865171637661878755814004365736665475560199363593899433268129320658885438034916193855028068352;
B3[28]<=640'd4562440617622195218641171605700291324893228507248559930541396904235903608900112548505130745862077381934205531027320546803164779078199969021232092371700174287616274702098945515551181846706388992;
B3[29]<=640'd4562440617622195218641171605700291324893228507248559930506872064831862281599019667625753445314731750845524595226071312394302627233375083745002988344813555811559884598870806781934172215940481024;
B3[30]<=640'd4562440617622195218641171605700291324893228507248559930553026323824633319148901729483006755232759974717371008695976462944913812209090017761077942662098423049525831547510056182762691616957267968;
B3[31]<=640'd4562440617622195218641171605700291324893228507248559930568289937034841063850437529528505298268496773040070402922915147935289775413887299313493644796972353080187715593134957113602484526946779136;
B3[32]<=640'd4130256301304467741875357498519697322437522291229897514861891468271695767598401827657168322372345742730896477426174731242611223261413171096383480340087071921390921183642976758696280211555614720;
B3[33]<=640'd4562440617622195218641171605700291324893228507248559930507962322918305691934848116540789351667762159246315170771918000487383409667842816709065323554525606537047712959736417658314448972810289152;
B3[34]<=640'd1140610154405548804660289127462648009681954885257558994374453535105007161580646978404911313685938816587693973461410048009655572276130204398461407482090893048616014519573911595088348319431262208;
B3[35]<=640'd4553529600790901868604750330284555461429937235209273856360327608686744198707174211550276464715999022439038914661060340102973983786365923792782840729823285846627937254942842363779891694114177024;
B3[36]<=640'd4553529600790901868604761652171995120544887342865198145619652518448460242200841603126363293657669029098987476878557325549480906491154320992777636111659877265174057281560211947130110325234335744;
B3[37]<=640'd4134711809720114416893456089346963104717846656952431262360201914325051169486713800280036091356498523804555266781282064106355493171372350180063889274661594820626668986193082648656664834596667392;
B3[38]<=640'd71288134650346800291152831933923017020745154127857782463538388624538024636394173583438591496351386557127824940456529590498079505540361459872513564420139383603342870328596118271636703488770048;
B3[39]<=640'd445550841564667501820307665330163141576785291711463616581527098308512855097773197642127140485555218773504994050105980243667847691142303957408967984205075608555737981289612537997146982799425920;
B3[40]<=640'd1069320931984592715629523790952906552546163565267606351655072174228697907488049661049209191172826739432136238354930781221069968743463765685482807147828266616807969752328793968448570440106875904;
B3[41]<=640'd1069322019755202004244878578719449173697711125808803400399980961466731225275685139834044247881115183383083981623006030694985838822524995892865038547507032293098481906348698083885629568337610752;
B3[42]<=640'd1069322019755201917184091950420014821883227179308801487373859978903901658413211251960916609774456069559160741202467023103094223711539647568255810181623144354575834866425343493621275362940977152;
B3[43]<=640'd1069322019755201941044712751919529492907328396786928086029378017570418778491775223392871222374491656936787516573870532507537324461926583476979821397015921388889001298618229679374709846649602048;
B3[44]<=640'd1069322019752089867688499313578416710393040226159502899500045327003409461582156103934683141732836888914849710101676823397170781869543190254630922324389156540291849961637599235274910006025125888;
B3[45]<=640'd1069322019489633001557102370131082497919271291015910102551642643613034262381396256243443468247482881879500941157273242396342622946510293141809357108370913828453357497754800619993827135727861760;
B3[46]<=640'd1069322019261393404549707279198668952493406910713075027458674307890353789631837803280375368474435667795998413748028522056305505635875652753628400474220894091423655430334111225028808758785736704;
B3[47]<=640'd4562440617606634434037901081094203584528799661529443406310744539396847854447293582113122610448505128531641174171450166452184489958087667716457759279159895745190956001322875155816514404526850048;
B3[48]<=640'd4562440617621238793208081109977060663597614844749510444694376221416736109883583712835255958042621549591292893045408024635838002974856513663713046709615315284797045341328964289334675874083176448;
B3[49]<=640'd4553529600789868512106822691272881919815143729842292279509175077456661587715031747581597758712033774063278368961898537586691117024454582535957817129772628364350329144802364487494959138879832064;
B3[50]<=640'd2272239674660566582753894284570342119444893314010740735962078447244696087743479007114525116508416912885320322521578510000049258346368843357656643232665699675243176698319386827388097790614700032;
B3[51]<=640'd1112206288255573895653345867592020210623164220973623738115347242633725211690265185132760769690508599672090032983193759557506900372069235209446858697434122803003820828039458018892190502839386112;
B3[52]<=640'd1121117305083755107281780850839391023435290434115040314177143561245018319483695667233527035955937204837294312344741451219230567711884407663446717686378784823148789781692547928100409189790121984;
B3[53]<=640'd1138939338745843414814613074872380683976925384876972421999993211198237178479686356341696179436826448156649160818423219803591134032731948318366920636540114151688146216905423806354644253102047232;
B3[54]<=640'd4553529600790117344921589832685408998362600250318891799354624213963908098282082619054623144374519554473011110883380541885810708756733126539994426455026381120269277613183732467438072706422013952;
B3[55]<=640'd4268307444869735576190904803957777642360099610863134299823347887635301778743041880362624524576124915594786764715071901115509731262189430046006908206920560592779980354080155128633063509485158400;
B3[56]<=640'd3483711557634742818438480147292515715571341681106500274689312627537184101023537737912629272405703469921505683281229909525323696068613267363541684354225698801764305345147396875350972186706837504;
B3[57]<=640'd1085194768485934039931208145348386699020705216273416448400287385885446796267686382268652429042524421807608948679399416413007417227256267503945039349725613639820693076715779409949484916865499136;
B3[58]<=640'd1085473237761914616632736652451698655617302377905694659194509706157937066947512628067468740505111413359769674355310504475531150177737702345543785587403603753734684050581568655685314594140585984;
B3[59]<=640'd1083767613446549873975995531232966125887263386893058211833785115870444980118259881068117551666394467818711484712342686886680881297069846370677761175485495757248692808031458201645098012782886912;
B3[60]<=640'd2192945548319513082766019660157158852429167473786564288349894746999645027352376813829659540269178858859318674085103635664404485145521987210877078477953084904370114478162000595647602540675072;
B3[61]<=640'd2303254190272850116944987996405993149695962261300433629919420632841525506404069477077651931298283853870824788924468958537357752260432733351933939297024029470210929763891722787478480975313240064;
B3[62]<=640'd4246656458662097691024507529444571887005222801881057486403213577534363331549692269801928611416639165386139875518861264562600578996470173705843428137685675372470000401386108596851577752387584;
B3[63]<=640'd516838976215012766931893277398393213108944209617180973317707549104887471321122942596405879268844238693052984950758033079558383292384318069067938659816897179757548258051089039542195482666205184;
B3[64]<=640'd3992065923100418216662124548319682086248335319561263057626597195448298580988772832132115000271294546872120636851045218413286925283736910567146982784707414414630265206668637395778183094276718592;
B3[65]<=640'd4562440617622195203043898162802636645702788275468911248840059282983606541841761978066005193446840468714918805876895049460034511791733551133733997083674674000447717783943612640007744600882020352;
B3[66]<=640'd4562440617622195211715920364453364371199157918701560358145103896572429641244728969359355874061778128240058845321051708256272800364480583317399586173993345631281666921341321024350047194235011072;
B3[67]<=640'd4562440617622195148893998390284812719831517579729904580522546920166468476113992849625871710930227512159610908658644910851057054321713815583798993360005412747354620307352599977128825120255639552;
B3[68]<=640'd4562440617622195184633241403148417891574131867169599931346899324434709756081777911708883120894503674471318545843871114669994059802983528203860378811758061028408418463493590491677221044661256192;
B3[69]<=640'd4544618583959604938708123607400498570191875095125611562707361680429806012126998155933809677536563932166928261133561604305760047223770927821490471756362670882920198311658153112935396467284115456;
B3[70]<=640'd4562440617622192145313602900903351089088902317221837753297926604658234401545765622088039750723913865372965135295478474608966368230497850844692979442255837616498469379759766571168944267081023488;
B3[71]<=640'd4562371000303188484122619171665219381825390639672655049779857968337854613011126619661703081248498568392091724738929646025743856771539476374620043377844847375384110753677148482299520373948940288;
B3[72]<=640'd4526761741637524518498339772240546865570976737618614836631739277296470434686458603281034859463464515312669588823448223006296675530941839131883636444076212317657109238832320005850406295986765824;
B3[73]<=640'd4562440617622195013047775381182147387102183885669002158439447884089396761433198106352661761228961181987158972155002225417731361810739407559207293590678815727538584355187639032737501015177166848;
B3[74]<=640'd4562440617622186908339682109387946892008522247163848846896661146331247417883683770912571610608777969932880575974869778963922988950471483500552192336302581627856949723057660590833697437327032320;
B3[75]<=640'd4562440617622194719033760630029132522678136048372890682695298474886278254972976043930803043176245325646767176217577326619517704090932419196838688795777332675864562934910103217828060904143454208;
B3[76]<=640'd4562440617622191172315803505710114095082040482592129520937696851182674640165534836677764985865869282973745950218119190028582987841433742306814501950313356656791440509067974692804106646563323904;
B3[77]<=640'd4562405808962694037535314009453731914141092865986324148766586898556310957612531960618821286510927125278176773800763910445185682776752167548792268866688804314533573041035039630632902788980408320;
B3[78]<=640'd4562440617622193239997959820864018840873060350120987626333092164544513617264644154663752363718181562133734029935624764436511461057869179229441492022194022516390090003460368990742817154202075136;
B3[79]<=640'd4562440617622194712108509388782205568990769363150757624034012654575905585653273800057721876636770046941493713132192811761082650846311667596763557985223184350274404173551467792018086269246504960;
B3[80]<=640'd4562405808962555928239131427910705577818431952016409241825385697468595540083506308072823441678115829134247540333444736229196282404080671243879693340495488219971256704299915624270219234223587328;
B3[81]<=640'd4562440617622194207554490383648956085558922578943419421474515515578007360690140295186286684770459589262731140651639964304524652146354501750444431551958924846120749768916622830349941407077105664;
B3[82]<=640'd4562440617622191172315803505710114095071984625820543150160505039077691097955937970177725992741637884763433819329019337238163080009580829675284055744685412952525672319298649739112216525640040448;
B3[83]<=640'd4562440617622191166379873870362803539697897139529600498029798663773551451131899872514971442986032984348825917183805132589851806867883386704376941760628436999810336547376010534922518662402277376;
B3[84]<=640'd4562440617622065324671604354775873556008498439071229770429502206883304014488946498973409997793301426517347620367660020944196870282090709341069982961766959344498198740960705609941509508327014400;
B3[85]<=640'd4562440617622053136229419760191633316515531705070178062345483234579784466010107460260213230515772852490130349245267054845567991437715644224126234588466565848771018444516782885021351205352243200;
B3[86]<=640'd4562440617622182808776445092312018705664110716195888412113756314530338310535973592482010399872565255813345775267729970154097192632955778789266720745670776664700593302147567933329648135094403072;
B3[87]<=640'd4562440617605564769933557139701225202593788397748780391631933337594547493197280609798721369961432668935300803063783083064967010891687979406175333639917913873095828930865201222846264671767363584;
B3[88]<=640'd4553529600790071123627766334716979392222595498008765429720901701109305058265676691818903727237294900731752254805204463559262268819280896903872753507387615821954630676323516180328442425417662464;
B3[89]<=640'd4562440617621623058340906208168648796784877389645623944843057114209259699861721608027900283819509682582772477358300136223123391284106192191018720344398212275601462650951143119792088340632698880;
B3[90]<=640'd4562440617622172044771875181710464950673740000257311954367885087976182517329639677851483332949030480802658774550309566486683802663341091634841175391427864461397556077162237093912415183371763712;
B3[91]<=640'd4562440617618021516137669761408613419276463762303578346164182457235332071376474260426936657911766242513110746153787861768374612146967071127144703686254321509237057995649025628303132149585805312;
B3[92]<=640'd4562440617617539073456556323762960882388024391471237463879550352682787214756455500032096081547969658518732766770866701088958123224682373187418823228124987697992188095761137556956431181580075008;
B3[93]<=640'd4562440617588492494154037549768781909411790191710175156406551126036914072406373712598972468186315203121477437837746465884052444828061962982005020039453732472856250002747868265694684158592286720;
B3[94]<=640'd4562440617621704372662337739563823226870176690019848196980362600723932699976212931489955068392955732854537756708196698388950699943627053940118591473120150983600938969755786223320872063942524928;
B3[95]<=640'd3421830463212297823284838823246498782505916666641624205416163041991521232029378521162955489623852153463027839940190048502136999185833815016835794360820799062737403815316341255518868696773689344;
B3[96]<=640'd4535707567023799180834851612184874323398520952164865741044080081533716818520806996668601744535925174617173887951696815033945002407161266397636489646989810211482753415699828285070131686228885504;
B3[97]<=640'd4562440617588739749119738212895648408550707335854308144928336950308007352991851568259394072274899393123298430721794733457463897114834603851197838858100943313513372016500921297392241190790758400;
B3[98]<=640'd4562440617622192176353568315262008501592687927677103854643771122848767304950719035590513144042851583388937221391006495010100775868761840909782617866762954190745396500492914534569253249340145664;
B3[99]<=640'd4562440617198943614334690788881819288193874048908492266647161990704444739510767716475396906176372981994960221346273185494355170477284191003029022377629580040373005273936463863782560993262960640;
B3[100]<=640'd4562440617223744468520799097790408439055107383172512874364972564021677497901769949842028071989107438226555115361281605659524862202720308457394757547061738780003598570971377091800863108012965888;
B3[101]<=640'd4562440617356528935808690688324738733190325758822075936380704173176217420294132718965997828693969966418829487211560233461524650086473646481410996494913406089342145847746011985510684304689070080;
B3[102]<=640'd4562440617555705618809073554549015240060760627542956978636566875734370381741021415790214546916011406338646260710043485606637673817165312453826716337329690987690689135443569709058142412768018432;
B3[103]<=640'd4562440617385600837045042267399942933985896013039795415066521224270496668670369047460722895757036370966972140570171568865287608034864886647703313406482911824355280225807708113169816018894192640;
B3[104]<=640'd4562440617622188724857815787572358435166539703896085807755864982696122502086043997620709264542243448180592591923462093819259788311414089234358501835863287759074796809973363495340510176551632896;
B3[105]<=640'd4562440613904221742288689604028857333611309964165992191370462901383885334453481139344881034723748952232140638407711821892426390691149169594632371944064050946291233427938416862940975861371764736;
B3[106]<=640'd4562440617091055587507825267102567159302155073483484396609353140074707517967346581172223401391602309978496782476808139057974668608144403692392106858096176410954877775197362706426655725016055808;
B3[107]<=640'd4562440617389820700552683854007952547500730266372002584300653529837721422173305621914253838206620678007034600595050627462684387960315395447235357575660861146846046064159780264387292270281359360;
B3[108]<=640'd4562440344517669292948653648460725092492310375198274485379633900634957568050737094235554626130736641182863842282439270711454883324430004078101281699193373265916819015286743046718494704784113664;
B3[109]<=640'd4562440293096866158350276808296603854635680833590507866468813560179307839492278227064048270862389546047930081544918385881783629436088814253727484801630245080956444729060191748628252355962339328;
B3[110]<=640'd4562440616688546142778644166871153134916120343678705752735946153424278913141676958653400844236474165037400823355495241938858076741238619577789765961011161230516511954429183603382717549815791616;
B3[111]<=640'd4562440613389681233859963340331659775252724628677466069990614118083678410599783182879928059744098375517050642091412450615673339583508004552494461946058440413859586108486367982910734052850925568;
B3[112]<=640'd4562440465293474632774080514497330504392310568891737472236674760033507346254572789302609557933138382771764198201624799723324286480752862929939168240985757587602260024464536389698507307323752448;
B3[113]<=640'd4562440613447778504093324029138157483501348493836518530143056750844322907227302327797715191647572638041283123362385085338697822731585857964931469148730387266071345244485616376001474638620131328;
B3[114]<=640'd4562440564724154537504946966728388947822523180337507056886079272518481847159816039723886502921090051185819843604119272290756171381237982529817573519127278492629897302000229956782030002411536384;
B3[115]<=640'd4562440562798779313546098502740140506717497383391445522776395902927252474589749512850527771429427648090705495072188276351453444973137665631365480056847556074304462350421731414293950199458955264;
B3[116]<=640'd570305069268892530110956980870457949978027066677884853628664275891262447674772468292834709286430977085585472415529051316714789585331527864751951816145147177514440938615486964909851984539942912;
B3[117]<=640'd2263398054257340526483275095084999776195303268773805561665436510550908509111760642749744288283554248554190018648349508702447740320417604240686950702933463376814955421550927629005285053423419392;
B3[118]<=640'd4508974244720821300697537326897059842612955039205201179944932461840705104005049253795578997293668387515583491400567350471724639291419780491540166824986820816623007935901550137415008698465517568;
B3[119]<=640'd3700288861521650630734321365435170153109729782146700475216795771487430757327233021554076783358092492504481883762402616357520496029367272456953161599463127884943177462650004762972324342678945792;
B3[120]<=640'd4508903811555197034786149829670942545643442198278254058875655935630198091754909294532131964390667238673633901831356512833429421941368519623504630586362028950695408492705888657172753346776268800;
B3[121]<=640'd516786219344605209315602103810024896985175702522334732211497573471395327611881302298366082384583506073024836052820213082781850261001935918732957556257657181542356962545064678104724335556034560;
B3[122]<=640'd535721586225799950807669433480307839184934613320045521453051324273679413271740990963963140786768582888644438804603183361176414301804043487837244979126937674496793694194566162094682264850923520;
B3[123]<=640'd3528814878189708465844153808838032350102809656170763325178478462978167169854143580144115218288180555417836031796392256669973871353223020022434955669856101239909211639408595800369007011660038144;
B3[124]<=640'd2281221124647350156373925685477879573183122097622990599804364755338726366893151310181666380881709014503966739160001204171389054685432104014646041195382855002837300741438206018929959732519108608;
B3[125]<=640'd4149484022419776909770176489211097571683260241837105470366801491294712732556864274495114532181928296001582562885393949653509149966867035923972291185326250116055120567510073488703488;
B3[126]<=640'd4149274297844557014265536118697570381187984623970874799331916045969488492103279085941923910130297590134351642767764236446563863335745533013491042768610734672482402432559563854053376;
B3[127]<=640'd271950951258161129352376002374797560993255412520772679893633604060779576817367084320589165435393266615859399704756977959626788165957499086434063946727743271719161668045372682941147119616;
B3[128]<=640'd4668038561510149668392577980101729724802936166865198595859860916371318715086518922581653488760192858894600560789469878504194026262432592069058256555587514338481488050843524295294976;
B3[129]<=640'd1037252259052777545712563599245007398026653044043970926029670013126698176567225633943196881737139652756321622076236227236978382486441996538743163300278539560612173160096286839406592;
B3[130]<=640'd5835128646222480653803919138116051217993296944719191509362539090363837729797618011453827321923120692269436768021235677892603749586334368226983809457565881371192227984749447169966080;
B3[131]<=640'd5964927146254586310696226213630479825114555863615227839528385993144089132133373612741440895645773242802847377501626868054209286632819092086530372947598168791423836265157924782866432;
B3[132]<=640'd17822033664661433355901034324809383145963913004781992962094768536722984939907991638856927077765234205626910552021470631448418817570908071396731535860184800728158884738447003491607070101209088;
B3[133]<=640'd2027256329121311866520621834962461629140928243636214983101958916732480029090276280856379094679238289116026991359164994592292948477818887552824507744719004221920103834595276916553626233442664448;
B3[134]<=640'd2192110140500757390971126397856041664818321567549327526951673786260913032014260965705300064902219730040183297614448133627399886599705334824086922890053791830869382860226220282819148039491420160;
B3[135]<=640'd62359713491638894849665984189364166218191515761413184427399426316975127770955696815225896472338578738141004472116925489010564901436824240073180400017211146450610042454596039752341025070252032;
B3[136]<=640'd2415338073854593882725459268766774956965391857757084347935373834269948212068444987082233740808910603235299682114586018780926324232523613043926166213764183137151754814852735519623153443944792064;
B3[137]<=640'd2833211692783328285677575649050986786505494419014089304689624390130340198824878967579100216568339214651113914762257704194757436401746079410342813949674750852209479071634274989139441220944134144;
B3[138]<=640'd552443966124751700405155890267171051322616722068683577022139166760150190939389776254759217386631062411481208779922829027596777583265123142897313502131619632184658493520433347085004945804492800;
B3[139]<=640'd120260860270400346897983178461431676810448469138068291823578218915119969511957075204997721040591363568852516449373079884390294012155617686344742166394877006548221173735235993313494495062392832;
B3[140]<=640'd2352361697470001558910204798084690820672895640680248098407888100680269734465448924389061557465260304757125159628653797533773102071175124692105604588738785222134086234760140180806238930057822208;
B3[141]<=640'd926732220245279389461415963844196368447508320109620552115849290720128456323321008742537822121850844050700162734088492134829498695264830461002381704695585866440686341243117682110833232919396352;
B3[142]<=640'd3199054905400710516344753799794704670198713682234025365872443233718188330610302040027777778134666877484365356932398296605828719312029351033721903103102741593814808105511084711098080936272592896;
B3[143]<=640'd2325217344337219747127307640808236546544997312536270747071154195023821286869892372431055227006754673107398469369444717646354739282594356739335194098253617811522531583923319506597106729485336576;
B3[144]<=640'd28891187351587573212852249113374052318794618860086859711809347869329556886093818144480153065187513403852344067386902250604031889372692226548628417333361203696900225893871712083829525925855232;
B3[145]<=640'd20045436771374820350322774217224900799787073790513900683482145813468605484264002839343593522026788975831936649204660633763775896128911052055980977196504946976455510589238863807933996244926464;
B3[146]<=640'd552578332285396745256573892364648082745582688651760398940986882097767972188536094919176417165164209525827071960051853598920908516355577230649397931727864982023923048592427684336804084842496;
B3[147]<=640'd65265331962930325030511643117131754400174817036194120382635802494114946727004643900017619543596873455837104802796089483542696868847678054106218472022301912742763424493798883050141654188032;
B3[148]<=640'd55739878302661010596654817145521365141253901997713973229577217095349763936932494420384449734153040618674558483427889280135681317239017706793129480134568157934529004940233679839119504572416;
B3[149]<=640'd4142876343970783369778788011109255502503296588028076080914517765744063919091566350797658658337619439225175764548508564068987860029128666980163506646839645645145005506865612950066752913408;
B3[150]<=640'd3544354367830957826435916813261738508073876204143691194686200409398577201006900742475842929711717238368160491593586998523610287143748266555682750432827689088903869480443298420100379443200;
B3[151]<=640'd136606202043131169187186979284009534066563627883773405025622172214256203903202580374353235918153742399039677791060347154161263432301103598967581776508817806680034690062036523177962635264;
B3[152]<=640'd203957118917958345985782251688448326359603027840423446575827915515660954215300106936839042738013883008969690943532957121692635302014793002784458808007878203739465415080505562212675354624;
B3[153]<=640'd3957286423569672544968459330289517826830455570792212428899182648776159024422462000059779086755040759128487731188324602825447460234988622411907135651497388058841481025863811072;
B3[154]<=640'd17822033662586704030194075252635024948777301476198695249033444878955351754277643828487353070582929445051615489242068055387217329860896566133509592807921538492711691317541046107267221052981248;
B3[155]<=640'd151487286131986951113605953916726553518688507813080065231473013272523710540329933872838954343718577536767128301285061927413693037330820024888646650258405642462826508082223302776346717391421440;
B3[156]<=640'd441095333149020827299781851561451153218203840332950134297721098886935931961906366998327846965342548688502950296523889413038912992862770049063759611597643413865644022270350603547847128185307136;
B3[157]<=640'd169378937113568130858201078401979411198135594035656769282172479717852624673830086421179454105110326180228055240073308611464685086432246116186364309026608057593439722566583778591451290995261440;
B3[158]<=640'd2765130293141723204865171607250113771315471400039936324860479400807774319115230889788713271456539036800408497953552874625560823007764684036705568305111784916537267258612940778627237799192952832;
B3[159]<=640'd444471773120253073703762079639128936329317165086116780864792382767644041895191554386506669272827948835842127503533559755664685908440705125665049187644052125951448621375767462887674452956413952;
B3[160]<=640'd231146937384251427656044696486373332850457619481468097393682315260098874208142366121117297376265947178594908749611425732411200562455387760127566871207817545157210940521709401958195221495808000;
B3[161]<=640'd2423257043893733511908337454181076249636095307587050295484568089612035389327852057130264985145309458455018068799411571629250557474224855121467554406130626442472223826926197055888464717497237504;
B3[162]<=640'd3559414953195463507767481378780504653863763782350409180868259120480897511963161167143745279728636328862623469866529418618514463728706362959250469114351175928702874759179286710814528421360566272;
B3[163]<=640'd1962332740370230994583428723140603072932879961024272607579659563990572712765605437614188871065854915911313556306035457288955700865786103375186312129136548069220289152122990787842588465443110912;
B3[164]<=640'd2254764911765238510093064297336543451634712505720127369291101752578896474926792157077257100199968375626844113304193317163055593782644187213424765582606434757473695345539457078990740121481904128;
B3[165]<=640'd1844705986147057654310094351153927636647869125890232189159683015257118038061385497283603795324852220485770681298196900924835419935520757547846022061145449791475408292368947069221703021815136256;
B3[166]<=640'd4055765090127893613791298721641192853801124125977823240732925304107877311465752865490429023613202985572555257258415977455060465027462618739246735741450335929747608433982165111948007652578033664;
B3[167]<=640'd1759925038197870396791605963444704634449788721020281781089103022050249338703688532232172055923214257377378764375549945766637330325606048656099755494435079849697838857857702968449242972502884352;
B3[168]<=640'd2788034323106867757788843427959343884663594685999487210803437524733428291038315145966341208981225909696276765682641993627265490205709424530941566686921944483019794406845840186767727160920637440;
B3[169]<=640'd2352369140841909978192463885775481748098851062284868349533123605930913504078584337520098027762970513826869720186331523745052311571159367046115550813744978561322734304034415663801985753572728832;
B3[170]<=640'd2919332599604657950523467283386592070994061995765547694783327478349009716960082162906413259351047218457353602742934364301927559055110440838986999991352390096369261042515146761702120449759801344;
B3[171]<=640'd2121935863959291809606478946651085778782728232980357816712040981825708858961733570757745953003255302241166951638334635516845760856783661119202548530379393033159216994097721089983789472003913728;
B3[172]<=640'd2108569342849523215771215581857322476713222674389987622098722104219141594864285000607944784069107672830056757563607627434962881617732664023712697549459927850172568117579348430799241474905996288;
B3[173]<=640'd4330614778609847445252594321331801878193930355807064516190118855385781260322969906288026611992027346088275970694145449749361721744281037910978163875560208174983880955440293140772413122461629440;
B3[174]<=640'd2325357536102453583107980004664894607617443525381393387268987414330353331164529923554399922223082335559975130001778870174905098807885303258223068489363596228913413144829963730153718632339667968;
B3[175]<=640'd2751415543419707459557821055525936755434388144360354863030860295694416473412692961899325066612392377117997913891640372467323299086195846591579547089903540594313297790641986258244327716654399488;
B3[176]<=640'd4445761854182069126164490458207128826606678324030339511023604488221673619691187616330337488020644371032951708171521420150675658246900138080085190227418018030681826667826221598512058848790969472;
B3[177]<=640'd3412500790041376694044961734282889415208645568620677618434040585637004385934775994456864517184325693973668495737626009445415905388945528075323006200438623836928752560654721153328263526447283200;
B3[178]<=640'd520754116422216666599425043224272673039834091965917343237935213760750825921751285748092361509981473607319723773382373410178749181597483921920646438187011465443789282325115556794824119067572224;
B3[179]<=640'd2717860624481957746552643086696880933379653045102073751184576112201530083437337263028340769258044465873381528642327905662325361316620231199186052934942308885537420794978784435251011276813361984;
B3[180]<=640'd2307988320301490463837404631487292048475847794185571007225942163249548284715862862182637772222673442959577306423417917108173897129544161732999521854374749209885077635862847367037139272058534912;
B3[181]<=640'd2299075145439934237000750145563975078528264361785210626432536271214465091287727577735425783034866340785416024669104139510685661711325455831283471027549300669645008814974124266879289773810252800;
B3[182]<=640'd3439657011452583682920890811355441940047823779738865666524829467491289521163493252129076840221624044450546400634965048663117420820034997592080304513173186386265979033790106663085986575896542720;
B3[183]<=640'd4423206992235371382782118867706178665102743318365570575654022696599935375771687783334306975131275113408270799008841767456852006804353516043001195401260630194143385461448460275745819556438867728;
B3[184]<=640'd3992205300909150968709054452547368803377386850082202094576674030898527928331572483954479465860031977721679149976528836208083640940774485970941148702312728890049522909745344124401419712133594880;
B3[185]<=640'd29772774206721124477326526366958437718604382046252648821361723350585345797392685032181465749343730488489279895318371191268011889610513147856595741118183767149091856539207806972445320960;
B3[186]<=640'd29747877113307838519575451974533778286437267951866316128355502672531392372209637797441741564664977021257733359614348405302624074226066672831877303573049845805421328066998785827355486080;
B3[187]<=640'd137037751662294792454872269697730206666810856334081774274151737685468227540195547578361954647665008716879483425847227540976123457633476640944313101291967539444238629563913327484445128384;
B3[188]<=640'd137037751662294792454872269698373781447049297617563229345634808511348134668048997794358421684520731060527587396222640128834339757978767127142135664976665090673240312903004958711059840192;
B3[189]<=640'd1037378892220248239628101939107317454875045052981936375066313568112063767622947435038892346784857940762006078738382202469619147830142921363145376428445505773909415952716475028995264;
B3[190]<=640'd1037378892174945948489521497142215271621506785802355806951145337888213082956936844798953656373806360051831966488893239780554371441676194721608866450193352683930699199138707300941312;
B3[191]<=640'd1037378892173073709317832690639903689080445645274379159589066078319931950097335892674727656294360185174036279366257409468659179860911007469195499846342424594906745091680555136712448;
B3[192]<=640'd129672361523285322225588505067547328064063962646405655877971623376880457030426661697939314118156564374125075265050530678989389843196700444697084600594856316323993629398701705231872;
B3[193]<=640'd259344723055062002320928914715534850256675514271784656388323034532732119813430619957806706800543812856148756121349049040333142928756141380727374564552800646681559446631918222691328;
B3[194]<=640'd64836180763758136758133313844630076448032576480075340703960640040236434603620550812919214569101873197426212932727611852362082439647009997664758135208914143501114237005879735993472;
B3[195]<=640'd32386432090483100387904537910724068518101688926371126623255887323795505015107453184672582684422626831133336445667851635184466126928412199147524045898479506991570586724313981680768;
B3[196]<=640'd32417162892877204328381477545713915762137676150940490025610889558631018727745090367674222076599042359266454500281241682523023551647517798257344926848558449852867721740727370005248;
B3[197]<=640'd2527747619355312476165093262532130435090206601086157711980497579844457211984772729708239712968333571078963855262372698224690310552088388294412392582990346432825935312552382628608;
B3[198]<=640'd1560217869743857191243159299263982507255475347454016179293327044628371220122183058355089123386749347048211443467387251152513457400131888814334065348399928291324379206833402898278219776;
B3[199]<=640'd35739792184470758683345451861935316665600803388974531410166516063378853802587296181151263988720174897009673406391387468641041897999273236282574802775154463664442815155025342338195010871004160;
B3[200]<=640'd27010465850996689497714896012397974379118583570004922998531775943678715385374643576536109266847193135637968559452588390523693210628223090839778243032345038052724403377451793916580032583106560;
B3[201]<=640'd17821659739364999288203640158430404462747930888584233356608536208760884957168892864669780649728131080418359577207499549265796066650897804147970151282755239884159687539246357304372415088754691;
B3[202]<=640'd1122788120741924725699120114123695224614032204684836987257490738183459923293970890010133899291534427592916215908450399523913688043905047016565637090730809299189419823378216382875316061766352896;
B3[203]<=640'd4562440617621676529196993750341985903081947016366138555530828986253476097314742476577008903005097879219906859807092317717726738374877015795516399378591659084892846808974012456521026301295788080;
B3[204]<=640'd4562440617621939101086161099089099035424043391822426738438272057269087602142084406670974467590834404358467128229757650214404793830245247270564851241672769369657800095009667588644701499005534208;
B3[205]<=640'd4562440617622134433733108570423148215491086609719624115673167265165160828028874850816980928292197806719426492203654881173240323678290848222781069770925993008719452492406035487287916552199995520;
B3[206]<=640'd4562440617622195218147476937134836571358200899745524778826625630990955781611413272120489557048103858375158419210165258145539938389633756919989809398210511611291606820212682249192564810489135232;
B3[207]<=640'd4562231765665211780255515544828231678561349947471778127829690093517430510608705879835375932420181204549882059859143280145894001571497738523371519177407142566958830967664454628211355472636542976;
B3[208]<=640'd4561988105048731102715940566049676477766882364359381458626836749299387306420760289297697068553749428129114615686005459801211601225633075296173768261414428702512534573093155170431779023110504448;
B3[209]<=640'd4562022913708228342610944937393528464486427781797051755055416829746454548391139133051738837371202145340204193853448651520589758974394960739598706572340028992035939382198316596048987896810770432;
B3[210]<=640'd4562440617614933566272085434083936534743244516820928900397884340138321737748051022010092147205910675036378553792172383569159673351723416396166765435818040220432589640520331727640632030507776000;
B3[211]<=640'd4562437354163059549667024502324582061322647661059929448841362212406896633655581185439613065517945716397878249465524567589002339860104695843931146300010052258493936573170088178368065975364059136;
B3[212]<=640'd4562437350069562440965917400827242060710079186264332509063532031006807002467557351825411072989957573370848200510076834073468993836649542492667264626786335354955305304823160901193027760411279360;
B3[213]<=640'd4562370945069126394871835508710147958698454784285501121422632857462163299128234168080727070317447389365481094991587485265278792310541961701532743140496183142703239714556110497955736937495920640;
B3[214]<=640'd4562440209708291702182589935407462662892045563695564568441107143584687809556736460725229435534065543834072883602834710239393949796641205604442572565168087564009506033471162108364047001167073280;
B3[215]<=640'd4562431507543601833483803649510361131878863966155168100999700815040663837485947612668401762578942720759941704334661591030516656008706375968907730109707445849230820036269576551570793761920573440;
B3[216]<=640'd4562440345679542936025416775056776933859444510311755394552563785792439201358996256514926021452732923797154276637800349506919576351986547322664342093880153504246629577363373738500946398038917280;
B3[217]<=640'd4562440073736890578228465903941263202840320632635627469084473296766537990056372088497071595989920058852299285276897409102001779182584757099612138762586990158929711317530734369741508882952650752;
B3[218]<=640'd4491151395201239137525216496628733768207972177579359303042027647095650311893903705909486254780129761982421237862038318439189649190453458059195248686086674091073908315841959447736496375853384784;
B3[219]<=640'd4419846943991753006148812308787255161231748906774562494077971724536911508662325465841648509297156983148704768038837449067305159769813252343572068424535041339606517948823295825300423667600557128;
B3[220]<=640'd4562439529851585930891469434372425374122631488248068265336226058529880071550873367719818453675507532062710268632187792844877627416191553405057950846060123305060517953377516003452429275470282768;
B3[221]<=640'd2254225105600378981269895762804953468963313981575921273561431678687692703565126710777577925971317927572548200572368587323720569458200366476924450575787141711414013130504693570214259039709493268;
B3[222]<=640'd1391789441337630116729995841267672119691743457094854157118814547993174420508121512144466419567599196326290233396228335194565718722486764638868083445295144967622804110908062796374958176269185156;
B3[223]<=640'd3537673682023459964456121963466691434364722552759812942359526893014362184437420183926576847856261105361008962750841151597577995162052848109947272208472676228722248122216058207346547366404690014;
B3[224]<=640'd2441618611774377909976422559274630686399090649832681570852550342136179797453815163807975042977982785094686085899317609352850714222427934593972872035001872598428200683449935049781303468045679493;
B3[225]<=640'd2708949116713178411068678708074700233812350180310260866197050926122449439895242809011852814169462954433220668222769307852774808604230114772726193610953292333406262289462924141277844055128445826;
B3[226]<=640'd30191699193445311987943138313241362376184060498610189944709039668957629008863084446720352559791912430217282066261389922650916476548647028332491760334418028572667476906147;
B3[227]<=640'd106932201975520200436906233470856573499786437911280722771753309991635291782557667884106967451079678799575049520824215308935312535486842833778587526102960118302525241116656360089679029715857030;
B3[228]<=640'd35644067325173400145637927131895956803651227933836368632361771628538315896628035720279652668547847674303022372941179010882485943350352002353550518224521501346567021588715887654383408587386007;
B3[229]<=640'd1886981187735255591504226758544043255222984944709942280378844813447775116574742538541127010671963503083928154990852140776444339590873302392309287147570113989285923805863;
B3[230]<=640'd471745278396285916202667908663030549739228095959707781719563981944395281973396440828347532390768992503836064813638485975609278138893973240583890515827962905811038888551;
B3[231]<=640'd471745281794360757762732804512250717321341289047986311718144342363917742562501983789175558826313708236530542191687453500504281754621032627570543910028731866769724122851;
B3[232]<=640'd471745302924207955235575681461319933538473933564765530156798496391775259901058256517859843582254507381360698132929880864294198637640543653113937632509024223069326173996;
B3[233]<=640'd235872651544481548311833679417863597641708083024137003892391277014859806953824226339248133163350376458775444379506081272973789825256093852599224908246729040795700794225;
B3[234]<=640'd88452244276407444308358394843498861821159957710677319459217929661515143852439266677851088654364316312293326721972832439581427168585734671942033829728825497546104994887;
B3[235]<=640'd29484081443703766887508063699691608751761328207164680506837630608000812212138588657742403992999925640205462896482373730304928122598087654167658806760211946416532812946;
B3[236]<=640'd117936325775250821307755388847246821053710303984998163363407786491277462889309992722500008768936499110867844703645941872512664128107921795147958692955617607983577910771;
B3[237]<=640'd60501335122920126982099507766213142260124421124186084687235838068715307702226402259916828759519071607385226158699412575059079420516240986870342985723364146722218522458812;
B3[238]<=640'd120884733920064942807755575401892089616082640018079597553962075685169138083009595212663916690366788811099589708459605794397112216426046886459162833433582838454836588015795;
B3[239]<=640'd7312052198091682738736292230276372680228992901596075563528635844937543277413149928943861185097127519661472256626478069696908995661509726636418780582652573104073861247875;
B3[240]<=640'd30191699398572304002316576762711951979285741596833018889001546975312069355318684326455127359399035199962399436162076034714038588555278018152511420841378756975737793604321;
B3[241]<=640'd905750981957169897722357239551990334672016331797680774605006108045867184789044248126246458974375588208123057755605036722556077059083770700639104461877960634762589940514523;
B3[242]<=640'd61832600368276133501717822324969200409208822716577588155690881465082795851029578177533083595106212316133419629822772824368120254164202471086184034769934572555300635052289406;
B3[243]<=640'd47796600084677451207185408283081848175739346211360336021454101540647640673472965471663010594186176921874674293587929559363916145489559986403235251508470063430850533291657269397;
B3[244]<=640'd47518353383020208606367342946934745086949823439462807781847906163408041697447549479364696844146313810522925685167957051286974934731975981845094330463920583179797482873796876500;
B3[245]<=640'd14847553163432306560316190012978209727521585960616301873954728176181635449014220258337992510648951576865957842050531724301606414861134906124064239282068889396369633609589423439;
B3[246]<=640'd15550898992621447579052420033119074248821817947591158221051639624614584616759128643886224774878412873986862115099879362983401376429349671806786955778177426870305501423461936968;
B3[247]<=640'd1978643211784836272416981128507464535015767628895549450773413448708496199247357335626437447725876630253767421024563907032690330313179666151839887423380548757137068122825988122;
B3[248]<=640'd15595146276120956070110835048615860896207337179439167361127600965977438871160838078482285422780789174765530130227374361768445656609002604689703307699701090889327969493984049266443097139672614;
B3[249]<=640'd3674682605374503597385776202829683960717399794697945565042391153811655379630323871905537955076118867541221110132913629594861913332194062752681454707418427395676194139780507130169687569595547741;
B3[250]<=640'd4549039250785210313871266097999632759466937585158811762504791368703670533560406443719507081517865401931764273535556512853266830178646638994163823807280283539685833309926894079390333906949523470;
B3[251]<=640'd4562440600625779511821207224748229432986678398698609907853605479637527187774069347010955578025961048117299597962095658184490543614925454001118236541334719672992064609834186187969984788629434561;
B3[252]<=640'd4562440617091057447432444226912365634834819298490208849914648861459945122055592140401029724085698818555661365309266443724409032091185152141811475429910442891094088746439791322991145620791724105;
B3[253]<=640'd4562440481567878762000320176274152468343398618077679597206990769956410128604669434820822458242638073123517337046290008027433847064017202025751522267886081743970334079626289604681069921524586792;
B3[254]<=640'd4562440617621935937234699320755145017174193775675113192570788157091368276009820802156882434826141742523196190501145762689739965935923260002096693957613524506847678651020329888996661783225363907;
B3[255]<=640'd4562440617622195218641171605700291323177029092216322109063056160847157231273400466370068694624582215909664224601178405836386940456954990146352217243304639562989759015490285360332005882785702021;
B3[256]<=640'd4562440617622195218641171605700291323606078945974082803350360789916167773334837147284924877515217035500127994344036784592373709499179599036711800378767996737055432831342937231214800559226425418;
B3[257]<=640'd4562440617622195218641171605700291324678703580369479901277292451908563358464529893320919746081472720861395405563339462827891254537378905821591106362734247036495106506235604884695247717293803667;
B3[258]<=640'd4562440617622195218641171605700291324889876555662537109340072192025477418508300845853079291495235266773900898482478059547282324203944206901465348999384351253449989932496588227215559224766212600;
B3[259]<=640'd4562440617622195218641171605700291324893019033423955321843101086915110668556386182125805674446179519534054953498172771830729087171083622847489270039598427615827938827116887035091014655077703784;
B3[260]<=640'd4562440617622195218625954989203410870160977670202448052567714168973082199435025599475759035890766305378281052495082259213042318199260854110323026248912645183376088030542400331741115520030123968;
B3[261]<=640'd4562440617622179009588361034185832443809835264951287993817756760819614377040621803316755454425781545326673762007126777935723411838268241702350139772530556366902701117736929228503906537699414537;
B3[262]<=640'd4562440617489346082120537243996544765284257991740927776025261237759314618629662889456876933961561022928676877637254895458746253597231136216300024770390679798174103631104043618598808673607927589;
B3[263]<=640'd4562440617223582379552871621096296803715247047304496939040793014238247614580269876425512144253233209223185950932276397849511550503592331835279351974817271451932817710885902360027225755292140193;
B3[264]<=640'd4562440617622162800674454923679348184204352418712456974203591673558613390552080188548555621254189468177473346165591058320872343491239848171748305370366794763153871483915764753544985040910593834;
B3[265]<=640'd4562440617622191166503539071092150515099047384105716667221500182543605534640724828288526960033213643434325095224321060025883750594164591238761365790888162196275951973582864432400020741321723367;
B3[266]<=640'd4562440617622195169175091311072186250721461735887840854224001733699961520758709616520155583703361483586194011107011812560794111289856386808806524724717107572558666159517822622227293401060081739;
B3[267]<=640'd4562440617095206741393285499954819002061914449340289483929470928478774757298011110494298987223630999742651270822382333670955972868603442654192220211290608054717946434050452633247050829566191218;
B3[268]<=640'd142576268238936304395112539389978693495861175980509239567013979823439580906677017122233821772224536945533889387053910735945992481498515689390862277414643637545013920227006032900417174132263448;
B3[269]<=640'd8911015769275822693770522905775148478216886624811285789529467659418616183787719715799099833853878382170667851037977268601727714958810002160482147600808240496800399590033381508655495061292417;
B3[270]<=640'd2227753158222841044029777672657396445020156567116245049267573831353995245950958779720120174682181157135020073217068565399662570855054229086843466453665310238679079491720439372647624943619776;
B3[271]<=640'd556938550108033894477984389357906259737484477193317972709329982816915703055767864692928940635225361758656354042254841705716108577181504188688348815116497535131395668120579918715986392305920;
B3[272]<=640'd1113877103781999608303659557254066562124969120269604461463287508175365954487409011344538281637257007262620137767606719597952714258429368092212742288835148075591091097182352210093749766333712;
B3[273]<=640'd1113877100669859774330854382968979213663069582339688295554357872749047063659595564265574558072362227763775513004068936092899853831557519191051803733301889604042922399008360470721642870419058;
B3[274]<=640'd556938543656803262700772864352695684160544476970988912521133256493957737058772182173719036074836182269249265413879091975023798308955228935494744353985360732900596064685453950447891014852936;
B3[275]<=640'd556938519667416356920307184849287654023907726893216359826087520047366710044512379828356248461835140635693968831932977124434087939011901018345409603632781492660261391638640652107356755794130;
B3[276]<=640'd1015855918767312231789045834301751977562517561031141768739524639281719425371295442045737210085799717968658393956568923962807203838089771547661993826413356797806378093323032400465118567093998052;
B3[277]<=640'd4562440617621935873918116543640384299401747809676645809133976361527478859531564745294170493756306895620081948680238721297069717772096859678144718911543319122681032323550187109773113544884567132;
B3[278]<=640'd4562440562412890574679560292692704698482329393027968205155693026685206922009476332648199660488463014105382552153882984366164561374524086721534678384793575664881741820543731622074215394755748920;
B3[279]<=640'd4562440073736890574271662547561967815165354121745208908344050325078671026671015083156234593770680697346008094092679023625022138676243676354760759831401583067832491309227439555758194800579731484;
B3[280]<=640'd4562440073736890574271662547561967815165354121745228721153615252111427683822775445325276022435033484788842097485869244610208550484250156467327828812054640554055189292107760297312064699332625179;
B3[281]<=640'd4277843929802154563114355797710650058975023709971845766001355432607689807404023145935697707682891855302662559238353449830867211052225533208018445088411977181615708528806601310116737716758708363;
B3[282]<=640'd68529548385190558141325428762225712172573422421614055424592437890080713922645154400464058949774588019545522858207539896826398336074372101887876723890783912668482504740275002664009293052189;
B3[283]<=640'd16452530465492177649008684286169268200161476414712726923739401300259681297144578400249092202330061283279687213466055484401840039801880389187938002690380922496205736343428616041435734168962;
B3[284]<=640'd135971326161092377264534580877431968596375838138306243052477374743283938219197503302020132708850962341217279669014769654781713445002007118151454150035465525165541832287614080922981685049;
B3[285]<=640'd186070713419675363980626894819329160794532062202678793890859104290773087790955271584137644454160207196629725442919723642926488070276553732;
B3[286]<=640'd47634102635436893179040485073748265163400239954371616014980064623351509791599631774925599910733247766437442948664956779509758648595788212229;
B3[287]<=640'd47634102635436893179040485073748265163400240130241156057087201006570605367641520027027196151121441605786972433270118711410317343577903047151;
B3[288]<=640'd21491167399972504539762406351632518071768467752802620406403102209373142470936949796908816987504445699718905015478269710773984727121002797445;
B3[289]<=640'd21119025973133153811801152561993859750179403376130713559538979227392655155422890060165807169536201562600453361118015612414114284408648305717;
B3[290]<=640'd585351670235566261830639000828755556460443851869789092824291233800603952216898953595708946952754531761060687833715099962832937826708063877431947;
B3[291]<=640'd1463390339831720835098436339685578050900757301605772889266134008190969295161712805781374657676425293827737979370721183017214207802022342520473190;
B3[292]<=640'd1524291284333980581729295522359944485228807686848130444755447734192076044345588681699368214386470687441288263584114588539519703095792366209045172;
B3[293]<=640'd1560874275157996115690798614896583152874299071332485575429578479812685869409882810060153051531745784687669239226012097563667191292985674217080538;
B3[294]<=640'd1560874275157996115690798614896583152874299071332485575429578479812685869409882810060103227033728931879144056968534709287570629575226050414171688;
B3[295]<=640'd390218568789499028922699653724145788218574767833121393857394619953171466573436083569631357959950740646080743624535946148416241657018563433632403;
B3[296]<=640'd1560874275157996115690798614896583152874299071332485575429578479812685863667683769218062766203938460334254552399593464022470877808794695363500400;
B3[297]<=640'd3121748550315992231381597229793166305748598142664971150859156959625371244102587482172693819740191767426503469139548054605231292972273573325716240;
B3[298]<=640'd1560874275157996115690798614896583152874299071332485575429578479812678010474138675806655065024462681120501914810646599636034123846765950345475472;
B3[299]<=640'd3902185687894990289226996537241457882185747678331213938573946199531660395982877033183953588778732968967348893102283602943840799823308209099694711;
B3[300]<=640'd4682622825473988347072395844689749458622897213997456726288735439437941816140411113991656362795891235281568997158620786064053083635395663455968034;
B3[301]<=640'd1560874275157996115690798599766097337893790554366516953224137169564862250398273976434149647450907332517351244827235618569373218618837741752066560;
B3[302]<=640'd3121748550315992231381597222227365459694039470169703591630016483123868084289261384452405272315819896127014411145776054217480204857626003081864966;
B3[303]<=640'd3121748550315992231381597069644145003872094257297377252888287501931387618075177585164194488703528350202011479675826907922897696274959461645874556;
B3[304]<=640'd331961245510479436680992629095292892082556572854552948115343382974648764311719681683876066210384222795253797230472162949674923035142381685579575376362026505916090338526388365861068053;
B3[305]<=640'd497941868265719155021488943642939338123054422144250424115169669464543921986518603893643586893102428553796072228600015722372308508213649360447087253902023757622975453185284460400873803;
B3[306]<=640'd500016626050159651500745147574784918697389989554003145478399338259669668661014863738078754480361065468486450476586378068647456307748824478793279219504788992340290012791408076111768640;
B3[307]<=640'd1032710687205257122549775507076137731458612774618125982515341803995573289408708024231859176239630099289657665791038330295745194823432014762123945585604708184701686500281926799379679408;
B3[308]<=640'd8771783255577084613319442293183890853466839185954005627876650883675521875677883229615766650800129286087413523976150288620509480963190255004330005622670876363811209166142442374074176715657249;
B3[309]<=640'd8771784317836861201662698293616114865186550247089207998240549777834827910335813689822732444562010807612507319196592891629529626245834811489786595025587084882749195287089737952276997647113225;
B3[310]<=640'd4562438714023382535207721371567438791044496720188106822537022874167631551357246871495199761437543972451253717245091113647843439696088092488229843646697739500729614887773478816335362570510402688;
B3[311]<=640'd4562438714022604501038556185387717714576758531440385035968580421979347966331678413116145698438039572088020135815366997712469386640886383752815423099256135230969180206529180563745149711876991105;
B3[312]<=640'd4562440617621806201553690594726127120951747822147946408363499873243408373790999535304609294052735220878426668048249761702917582676727461803552447522090320305976196781531076236314766029822150704;
B3[313]<=640'd4562440617622195162991831288993590462663401926858690048313052111888876116025113151681247988311315030598304563263667080287976929131578685442284999025235985976676720789753875403765836277802132048;
B3[314]<=640'd4562440617620104251811540153147250671799046200663876536159424031904597672685476141304554759995750855194373371406999603394631088206635266947371275789737729578987414591389656164681302625286131715;
B3[315]<=640'd4562440617622195155309187302671873738411130752449553743860297584490941121774522593194460234552548008411439675161469360223640784467183380664817546864108072295100055293946266418499362836104120846;
B3[316]<=640'd4562440617621182153316737769528782197567395809559373599319025505829288244487200690855490860729399888955111457266863115454083842256598817482001368806859932031269837051921344577707050934145802596;
B3[317]<=640'd67985663080546188632267065493026257189515505266221361083045030329248432277890248249598738121696796886443104898000674475221672998915167931962461803411545733703296462984379043223436003553;
B3[318]<=640'd141671244153765369734922020599882949669667467081556760704653730612052628422111094290449643781360003516464231451055987511335739446125600668227191953266266677561969269908968998851133461705541721;
B3[319]<=640'd2175541165898081169447034799806552842518514669476653689368778964945040376438204396468482953675640024221669340474231582843514846349637747352076800024487183369949849389598295732232611470604;
B3[320]<=640'd71288134650346800291268306339067051951456695425758748915299802684770910335451239642728520633783717721127741405146865968145820166573482133004623821755856365265293549614054339228243901398533642;
B3[321]<=640'd4562440617622195218641171605700291324893228507248559930579192345993774704543282465387795965541130495844456657245471026559377661623971354924628424182163340306875561905209953967360068772994244780;
B3[322]<=640'd4562440617622195218641171605700291324893228507248559930579192506808601676671613700784350679530020606661109372761754684733042464220590468769204610506145265152442354432791789542278336956705293896;
B3[323]<=640'd4562440617622195218641171605700291324893228507248559930579192506808597692219704158339289052195304103999829923243123162495860822389301803726519590671044761540037886597287125942546883469499716308;
B3[324]<=640'd4562440617622195218641171605700291324893228507248559930579190230446778096000738580126835486960580642255033205886688452188817326258098264382510634108962886118569954433157848153487374767305032867;
B3[325]<=640'd4562440617622195218641171605700291324893228507248559930579186845017080996026518145863622538580087862305069911795795216860482995839676080141484841286965581455213833629299321798407255680612974721;
B3[326]<=640'd4562440617622195218641171605700291324893228507248559930579186839471741607782366698310232426835385232084332280711499507984004843775722714727687047853851325905469213306848179009209656725977837670;
B3[327]<=640'd16847391196663989912584892709037330636965351848665641833495765970126417773180409190954477631328573814080769118750881141390542154684975855580453744137619647283043658975999999404380684705734880;
B3[328]<=640'd427729147826506033632727068472249122916451199915073670449502861603558905384020365059677499403915002239687559349181382815227728195298217415020079835272142874240031102636018426647528990851093632;
B3[329]<=640'd3421830734097022750562166195060621751218091376550053712523159985195846842417139087632099575627731259909315085405357185851504660890897602171598665798430161080581443726918380323380542998150925504;
B3[330]<=640'd4063388873846202339705024577399365476210425831802059799042330586090191768457854364431874885107038861299607514277662936555565871809745910211075411482703632670762732792712635564860457689210831497;
B3[331]<=640'd2561917338998912893251895712085651122645254942945910591403742180509968248892599381154830610682708589352416821927133970391415090747898679061500134266526260741269490470886094034431086765160021041;
B3[332]<=640'd35636996816213086650871986478402718273990729854432433500956879191668145752816956613379432260495807560066118124131580552384771425520335026473515532941344811617480313230329195020714186050635374;
B3[333]<=640'd9467955383249184413684071935657342837302842361233583840313265723178326062201520526879354503079183397384893031810029395876534868817471817636761533805742266716172001499238156136995031385911839;
B3[334]<=640'd17404329734405498785870883682929733465461600444348504728005834792419377068626494867385515327576550752757898735519957578680982471269024451913982437205122156592300588062511369291265905159215;
B3[335]<=640'd2281498778087075510926896904971185777559088242227042515128353910630110136230395937193220243678957842198676468478859867437377706748070685991905971706225952869621736943979443335578971015160796730;
B3[336]<=640'd4206033932957030854361448370265653068445607665095733292040146082948421949265014957285592037566577895349250062897095313435648064298993685378905107457833850168316936329912144291274510158957647918;
B3[337]<=640'd4205999959242325016054308837313425958441829157438128922069999060793716275213938206948826789029016933252296326235336204514547932459729916115478851371627720396170879729303808933175778276718025616;
B3[338]<=640'd4507861149422996553764584050664121410477574371353216121371281179674823462744578083369963869575042429173048115364029180091371467810488270702787731577945090145479965910324579681789403920947480602;
B3[339]<=640'd4531112875064056517690591843496552344543750916633750341097231517008377569320163219585269607015274638969081273708000203328643921461235509700833626148700038268453136645709292100581575598035963908;
B3[340]<=640'd2049534143140155248649100219074827876703355474988482433558478015251977689335711351327432122529937335320375294703553776701431898533298469139211932374151296316967279118656922540559023704576765992;
B3[341]<=640'd1995999232163117332529097673031703924089325949059973194403058049832371089492962660969027569031247163701526445408458255766635385631929295689481506490920545426307537942765335938497574666299140215;
B3[342]<=640'd1318796103033208876619426108573895428073141038199747132081590092870297809046651052131335961276754062486804119670634131338540615519505804263424974209589095122865170338251425964753990861789948998;
B3[343]<=640'd908895485745327506908841356830750235568593044145030621469291612570412596867349828183479251788460157815539628766058428634673241706269474739954086417379788201386173845239756552845305662097340495;
B3[344]<=640'd4385916591275850925865564541016360097538810855452855176500958724497441229459962415603322061416336249053173648724210107113630520870496298829716902410134893899746972114814868141561278369043249;
B3[345]<=640'd487321232961355080116091937864716175449411003887022697663182794575423067801463766538041235508178655607519115191345553095102574580423336087416456325442398570460972007665614587076901673110560;
B3[346]<=640'd72332394435263989748659931920205729470276861862659511838863846223409289564240532030353750372467527040938712695620635710668463422899508638558755463866395767487868066948995840615766779281014866;
B3[347]<=640'd4420971698803783685027945034991846663594756951003607079443959165011637492478643320959850071993566587183772680347043766464019790539977034792931215363101206922049155261357006881193272497551364;
B3[348]<=640'd8902314666419040124263608079207225847941918874579003923382785693920047667123270861027770138529773008212136730870400146540368831071623941009738789637156847473442242598512043284992958072503618;
B3[349]<=640'd17813331497712390160672146371590607341874005802798847537795271080957417508233162469848924831336710742082434553948857003578287104452948688760036038198743567440485011293415377977168455097385033;
B3[350]<=640'd231682086531189945990549530495379841019239176106895514129209770204217086708089929060151464401016080578039902983739531450508109944107570679894783998507923821761423875958486588456336564854981444;
B3[351]<=640'd249506297859547194808471234391793469128475401295117882188919858698556856222903633891449041303262954300098650698378522658778993351522287739128389335721478726954860133932967135645422017627685121;
B3[352]<=640'd142576136516195396390761940281082465787013540446670184550704031167575981406127221252924020459755011642482129456058741921905686567881005343076291502029028254616394974197876223129346177934560687;
B3[353]<=640'd285152504608555660891978909222622988447991755358254476266547927923097679004398409921841245795775089526858690177742916250631660279496133244580997093856149856472721520292635530921650731822749968;
B3[354]<=640'd213864395452832516548005611593480665401143910526503740317575144793691757223962894347610146907732469858949122577842530792894928898135973204271128217160557754343560291840514805266110976386138136;
B3[355]<=640'd213864400664624071305757099653926452677652580062625174638169874175727020370327431619624594528181344401943026958769257885480011047380248762060910616158572187770135311551953574187081748030955810;
B3[356]<=640'd285152538601225110717028584503806820808415622872228122198289359988434369835758106690309447676053251814227609642061623139328122421227966389498641964069740652623380949560795136446422817809901860;
B3[357]<=640'd499016942552418496316265970755617786721437516788162648356059593197097255636609044811814750349283622302367519818968201460682011046258428958526309255178042497260738112503773464046804407779590412;
B3[358]<=640'd499016942552427546883232504524845217725794483589452752379973045826945856296608715743562290312321574562672379441686602290081499979243022108277663991390134060474833751197639582919049485237250465;
B3[359]<=640'd499016942552427568649274039506574127040634781693080605378506404157133761904006139204694875727399664095098627026765659424274936418510621981555282248049139420417567316636090298380600246085625088;
B3[360]<=640'd284743468866615343847903920642670261326573744738977841749273263541288259411276733199018767759448188223365010617898880690234762131899950367248597422583494873072620655636389788877154577601806336;
B3[361]<=640'd352368382619953577310482357510571727022634681833784079240284201172154798157304974411723027705883809984674806864888075158661145818020870501657913226246812244609300393449892924912847160193853449;
B3[362]<=640'd385135993920240519938082537751448231673348805791308154502290934458454814392656576072242600284584699097881469433167499662488690900935906452091876507430920893501388554038316336664692989725386496;
B3[363]<=640'd395047699446784660943409256485956403779338117794043704709423197307692292696064284101447626294599525475801823814974808681319762575618184801599742537480167121947016981288606665311513914095636736;
B3[364]<=640'd303262767738876279065639154594586742727938610997555629254253220939145112256514115180531370154174882185721627887590435236484886283384502829714836538217530257132203401673361427602840787378897160;
B3[365]<=640'd392085801790617049502638630818246974506323264047085942860370769836614239355893537964619468674187917439051336252826056574437037591338744028465094302148814156412617277713026288125773559803937536;
B3[366]<=640'd463372907112131833174792940980257753905405451708719305268160624865340638311993866603299447682669736803108358989255873510635665611744349441255788455060481706233657188046160606409393231362129954;
B3[367]<=640'd67729171149444731311701394312615716782861045312686941080250627698425592855700168278032236151694838688799474986746657720384035212050000055126967264449639152604647876217013326357093947488;
B3[368]<=640'd12754145459748280680742018210370114897709372898794684238160733842758251260336992620494983008440222314373099089678923052975904106864923798493378599009816569204666372523087580617517701288;
B3[369]<=640'd6108553323164476429622526048476756783952740093468729929336056366563358491783133199181883561354584470798737412162138194713655619789765455494882584796090470021641121759252073485290184844;
B3[370]<=640'd1610042194534396671990187338440144458576105713030837653585897769312281903898107396018996747560974289823975506849436872886140388696622221234756976281765361720127382763781752030095212704;
B3[371]<=640'd618277867264230531691920944951357261466387764354788067271437311954307459723590618385431147216023355156652526371002268714505074742683270487815166426147009678682530107011444037132484840;
B3[372]<=640'd1019775870998044975103667148584328000629029536271407568451259008160786014409717671519619156316755806837573914604087826759059154661278778568559084795537507268590145988074466145989558280;
B3[373]<=640'd22425372411892710899490266346495789119940496085333141118416044118527127523528828363159067160666590028116766015503902375702507238841139499036617718419073194456624533869038240935313410;
B3[374]<=640'd1563984890472351173281385863329165827736101173877997527131234271224065813201003569683918680118854974622746960035825639212546457468361196396199980056331426265872348453554746950680588;
B3[375]<=640'd1427306152692637894257583805516168696462086946656095239729363768168923283406647602365631904127189303709492999492756263896980891848671259168558236889223539133261091621031855568650240;
B3[376]<=640'd781133188179467697535759258741321097389458275661959726495984332279762543626348143549449055812797725374757294212797203672546440871792652208596839448320640396919458429983449432457229;
B3[377]<=640'd162217078070493897760648252344417727409592792907072787337983888912515767944273352312278658127710527239634282741744661884160408557979529319180463048495846536577564547953331693158408;
B3[378]<=640'd15582251193207440163364476714523500128585370884770582960086804782365146063186722226679669293179249946656821816464632464771039027803016267669498982812266082004290241801295495168;
B3[379]<=640'd10130662308983248351678173541181553460343166580864511978132375121566477558548323915021314220797251305384358728369819707906105086489436299222701072166405530367457811870350095417344;
B3[380]<=640'd4812309549499177458274098083719505051876503741091594760413518596524708744221082500153566607322339585618331161191973279808652719108807330717194540185698207132531984607298294120448;
B3[381]<=640'd950738184014767939160278918317941411405762600321236572676110261629520176499721266627079729418023840411072409003492153416845737189516742532981945337542912360598560248440121458688;
B3[382]<=640'd221854889869907046852184169731981313402895676228781100733278593145327982742740300288184065335874526819131713193696019921670225061785095978320727556281265190505608815807169560576;
B3[383]<=640'd103940574804965825726862760685958533498776807006050496746372714078995787178453822123429914245642355574723773027969334019997383494058462033148117122553901236938054688016737239040;
B3[384]<=640'd25722602822445371729095889437860062626264668989815922152931128085769532788080807593864883483931516305739366864092810094906119477452159033003069768059171188920890855282977013760;
B3[385]<=640'd12861195972220804678516487283299324954776683091819118755754580931201009333809961614362260458758315300952813380395785398955939959399262017682215882423272277138200829479482294272;
B3[386]<=640'd6430590439970713834859130110918708757005551006363676254051579335679474862743770794403826182929899831980888818789701684844440007547178541075476680859347996072488194334250762240;
B3[387]<=640'd3153462618782940196753639265691054356410278465411135104842525893608119381784841800242549302812592987200856332081652271482857830483689082624352494723108855125912139874546221056;
B3[388]<=640'd912030855432073504849219921198461726246224312917128462928346345925919372477054175929189145469401920834445075893823356377060028758754659945035680872542026998460181692706455552;
B3[389]<=640'd230906130867494174019602148852043611901070434970084326542928272859489168245689329691201693165967469223737583456668006317483986768611716949785310097258106181122086304271564800;
B3[390]<=640'd522129892458594751667922073944609419627076987745742860435054921365434174469567054110829245730557058112148657440994565171944728241079388538754355173398908159545074158493221263299972572381184;
B3[391]<=640'd469916903212735260838053611675494176817843208407534738947261578991142684109158871424439733079578585355678416612734258442296839612173333637654616891760527054178245490956719899464784878239744;
B3[392]<=640'd469916903212735259449235439341084810392488029620406729289512744981399655726597586545009546688406948526504123335534365915769354200718173098759388139825840640242306585780846930191406055030784;
B3[393]<=640'd261064946229297365978258170400316061285564231661861807614007118081945609353437733474507680861676730773340024030683124715857210256911933514836322971517723830871272237173811039745511243382784;
B3[394]<=640'd69617318994479297306626556674015817802949660950392752482503445177198050333503983885700763487158676334877140055622722651583446417032847608808124005446385937949586692856699749441462209609728;
B3[395]<=640'd97651277742476921517697496371789438504278848906384281754753901845357073848940529505227365654425138566632116330263297504719601586240599205704124417091902990395494449020928;
B3[396]<=640'd26358768810862966234224777504822772405232992913550188473094896696458379728761251942929586956065619714565531998525502174886829901260106103842890927982428158930330341867520;
B3[397]<=640'd5203940374856298394037744472293026885694719858009697272697349712651382466473853977195980505118017669035430666523699544933759928371222194838985200870954613367301883297792;
B3[398]<=640'd815827956966554266653551955445810347888743754770198364985420690363350426471964608240757442039780528147858003580154244988819979259891507824774406428477217027753572322995095596769992507392;
B3[399]<=640'd1798530767977435871553302330262892569139134760073621986778798100615036338092890739743400323299096617457798562111799323436173233388993933853548659340415366403284839432192;
B3[400]<=640'd40886128564808777405664626495087188729279496453881422366049464754167142720421565036657550945942250894227016760394942372259357936144613226436856123104822485163719000064;
B3[401]<=640'd24128574462894072476934921449864025424360374366416215280933201061331737585307204757682461294962719191156713380268904137375910097875267986502064187832260927194629406720;
B3[402]<=640'd9213775451224466198364349927135264311946454213393745893719400076505004442243820456417124108494564227367310796925950300186846559794009689995924675686818436325121720320;
B3[403]<=640'd5999751436402806696119207171878923767078913122127159751620440611025479788431281092900362850295723154652249868900562681504975827671741773552414350194460331437606305792;
B3[404]<=640'd1151749171121290586621121574540988240306468986620041234720332535540872954373240944135193640640155851251929640207405414426024948739157259780258362293183032628604829696;
B3[405]<=640'd358116174878780132775412290718817482215185735436987043843100595854510593270604114021149898288119365167048876356114142499541524659700335792056805954575240098710814720;
B3[406]<=640'd21988441170829878714229983704359833568308823877556423808131458628914232861005178377813029587574871178817492489171372808154457400390009013157614784642420934363316224;
B3[407]<=640'd49488051739975160210937263838557729716053182532221479651376769832453765643552732077713268961532303546168182869013034180998377062506110337444819254235630412257820672;
B3[408]<=640'd12259540090130210143158765206350490722051834292441313174314208520065808888459973096495405839105336859310375123515320666873810081276867432503378617472971390383554560;
B3[409]<=640'd2706377832683905618302940452991104074178504247528477117422346215730613425650897336061844815415129536484688677680108873242776954627322285428674671472001985846181888;
B3[410]<=640'd731073494860473674286669170532835289962991809634462777329253303143372306336634032494795397998371052139526014947631233138524986188069494177400497085688363903614976;
B3[411]<=640'd365536745806634706283835914426238774209402367236469387008499328136950077668823625820181368526903774239488678590224375191680736866666972368297312504337625226674176;
B3[412]<=640'd35171790811679178874709909017623742201412528427819272767277154248008583448792395248077216893961754470503597453136506452327153957071420004691921542508408685461504;
B3[413]<=640'd9665635105463898478694516328523050588641941934235139398221612957163190018488989830864030181855238290139845784156052926719528842988210456989952536253589304115200;
B3[414]<=640'd2196735251260626861814705084979595155584095695602808058421885550871335804933437133981535060674254851965978085232156785190358328272626852337333250871127353327616;
B3[415]<=640'd1098434299498481621167977776419803952304586297060224133326003840697691253451542032771423776906878885307123964450383015074343369828980596632266091919114151919616;
B3[416]<=640'd191797016666424521678277847876448083506904186154354340332623540767736794593384007190008383952890067791882992983000750709030248562869016181453800531636967702528;
B3[417]<=640'd75405511797997166088004316606640465769356055674970975219043922004410295009141404370326460826191183916745855238706684724160260428518046717173311260385884504064;
B3[418]<=640'd17604451812014629991740694822817567821263365205417752638901504983589851079461518816744741295907694417872732514607929984399716572745884270611501715301488132096;
B3[419]<=640'd11798870978449286514102805091649837535594317908726140534049805727551940596131114922960659540539869577878625186165832846581517262572183366856166436579955441664;
B3[420]<=640'd1072833878844855400481831328085164388339278623236610309376233889198148424445700403447693402296169811574096247305127254771846570118853538795213159666785714176;
B3[421]<=640'd588316673785349889871860544944994660624913218008801604037573794292759985996769098683100388264612323202384273920589253683691629487026060424664610066818662400;
B3[422]<=640'd294552780460926430031266861782226721543328086663742338755205386735604778431135171974467061656304814391847953101870589413311765334473497910404504011520606208;
B3[423]<=640'd194609618420641426456569282923385297198980018845278395255245904068353909278160193792845770370513881997216431778338305673390569992630962237712587842327150592;
B3[424]<=640'd9268605506279265782923022371634591067579281418125253927860838517478083772435381750268280896236108398023309501468393044901877502555003407117156833858420736;
B3[425]<=640'd5237424972633826992021103840861772822337627949077463116748488285666831878353108343226988260166744588636177888673573693994376327721266696970593025273102336;
B3[426]<=640'd523742497263382699202110351574390556304285621707341846147460860652376552395721644850065356514817482916515894778837179666740712911074600540540682991828992;
B3[427]<=640'd209586505679787739810102313753050014764294857297753749967548210938687423262969041197998943120185447676926776693061404152382724431324688500030618252345344;
B3[428]<=640'd172261181780998364791930066870371333827248067915675813307223704802123244682923920354202893058654838852630106272849657134418266860377929032283646882480128;
B3[429]<=640'd15085089528520746119293714764124550070108670262484445806811696936728815402465463643453147868052572578275332195213908917081436064410569078044944987324416;
B3[430]<=640'd4500912774836855590227358776265690131379387743482983321377097753561286670105408289204790876403097568508705083153322864812610051808327451923621334745088;
B3[431]<=640'd2659629868915615269391264421241929170908922968654892536384151298011797825637468012326357225794933077562543794926611429015793410091206758634637334937600;
B3[432]<=640'd262576514064178738565969075271933372844643269726837580155528501532967944805807567245062515415906870962009154355613683192907297034556351304827593031680;
B3[433]<=640'd118251835085969785724735067014159366808514763281408640676408459211273747643649747569922672946137790154208326574918824411907600470731381382488317231104;
B3[434]<=640'd93496369081963967334037843905288453799775423070040362701536392526888322315382582451242727562022561549504810156458448003833836796058111180401440456704;
B3[435]<=640'd9989607554736719996424817805410323141743523787901049805571802513056212754741674616189980264048809379896372133143538364831386636540909703953272274944;
B3[436]<=640'd2572329951208106316294193794064862922878795840858765286930794664898756731369744491185302769678067181125637022128329174424383906937525564036154916864;
B3[437]<=640'd1423517340432658186896799967043970434217317740757462670731684500576423010347888484510329018491002029376483038125368400598414276829929643827045335040;
B3[438]<=640'd168574445301527909344339414129652555247413856953220926704299251469004776835350212292771491253653097421496334933700233148154823741759189519804923904;
B3[439]<=640'd15608784432136751820392219323928653934090316427872374174238456860503766785850843151372994531459139333294512987882861604989308696691834472129101824;
B3[440]<=640'd3902185919208575082537109740147551446973702898262765808235316529774990717369592055174149766495574837461175011988110799466707712102856881625628672;
B3[441]<=640'd1073148334127556894331550923015246924518928987540355513130720440148893828067361213547453700213008380609300858973090724410821327236840447105040384;
B3[442]<=640'd283494199022928427539115963867879844915261190195955733381361633661966051364098779871133690938222374793708434021543925470382356483580338223710208;
B3[443]<=640'd48848772252640533955106017443128857045672840110804777878161170087241878059538271804532008767120112818465404015479034324490173953175844689018880;
B3[444]<=640'd24293392344072815521310647387611616683963038143893598840291934773133928233472688681532553082669717562451276110506668196817208388590092557484032;
B3[445]<=640'd1577927047801169199988244775967835815268036712547777413131461121498502387231767973800020534194306428375662592;
B3[446]<=640'd536455151450859487650010068616182585360384;
B3[447]<=640'd34587330106315926162967454264754398477561102336;
B3[448]<=640'd1332688833082064660007289256600604206296410956804547494467003505198765369790173679473367176533971178849528435396710806400794624;
B3[449]<=640'd1343265728582708651681775398172127910270556783143567061145936857424783512390218950899794811794185230378497549961832982512664576;
B3[450]<=640'd1004805072561177875103996433757478436318171279730937236005812105558719896897916694095241547411949842972419467860087175452295168;
B3[451]<=640'd994228177060533892823680623281287643901937641531115018303556844707608885819493513125151855017802615691083719322485747976503296;
B3[452]<=640'd41591230024108295019165534594378250277249928634716267605075259570741865420545224577427674353645313780920972079919898231852406669312;
B3[453]<=640'd707031448922119830407060943717761769933836238508183212835607156060342408438157572123089780758047141280127601407188598088962353922048;
B3[454]<=640'd1039751135295305572341905319053656388788663903280472645698821633197616497450625125697460130571413719811643687180570598626564126015488;
B3[455]<=640'd1061932492848272091218532632526801058417719843506532744563599693144476284299586867807880580892769614860015570458459303110331208826880;
B3[456]<=640'd1350290141036836836614687707677681763575158305570037637646909482684991191974807806199015653907410501345811775449950450540899999940608;
B3[457]<=640'd1397425525837536252928986851862176192671766694781804190841294788580473057930987331825648597045980415225531386604980372704693692923904;
B3[458]<=640'd214524926879081553593185730852746716030810799992437180566268454546618893467791496111519474070433713874903195561513164536660229995267370054420146195133366272;
B3[459]<=640'd750837244076785437576145399899527383138846679224219671557558532742592209285109125087561195688962264199258133224477516497273940582566751506197263134933123072;
B3[460]<=640'd20839919903003640765951255182800189849127726304814424606001737109136104744374781871363986930235800774173521902119375463386825705060944576512;
B3[461]<=640'd2574299122548978689077679014315337359771576566618258138199121790300168402567907840712604186310925973246885913205374279388629280764278171759201684950341386240;
B3[462]<=640'd5148598245097957379829994449407752995207404569230065068549098627787715941650076980282608254262491343286852471828195620507148502363831892931696699141129241344;
B3[463]<=640'd3432398830065305238377700769616166677946315049521052058426701928062901670696542049209819783784728133299938820537013989771584342973270584426082489897869902176;
B3[464]<=640'd1886981224712488083074829900122401357068973050260218531972681059087837608883430133944256721076911795451753352872233009344015394436786400652013293199128199663581260677120;
B3[465]<=640'd208851956983437891480625692368658745414084534001922274772651464830483484342815586612432582031133428915501422029513166291229588071102861773436313741011296593151187581891326112970943047401472;
B3[466]<=640'd487321232961355083977547625976775336389441157616330060076779336262521171744836601087289018933074022455316574504544988781851396683540227535218326698918728102373981930400087612395411524812800;
B3[467]<=640'd526073061014528585640278901035463626532846305439265735169892540851535671826104537847139391879072700318370512951106478674791030177116176195429134715002200911744216050001468720066999447715840;
B3[468]<=640'd7614394317558123141589522214861809027079458185377908358033312855485658891423646744678036558856125793400859248848003122208289418253371217373951397539037871890170989179017066623832395087872;
B3[469]<=640'd28365890909881818463269262002501916169296759746711675790473412893263049071369277238662506927571058900233729130886567925734196825640887888322512510781914734964054525495808094109696;
B3[470]<=640'd3096695337307324813493593548902069209092764232187876607774897671977916778416285279296485549253797423121494282866085953870988722289844297909408487110951879069124453038091636517634048;
B3[471]<=640'd552483043547986528433867436821658866027953674442417976002533195964595235920932391206358208427135573043798334784175000924724258830261981978069602945569788728209268920366578573911737714783816192;
B3[472]<=640'd2437720042765361656424273317174365866515598671657093428852250411743105066961485425629884726586941778058477703382292741952604499724144585868302310216126716077141867559759829425140967100313247232;
B3[473]<=640'd4535690166179384358454411303477310050613255391324264702904056018628223274229160165776991281891747765779718023625825993026281343215849329260851064325058766332796821514516211134753614673081204736;
B3[474]<=640'd57849818123121771312898029941269012675476142848185188303434589869056144009648094948560245217020552387841173117082260543817305049369394760027883178908507670607825662196231080851943276461162496;
B3[475]<=640'd17822033048458395878430144077209414171392579920544243368989280676203959882667666742788358816893352906455043225217364679119215729975648933590885952432824102963280783087251469511320863646941184;
B3[476]<=640'd487321100630710144653069192900886609932691024529593742558874677013819593893833719583406443357217536384218302433574985859996177567360346455783252664155269391311623950957619980104335211102208;
B3[477]<=640'd570236543674160910926554441281350519961256647494432469576784163060499737549190741153190317947355987479086345580570225812670935423120640267183148705892012306894478883823649409915703950292549647;
B3[478]<=640'd4045605907713977620474468314488551879232223853201937860941234987322833916082599182783946149542302742573115421864696731733038121236433943958711984421234940700685188851129908450032494572108840980;
B3[479]<=640'd570583529595945747241513421547470043938985467009843568601896067172630987535155702583225435455069157787082995536952728357379495247087065396418412562525614595478326027677913266401561665762232861;
B4[0]<=640'd232421501095277224926907736380909710267726162562408446462992241857670737644375733769835649194152713847361165724997507307731903689599469437819446673138737620934798431808413088333428731;
B4[1]<=640'd235485008534003883635974162671035322861863660690492090291286093423862263398282992939417021374139486062839742804833472222762438125060033361464663708423299832126264748566670972775563263;
B4[2]<=640'd269199822531343101620110199564938816936719399294706799804741321010315447009104265205645812250874440018688447675469958272674184461997085974206633403082672999942706515880321264027435007;
B4[3]<=640'd796820452565104654056986474597816319526844740541887636112755313283598591371126549726876395714118515665542871898365085336384365579461296067048938635703924377012910520244849404389883903;
B4[4]<=640'd796828557079729508705434528713879553965719959559673566760792195597735082730075781794565839359438964187458898068373657911395278516064301245136705626756751825124419477632027503020212217;
B4[5]<=640'd3112136676668255816750331177856597414323539787758170861196869526617226134744069139591068184500963861790360378269603385398414173788740950075405176830049487690235377953264136997568505;
B4[6]<=640'd3759270815843378309122334489283900819100976283842806303118313561953859939270708794715557393043746236564381418437808090868871872456941928476955388232174972554960699391999;
B4[7]<=640'd2281220309010274419944184609377479914356431642243224004690778912210290467986766846652521385675828121378874618315254777087256949428336232845914411801672248715179651661803976521330985975771299711;
B4[8]<=640'd213864403951137655144957746691396617807510941240578235352332462232133168116694873753013579515460802755685829601900379046531169410757940959723372312163953381396396393112881651347641493077622767;
B4[9]<=640'd7503744700755774484386338076527174859102907339979663787699714348159426185816804228207861148307530230651654493472107092739481551519920937241841962974979608895196114190335;
B4[10]<=640'd2281220308811097609320589517873426032917288809638615643461433797148124130263474269222600342516537102900807071488871378731516663521859297530202806673537994914625595977814872887038217257297641471;
B4[11]<=640'd2281220308943882107526713561309131279245597120506539537159763513610097821091782461207933213223721731739372322340006251979121558788118643338631384221974505571440198652473495282595493939796508671;
B4[12]<=640'd2361419460292802595830960509772930569895508753771994505945312384195526333922168273525799708593847532845122570868220082472951879874433667237941420563749280229768498232094633423919523150866415615;
B4[13]<=640'd3644605884001054922675534486077108799079430381062417738923665833065810800076568315568822952292126363575829921964091602588163771612313534532800149291198522010095811176432052733488610986810146815;
B4[14]<=640'd4491152482971848418349905127374273809608759860374489017836184544193042454246104124746825352963875065546989926618816866650215908320439734182178735734030549327847441489760155102993797167225765887;
B4[15]<=640'd4526796550297021818495538160150062140878724315205969468125452381292475569355365334664293763835428384800549652241408887709045170600777172143013368557751990705496886981015278631288987165080420351;
B4[16]<=640'd4437686381984088318131512453005721128653426320036673125507786390019296164674151629219132682979605347376653343782329427240001792574058278434164955403955407110629184917962085010432979494974259199;
B4[17]<=640'd4295110112683394717548915456928789882126660714473005409784092065489401720761436253171570194958512250378641904635233987697243262568784561745049546435955064156858677463309692587045256410643300351;
B4[18]<=640'd4402042314658914917985817916437390458756430795052866048348088856545907111383983840252988356354595189681955181871196935310733408636939966099764774288861285881436250333601967704830729501303373823;
B4[19]<=640'd1817847433583843407427341811646209825085504504616813430610548950298855663958995735034132343226265167478735143495050771134862913968482970697468153486670060139180566867456007831641400093223944191;
B4[20]<=640'd4540197935192706393608371455022505322779530597960489336843192162037872462773965948979093677185562656579106564652879481038103304107185466271082433606429221638432023096951739063493810962793758719;
B4[21]<=640'd4540163109536793383823244576102978090516574976420913630002611591165961302257261291523629748346972173097547713340480203098773250906965167814042692264115078984222793206627606471159469050928562175;
B4[22]<=640'd4561535728446593148870476128064552015571270298151565872665346431205897655843745525570835867790232587625153938768046265580725759033900092471371581198986719141171280711239842238778453916781641727;
B4[23]<=640'd4561822903074273332871865191199320530357210740774609079815913646494623458983951142656024972419001910565620256866556575710581165190825382742011590807469988943092866757389994881251469327383658495;
B4[24]<=640'd4562427275435815859575622324042085453133253387114520129855697199340261086230114275471513039346160869083586956588943623028676561055780884826146730323765959932979293616102472951727019581272686591;
B4[25]<=640'd4562431065636532425657467767402416664911282553493641791849983412640522205899711101954656458081421470724599332576284706232335555213002689509156341148567191068334983824274109194620609381659574271;
B4[26]<=640'd4561883399558870720041255322017500579221654576262543001960559506713810458122113194190365894832689320653451832938284126291761854811203740204772609234008074386760943565911638894956661695844450303;
B4[27]<=640'd4562440614402171137428880863817190623468601915610089614215307944085350273672337522160695628323464477272545433821778730289585827643976788190245611474170582775338912547439791887285975661477363711;
B4[28]<=640'd4562440617618045895000625542187550358189247857802940628975386774572630585904294183914763721149025275215331952674211710278728231108344616251174489190153849745354077094515154933136961716854194175;
B4[29]<=640'd4562440617618058053763218569917902382020029854806395874039185669042904247852013627385781663927318314571039722317013349615691879683874807288076478160747211942997646885364990385556339959558832127;
B4[30]<=640'd4562440617605609554544012677650100105159919735177272839887669214500434357803813662820312080078181230218255070840964830973634828193063772729207380339339493911121180442629908086891269554312314879;
B4[31]<=640'd4562440345663206204910931479983800390220507716373711685254176670460099419198484392091889391499339956614239577437094907706430067622573113904616495362230632966792737227303749624081444353956315135;
B4[32]<=640'd4130238896973058643678416195758302290603691884889660543428529446849649822672778479999975953449610339484391200914735112306058312912520738470298318172554873206607264067302814673207203646391975935;
B4[33]<=640'd4562440617621965142008505264938526833271699975419327624189648205206791855851882594189987936529114412600545985627314873828950887656964505167048818916382069126549846773485577863339780254250041343;
B4[34]<=640'd1140610154353460978579902653323108084580615236401075261020668868293992036700586275234664920834510616435820543828866833498814444502527961302176608017164431613941389979024946093754322234531381247;
B4[35]<=640'd4553529600738619524088856500675903997474710479709457737815779128804257845370735912782030152027317221873616014212422433550129048247958438260516788530656078978649075637695132444801940463116353535;
B4[36]<=640'd4553529600790496579158405340588629672341447205510293673557492256787043093270197884188413818020106553626824335068457647969168448883704880550139141469903344742617425602714165861821029393329291263;
B4[37]<=640'd4134711809720098207848265147968218915581263338872152601466652075468542392783152196140991904554884058068789843955528142732647954532411358511212020274466949562129688619840001449009264408655822847;
B4[38]<=640'd71288134650346800291152831933923016977798410605138834295982688248075968199014592239586765400193086554073733597718331886830266095031006644633785277819724164814581306702175722941592013140656127;
B4[39]<=640'd445550841564148559107866432751306209150488966955906493146710481396888356193959441206815810754366157076759683030324474090550923939718177890965695098062799890326207764346524342558952974245117567;
B4[40]<=640'd1069320931984592715629523790952906552545993756578689304632543423053891813811453332270160602831875581666095524271680677668038949798736898563724326656350191690054523977727494926184280350681752575;
B4[41]<=640'd1069322019755202004244878578719449173697036193576887362174802559455792407551161023560394434542917233504584642930009257422728921106138566654536914617814615245036996810106821194864010065090410495;
B4[42]<=640'd1069322019755201917184091950420014821882552247077278191489085970130011021358185325201907816374822713770831765113529965302240671897973214160066434187391198680539697997607290092510914802190614527;
B4[43]<=640'd1069322019755201941044712751919529492907278682164643822139738424682065535368192582578718212135428926736993848803319171965587964106979222565187607743299194602290702367329172424915508822018097151;
B4[44]<=640'd1069322019752089867688499313578416710392962917802096573258642305655640757242112651628492559380452037323546847376063180871073907479173563765553946431399896073952347076130004945186292133049401343;
B4[45]<=640'd1069322019489633001557113692018356962543263187101892045888113585943376741241669666698680464925797414506595001185956335684106007684394347896204852326323748646991940641995833229782773243859435519;
B4[46]<=640'd1069322019261393404549724262029580649429436759238691314558982320916341051616024004096146962329564306442346496123906147825544081442139365628316824817201346477158287996469635388109451974876069887;
B4[47]<=640'd4562440617606634434037901081094203584528796796912894749836228706425605664148917591643999742503995943050230941500249010748627955193356224603196409433596749010448858766423687139669826696636530687;
B4[48]<=640'd4562440617621238793208096205826759949762702711770423252806277497293377838573957887565455058342457656046451910049306494316648188645563413041451139610049485962169311710484464241132096694049898495;
B4[49]<=640'd4553529600789868512106822691272881919815143729842285467832503877317791767869269113818385424815931368931030238949920077053438158489906700145119295471347521813004410659092310599302936576827326463;
B4[50]<=640'd2272239674660566582753894284570342119444893314004490522452976274696199261947475880000747377681603523497331464750330814176308275043179587403253528200797352781434478884263373198232967986016157695;
B4[51]<=640'd1112206288255573895653345867592020210623164220973611591419178034349052559582282572498255711765034779540545038069098433246856424156086234719361175141660801681965897893989331591729613243903115263;
B4[52]<=640'd1121117305083755107281780850839391023435290434115033478683421054478380686587474568284518556560941981517237560672001327140154200068008784042121970902869159719636718175308307890699896679087210495;
B4[53]<=640'd1138939338745843414814613074872380683976925384873850316193930166900290976160402780834051571235998076213118817508701038374243767778433211400272505317402619956066527304004518573593719142506037247;
B4[54]<=640'd4553529600790117344921589832685408998362600250315769860267920393695088022581801227458749451155116572971074174606311286911678622646275306473336135525848944808054480786097787191179697361738792959;
B4[55]<=640'd4268307444869735576190995379055973361068752823155782098261795931095548703398531507010114949374459310162666841293351833420633040563451714540607544468609279429947742017090640691314627851197612031;
B4[56]<=640'd3483711557634742818438480154663536076550914634703274344557586355720873679975383588523711568875356679086264404491698357913897332089323671130508918162770287288362652887156299360709397397364539391;
B4[57]<=640'd1085194768485934039931230789122935628268818665600901196092824664997005093321452339992371169206759294284926757043350671468310943012712953942596740279170793022013905545805173280232002889298477055;
B4[58]<=640'd1085473237761914616632736652451698659049701207970998138624314777216167631751677137327565094454204880444743913887748661797102661414568175575433316660334840482664451278750726836042887669296922619;
B4[59]<=640'd1083767613446549873976116298032360148915895068392705882233900908597580664307633767853898701518280397962941575742049559668148324799669582773905560253354090156307730124864588311410900741214175231;
B4[60]<=640'd2192945548319513082777341547432105728521516312855819351304121729908971731766808307308831522852030920596492321858835142456215925818390348393062641619104363743900382419654747169990236258172927;
B4[61]<=640'd2303254190272850116944987996405993602772607829920674760764209561346749769636535473413875834826403274585675704983818649076554096472409883970282097858041671581195245467502898364727428942458257406;
B4[62]<=640'd4246656458662097691024507530119408956186702259302233466445905076906084784730925288032872509819487768439353262195289831234984767928562100927866166647824026387482949243923577484315663628500991;
B4[63]<=640'd516838976215012766931915928543965139418932102695583699341023617471015192050627394287100229690446283008115274063611480823645037111968520465067535556799656661440628574732797437109785822075289599;
B4[64]<=640'd3992065923100418216662177862909953532115791741838841416920907654726717326737536195340410066223867380661397009078166106017072416057059943715028348446928111133082205186646088887740803671490822143;
B4[65]<=640'd4562440617622195203043952885718485373599051311006101000833609610256794874955447183266131177003912972541160757154414963917424529945720300148690904171084376391902952708606113647862042258640470015;
B4[66]<=640'd4562440617622195211715935461166855117957072111507959876298252889235964633905963659477613280492110996522306673512642250254219763063938983814133791831154728600423683599777481493329357059248881659;
B4[67]<=640'd4562440617622195148893998397713419181457217057729215258870726640889721022962530579380034752499667020188829804488408995707331597000679901766774350480043061384822991602636517271457442157247332351;
B4[68]<=640'd4562440617622195184633241410519438252795045363505352946318163908515410383907254951542678937244165429482457253210597051864224799332319070056678336457393544497933476166475522347284064923564376015;
B4[69]<=640'd4544618583959604938708126453535735455185904743800654805707858827986187417641723190533956552774980555624580614834855206147092117291240969160903012803323912906730286948619481074533749481829040094;
B4[70]<=640'd4562440617622192145313602917085044227232595459973244805099426280686076581737812465332488634829998713894044612853977574762015319104944415129720630104928455375058440386772035456637449215194169343;
B4[71]<=640'd4562371000303188484122623361629606808031981852122224277943355635293782302090052645348790746941020798157844888289123080291177588181922336546747519403611046078453493989223908996603643137947074427;
B4[72]<=640'd4526761741637524518498824354549917835304698594446618634081416123859053039846023642688893540778898023127081558684582210460735945515312399477831774446864347839380703886289053380197421989977128959;
B4[73]<=640'd4562440617622195013051641760423705152077365190156958737687830357194495714642511901669405339580807330040456071083668536580450692354027406588079661968927090353687524364348560079030098815635947519;
B4[74]<=640'd4562440583629355368066589665435887268324306228018934817823763015011830747160854299958150650629415774674732308352589813017445710340263011232049375594322671140778626939922852681856533703386202108;
B4[75]<=640'd4562440617622194719157429250890339239377562682769918230178890811885829201515607197964779845640462346216356900852851568343184010421075931155216226960924079602684280052933631295296417105562304255;
B4[76]<=640'd4562440617572396985489231826073418929339864729786714658098173181260726802122399566311031844756629006890554702929142320344470994086843009813586411255989076660534337003643609393227389385859661567;
B4[77]<=640'd4562405808946095975286842743755213646171234214821911136216579168420930464345025434103637622397393539471267505911863161319238582225900603956122734642555928939787105396389887482512325524821377023;
B4[78]<=640'd4562440617622193240052185056430371597220893199044856655385624309143925544368180883100114599632803321840484332510844769806420995266595496254779395455800255854928353902528706925585009817973424127;
B4[79]<=640'd4562440617622194712108874549086800020542477847162306821831605715804081475965717015923392018347784946715890085067364362352699950463802821360134998245946343513158851387070745915048136139503042559;
B4[80]<=640'd4562405808962555928242399679305760767075908438793945469950858149686334452710642678441768605927522094265589987966602230746988880975715876438741764270204588666760286348056324306081215469066386663;
B4[81]<=640'd4562440617622194207554854571022726418609692866748734067718410392569166479776043354166628696450591663341321638609398326829861840427193086882501156486485948041452381540881249526693418341769203439;
B4[82]<=640'd4562440617622191172316169580065214625091690102585437556738566497118399352823838996383655652229959998444941973248175393834117709884726098479621272092280955239274172125000781712276057038604109683;
B4[83]<=640'd4562440617622191166383259114614664858216828992844659781921830404424705766851913532613427858010475549158007896881785906168586828832378386382600622280453455169833203930098633760537481752508039803;
B4[84]<=640'd4562440617605467262397533358460970074073293317210638374786183978166880463165264480501739491606407912584633337685322422852809572212780732129898351982207502938742927845841058454090405175766223096;
B4[85]<=640'd4562440617622053136230869433479260783696829359841186293261033667363182083778707764720134982201619853623210150594307138334259634996427964386656069104715572048634446680367453955943412149736381691;
B4[86]<=640'd4562440617622182808787798114776483713966592921619185982844426442168940752416901865180277898671732395880118166496180899055090758331452854466385828347301567746699153664913990448006180925842883363;
B4[87]<=640'd4562440617605564769935342223857982077438054063261102937227752102844249877919239297394125005491508134339026058991335971538516811908692188185188158439295559299495713274764797995437585180626224931;
B4[88]<=640'd4553529600723678874533297625333370395146621374942192682296885700902152805137145315656269076540199411964230957493989714814811976861258896546053323651708911540008513233583826240013858861723091008;
B4[89]<=640'd4562440617621623058344548081901403212284796418503864074776281400157353341153785237587174255731678760031449677542098535479173199859154972920265158003921846412856280190389591439178830546164711648;
B4[90]<=640'd4562440600625756274635697871936080879882792348474779600316763000962497848587846130583978290465536058345837272990490922485955133558894772233211391237984116170176647611078097528833340963347702112;
B4[91]<=640'd4562440345675369193953768134836601870085223218374967274840849059054857817018906232772765621141305962728776881717332100534314780089063731995240657015572583561560042593025621215597685693625610737;
B4[92]<=640'd4562383917574529897937056049603667648456855207647377668343331388388986766591185494473680447522536435358661241334003674105361622486043163440976600239705347576022741750468066663816648469631688931;
B4[93]<=640'd4562384053516809479726069172675182727489519618224626885312416890519872943021747034447519265772965164599054256134434764900547363889073581878771749898831728505602865276561083959112395216358678627;
B4[94]<=640'd4562433819055396318044448151605744191948111095779349552687854715117466130706697700047526770402813946337106490762343726821266003295666914731119084741907713429880967375003494807228545926837501955;
B4[95]<=640'd3421825840187208346145525173722527082211071536433687172696915079338254895708090561345051711147917957219758736757035712932285799873094492270500712108772983039211020357308173941930287554203942913;
B4[96]<=640'd4532365651022100024784520324835867262176726303385582506653073752651892491804669285194609798667526860827984821092392078406524200786992321932594189951569078179875978793784982837714051350388474624;
B4[97]<=640'd4558542047725048908478813222562219688450481616170482625323639905654962191464389049392674434869617362903156101780365248361307111260719825740746482578849550352615005996292690616280499463609319424;
B4[98]<=640'd4562440617622192176353572030256356547312601723844087179569592980247950460977989196365351852823945815907375662843413553408908628494818118994738441123560756269191248795375580140067789306068926464;
B4[99]<=640'd4134711809296862812587084488937193758022480420122497831484683480530449605893906929112482446644958860480831638993660869513750978349494043488657203118649370987624969839068325619442205908338083840;
B4[100]<=640'd4134711809321663666773195864249649284640997833819068296598662511583763250364768896302832710332102575672639487505268062256158725848123618949125237104997696808051924866254815340927749951604130048;
B4[101]<=640'd2281220308545431326488111490087007552094397446207582770217600750738545152251974128077527291639191517172674061176913725312881150035895595401614504895209111741312193922507093642466476607063228688;
B4[102]<=640'd4562440617555705618809080984537553164859706788340065966643269993043224921157673166785534210060742249569526835052511466560017984141377720480829318457688544074880442103371813398605403169304510720;
B4[103]<=640'd4553250995307003408727626127790379927415972417360797075637327670127970811252510911808725534770975426316110063040607255808726353782654826419561290816225921527900447749147668268062869348403841280;
B4[104]<=640'd4559098986310453718595649408971772082804594684779914794261729197021371014482635554309407231087469770224923576929715532193823951016775594096670128140591631548014958530347704525153017196889768128;
B4[105]<=640'd4562440613904221742288742203630181401654580827659685061102365914118205213603683482028319541061759675119539616895533175824106895315199607147676701092126370517850063298843512880251204469658812608;
B4[106]<=640'd4562440617091055587507885414657562036788678463271440145585286527194224469327062763182050671203702298306208642966185097588570454478013300341331792353484792006840852272292666497846705195753472128;
B4[107]<=640'd4562423213060072080728812785503278936225951793496008068192486705143565360932774709601097405348523638079347754392087479893120882821110390595852124309055198090499737190536680927172736162859582080;
B4[108]<=640'd4562440208546343131856657436225374265262272259078298424279936886586052859853722727140652702373283271116552443747144698038769939966461078983077580063781768248591586107547821010976208438492136320;
B4[109]<=640'd4553529140294246647222235183685291067680996579473288181705408190689832779265327745403929634630909306079555087019694343926650992009708831992617711023914709030150881314032760219828291894704669568;
B4[110]<=640'd4562440616688546142778920491689678946580062772856382866881309033983800715452189275348015739162436534155568789095750591840253709975028171339927495754517840711223631348737063376057669378476409792;
B4[111]<=640'd4562440613389681241774571994107247455711900936447890828837192320570161812701220977017896428153384484411781838804056507652802424381928034543159683467511509018007998522473881983760044945344824064;
B4[112]<=640'd4562161996017496723500027504303595456996557016594252509948145477668463813512916842933065353460967269745310640594910749715429285877349527075232763156364439421181434729718366472351408252551430144;
B4[113]<=640'd4562440613447778508545271373561515616600759199023162718963641129489748068828074514758774844914291156606568913498725889277922100344083084041718918967310612899511662610752341812611340036795793408;
B4[114]<=640'd4562370947405160158871261159988375371622946773421904844305833321797179124127524685245114586032205018441688816006537217676678721285223450775373009103070825041211283142344838556456297041699602432;
B4[115]<=640'd4562370945479784936891055907554506343895293743239106172420689012047339982704135487269693282848630353557603402739219647968387373186894792294725626864613847302975212851938303380582489941052817408;
B4[116]<=640'd570305069268893327009512881556490496701947233354146950825161625601540091305184893342392717816600734406959196451014761529198161838450421377241105249058103254982861081635200267795587645030006785;
B4[117]<=640'd2263398054257342344361726389916050125701660076611572788312713034921445506492220442617872480392275399006121506470163635904833221720251568189968691368618019582162039688495926665951884089917177856;
B4[118]<=640'd4508974244720821787938428637198416624197948055873049375197010663004700405242431077755626572165902838998199425587787146340259373586048753921893687263284327669451102603431512622780072670689001472;
B4[119]<=640'd3700288862052788825929295519299367692863083303718086001384999483988969230749504889337412280251635328053221581355311029782122349569849211776001336203391875479040741034683148093601143383323082752;
B4[120]<=640'd4508903812086335437429404413596113015782854464452926187691292006750105385295804552743928522903857133549456882758399394196739029931819851310816877055842751841596082046573185106003480414969974784;
B4[121]<=640'd516786219344605209315603630532617164879577037857678800649233655607381683205053204397221146591565372421283432415679041137706309987446670937588901394863636717347075033425301022622592480261701632;
B4[122]<=640'd535721591006041886158574783912765807480288818539725047879067442570706023241001725708570602186254608236793779271066338444682028181052255578824099544256613526335029764631063669640901300474217984;
B4[123]<=640'd3528814885360022741734937291635848502482191016342964569515850146204890308805235706881970571539793144445907159116213716169221554599010636556147525722443376961721150554766132533802645259468955648;
B4[124]<=640'd2281221131817599596083945403054048152025855710723996581014425680021382818392185766515480391867225995707241928154301068236199386554800875043963753492322603772424351369689289932943092611650969600;
B4[125]<=640'd6908821822801460000887502367827787677446750033250404854374925134505822967916851241656471890507314477953038477222613774826178551518630516368364574676901707253704231768457392925128589312;
B4[126]<=640'd151444808692259097541087346793687470248104346002926957732536856503404954449555696452079027107597939352529918885568381627108227332553306501379306689968098095492642891695700537174903494912;
B4[127]<=640'd417416369036895932082420899030422500522319829132662478709637568027109004667890804282654337286773496289062255482335223452881205525763895297870501409980969509421826422164932599704724576640;
B4[128]<=640'd2281256100014128983618628214590768506045062515224870975818109526664835795900913008934098582540274264088512595207703130649712502113845805095240069477351437342071598213290966409967197077379227648;
B4[129]<=640'd516828131440498012574936013113195197737953559408740873449339144534748677165062117525221453056685557741628151568518556677203576294021568658371618499785059666374675476755153056693918269639229440;
B4[130]<=640'd1140548762959268705485605120698416798830948953687766590010178731214685887837999450758262124260844275284242143640799289762497685479894722751489889471384042270959144328059846165304381549335019648;
B4[131]<=640'd4562379693909427685448149008115086049759407788950768831537140787189446944154977297914309006868328854512183519068640300585724749737820229224413758176928921765799765258733467384894479375550906496;
B4[132]<=640'd4473330286982273214021183569804699382933765563627362505721033865148960509411587792337323389920488543193341481170686849932820937537315811625897321752985873385769053123457775895786040119374381056;
B4[133]<=640'd2535180819310832888789574285475446110672306539276808785829991862867716138148346014973974416690567660652829934061684106392605068768091900812467120337951961376282653826357047596310508656381661184;
B4[134]<=640'd2370328298066614585679530034659509943824337590421099028573486011768347140958217490064241677433356406641353228732573838324004602842187357892990594902789212685890512786394889038149540612004646912;
B4[135]<=640'd4500080631341917386563041953740015246584704177836172473463873274062606757887986870187366540830798602098324300031317480664827561498458542064638353608213922588073682938131795049614312223778279424;
B4[136]<=640'd2147101455716088803347204740369440603439251451595532222514596115618843915190679001061112226112876713908911117236619965086256827764396670461219113544278466944638541051881740639071116665886343168;
B4[137]<=640'd1729228924824602941539389802429318697710915861147859675572986746575452264247364564412088540756331244944057522933899658788611965586182809474117542934972585429672717463628586602316088551713832960;
B4[138]<=640'd4009996651364878032338980751185767389090001612723064795824945980306685236880677003947380690068809787382038786135757237642649510193461487592863072609703590323436969362068097416410424547364356096;
B4[139]<=640'd4442249374538004877074539212667824136632948763590144470932884600742069965284245272447104426801583151349725646725874051090040497893703737774301779423042162834175210538372429490692631987711082496;
B4[140]<=640'd2210078920122709462440294029592529592193832763418128763830591800987493838144175189725947629794851055218248984990098810314364587565473153250700861379984685923614480850491451222276402083604136960;
B4[141]<=640'd3635708397363430409151858430728887754792496151555783309149285902195833395033998906871843620553858813599912844894377680788543062446821511593594209482902975899967431562596748765341324377107402240;
B4[142]<=640'd1363385712213250964708975240751046887937407266196035053671922748408060768668714693498550142873772629952487196901263410218791159438086943905735730652559267019252570555330647854172945632523488256;
B4[143]<=640'd2237227624365370775981406755519241549431924981145053265120358512336395146285866896839134941626915527784520043368127510608176508529252187812690263232246737983436853799108993423983385378371190784;
B4[144]<=640'd4533549430270089399197465963924696360520536879728795416943112759805149407112764187925407010646845392932193304159438189934870218543775758178467046171213410315267158850692982857527888235472708364;
B4[145]<=640'd4542395180850762138930783238319481764158336693084644205753759481380643359690828125920920755845594725460286170564219867424566215391028321565616774710037563746797340000117182796303949877704079364;
B4[146]<=640'd4561888039288743755040362730171174096628895676276886856720345232675186067751965607118939737500480292622773003159913408376423861790116088965722183426709013406318450615785308627003506225079072960;
B4[147]<=640'd3956426207762057656285836023532225711428239945729951310311272315573182992975724462726544574242954243055714221245823610874660842458531935700790443544129233102019574304978246358693704580208583137;
B4[148]<=640'd4562384877743689992054091887356161413306986071935330330245486316640122791570111980567168805570010935508425309971544291766701596929358181250875538113099969701520620023486399616893815841739433969;
B4[149]<=640'd4553525457914525598696934986177403393959243805054621772784790288185238052050481965084364799546871903054571401146823787069083601200445954045125681743345526807418382481524592715257813012787986033;
B4[150]<=640'd2285672272871307099614442360124988029854359497678768144754895170983715937010922289951360307809964042991243464624371264934491939859035971122207287074003516337191563076724540375718423806338923568;
B4[151]<=640'd2284701038153061436579378425756208933863185389985945488862325196119516547902543003866109544952360765352175626250838861967326261485216421096084005341689411051815743580879281360398559621926600712;
B4[152]<=640'd9606986064100491257660310119468464346134319367969559443436393809446934589162702864922687201331372528993170287231919829404043250878574168056477870553502448962771257164619054009816126683348735;
B4[153]<=640'd87021648726387500882567405390807533166505262921136174461552229796231979275032886422325105780279575784634708864762790273966984437643924199572564147058939329826880145991942754642261876670456;
B4[154]<=640'd17830531870179882857170624360862677733246046796512052931655866035879590146543765219137919812619792854205117356535615326686149117374299305614496613490123265347973194573383444474246196528869372;
B4[155]<=640'd151491637147535834858106629397278852933310559992801183273788753719689182486749235373757878342024513490241669146827880713797240083674275210704032588774208699510052271968387880020368585719283487;
B4[156]<=640'd441095876533294134063545224876906124954222880645788936420619483164112266477028594001451864227209450679424340752294406808119049400208062207891039988527225823603448511279669051762542802146164255;
B4[157]<=640'd169378969214356702374533403802700946629088598730604009380045882135645100495764618401328849230504683515764093362606921850870897897390989805316173251485610392403891419656108129799021251155459839;
B4[158]<=640'd2765130297390834207198288060036599306351943601646436255152162919369599234238281052895861177740889782785687120486042737318379643275467309125518664455702629455369690780449150112429327831915298814;
B4[159]<=640'd444471773651528811746360797134212262147783376133131586721923044783653703920626844672814203632999504961502283585950103835043671402900258039801813937358100186145243746561690980350076198324273151;
B4[160]<=640'd231146938446644897208921830304118747154855740681419312377297321070047957835856324244555808985257198214036473916695928728976043134476248038370626364972006420021709252223416201721945377665432575;
B4[161]<=640'd2423257052392040265820617497913674390377140384019327469936832922799135300008169906879061452893863440425515312403266851014306784731311168584805411488254232615464467445480951323701797337817938431;
B4[162]<=640'd3559414961694223545095862787084840548202464769824948147404876786152640461073566611511873435396561566744635475617717256926746823529089140587406979885355125689939598833538462121669460176763091327;
B4[163]<=640'd1962332741432507011875254309077173898113453258109036249252275769684816452367506863282975114714354931826641993989067097782328386663125676476205324630269428604646551354955675834556845458448187260;
B4[164]<=640'd2254764912827514495726598494715832334242617216148195189911456621058902698770532028499164144687970018497467125924869507526822627274817445400168302608590868501760905478460740875557803368701231100;
B4[165]<=640'd1844705986147057654309128216773377155103095097939716040780233432263295066462503993779740825550913245183358052647100312626523090819901454795899619803614667221488845497570548734795954254451310588;
B4[166]<=640'd4055765090127893613790332587260440049504059785363226094076433752438642087362359240280483330049402525632235072689269175580020943329356694920782319234399854717776382570159320223078648358258081790;
B4[167]<=640'd1759925038197870428449897352002190492492645786992151055430697545990531899605711651662832788160085551715640243487912745163542585026860523530299139703325117335781163903242137663870546197769879550;
B4[168]<=640'd2788034323106867757788601894364380594956717249115549846103736801823677872201768687768519694057934301538396621395549764598118450564051947087753289594732789496856130723319673360979680308305592312;
B4[169]<=640'd2352369140841909978192418598226384013179352147601504256020087678155165072488360641688045883286866511980930522426158734147393184777165097010676933242056767618673420262599169145041419191860830204;
B4[170]<=640'd2919332599604657950523421995837495104926874318276950490434425562054371319769056319615833557571648407655209403272761658232375617405540907990431801591732961662414018951641812540765231111911739329;
B4[171]<=640'd2121935863959291809605731702090971134194562234894694546602370855405371471956934063791590379550168719357359457558612186738365961426000946633409259029499765167760965494867288043172383922930321392;
B4[172]<=640'd2108569342849523215522545423723406302343389880731336561134214055492426251384306475765187343772229774559345929533917957746306059891133682218431682710012175958494188810238968474404244058238092280;
B4[173]<=640'd4330614778609847445251403400314119130564047311759500741141821382573913199739915954617454955826327737478365211740306850209235487246756107500837404942526333169346848244471123446704831652234986492;
B4[174]<=640'd2325357536102453579150482357135757832015057703154110334351111151409120157566127514972523825530652040083619689034712048704363099484386603197032252557116889653731332032264869797908013185021051902;
B4[175]<=640'd2751415543419707459541608953245224565464694466289522362852818485111767215532832793602485500308269922080189640068898942575258046952841062523469860315404129678672649000831328186701647406010744819;
B4[176]<=640'd4445761854181971821437218345490874819528267423818893062577397391363955573518335371010260320544778612135341301998838476069944939058813866473984472175530925395373529361662665268307071314125915001;
B4[177]<=640'd3412500790041262277514359477504517282943190115360084621368594404526935146576302110612620438338279765768116184990559696690328835999560510651635931818051778944318000696563884903770056626404361215;
B4[178]<=640'd520754116420022237008011789441504619244817759819449749861046288215636412666876177095288809683205507062590585571066070800647540651498912728489666947124574920161154162888114194275201404316452863;
B4[179]<=640'd2717860624481708477079856302328029262435878616760434238535846704860455738077083884222531489146806638208177049912379707876244515512168125957854350392477152632710078960041039758733239948516793535;
B4[180]<=640'd2307988320300979882862481193639386220037532815670780618323171528215365933681092069122590239893639657536507363821219422309926422211070858902378779484437377056026159927331295066628372399722071039;
B4[181]<=640'd2299075145439424162304395581171290048718582385269307352242742343336939263441724234356622907049211309656421467414613122926726208575226527633066809002575889984207243914650500978587398641738056703;
B4[182]<=640'd3439657011452066704228251376630724111951710400144671530841888957731850891580981490809863584073132336271751154786365546374616520622107542899818904695131184246236835127248710446948458697907503615;
B4[183]<=640'd4423206992235112038545995534985423768251909685837787943688391642578511247977086833547128995670991292433741466130476568583472354534978667426342979540180768350726326784869277167469075850418192623;
B4[184]<=640'd3992205300908891627187829111712805831827463898580271937676499268177499962963079412994880964803997022423168991474894819861558001640641648580301855985223812452988756287963818638860855038250582271;
B4[185]<=640'd29772709373740197780875575635083037052831268061474946692190343661918589148018375007053731231554546560569840254694141408813703305843619609448663105023610010041301690744922304977334966527;
B4[186]<=640'd17822063410447604505504305796314652929475807859601490960293417436101899835243301952543935406869549320109401289859417159605841235394237806942111462352032787799467917257757067204644855626078335;
B4[187]<=640'd17822170700128088166246384349695296197373073337016887609713231605936489437427250524824703500364440542733308082587674589684248204136585929331419517584255439325928235018665942196747170939406655;
B4[188]<=640'd2281220445848614240630149258743406173161582511857456262734067650544402369161091620486645517944467751529851510877388685781799954869198125139158165163381954453698643728745075838293060804734354239;
B4[189]<=640'd217206035263695389402509002591789916538835077045580510124505626940299270702389385721930817604789782861979286476121536106744600582642176073535595426299794892789206038977825205843710762874307391;
B4[190]<=640'd251736225485050702950312367855365937779885394889386283485922135111381300040123930335935621243062980311665562746265759817168217070858264096803479377910506086027312118252510220494806074500579839;
B4[191]<=640'd3992170349237636069285238180027257450159420944655951236061209697690273664910526217970552658700981610772054941061472632496487978253383623822217714706278114945900917712641926960300533758212178175;
B4[192]<=640'd4277567636129767626322807041834385854687562286514718862413161523360936666672920528410535846106129756161420300054742126440432622529562645422991638962044367319171666778268128000004857258307518975;
B4[193]<=640'd3137097260247641671336108969648380910612918715467363029082456126585406022205319202958343931986665995398761189748164378682607736323214002210502525510592340176240899931743018830565682174377341951;
B4[194]<=640'd3136871544594874713778342495925226509916990999727040005953481012604803308091482925789914248078901048681592380336275191380340092567372498146266909377851420351347124753066131943088623491485809535;
B4[195]<=640'd2566427235940906876080833380526696683474305067215312580176232288316765580446902644704065254612114342127938329372403202692468697948396859508528617072070829735878098145762023451454285751697638271;
B4[196]<=640'd14265023767910836156466421364360772887936965139056423757947395404328292391339089097274649402289136086178756838683215860827087866116306557950009982948599640109830281223547151704647066003293439;
B4[197]<=640'd2861550279948560868742234955953521182192118567596438426457263589062528345841759553731733580140145474811754618352226869629933478325842012238923078339837679917754575518924837607626691438192950527;
B4[198]<=640'd4403991598030315573618416151795615500735700176128400549704169194247545452830902179331736360402832429100671972266934219070949452081455109916035056371405573224284108864940294382245951892243906559;
B4[199]<=640'd4517789808606402744122283633936554068629830594013791540636896012741661965514962340199007151410853698313651734013129936590174445811800131122980692654669103169220254377218837039884385711135224575;
B4[200]<=640'd4535430151771182515998858434510834869615024105965638298382154199661285099386429365702131931896946288559514493363985217060654835393666540899783776531138096895652664377869226182541259092110278655;
B4[201]<=640'd4544618957882823268634303675133580446350570257535926672740901565190873309458706911115984803906054377370357365427757749368351784267318397539781836569684238991599337739641949615048245885156786172;
B4[202]<=640'd3440766373984182098140301462486143928266243188384171161835357567806017656222060236901979816567674615445582292574772283559409671900676312753007980388638031551342963505198562521129780935183630335;
B4[203]<=640'd242572979174576205826702937739141691622481265664173021279166012795450265046970018746336444770815297552480282712758489830666650411839396915644551405348064665456968315478453306070178927280079;
B4[204]<=640'd13642819114739980464455907984943750409772799625874175849182040778714809595836153430673904738495800349718495978374879061998046273807677295746630791921748313134207338742797078612223316940619775;
B4[205]<=640'd17819960564669271914521656734692552436726291841283522866137069078517911018780285053109893438120218533865993769946601197660315801101073951091155823545211563506362104615711122870503727361294207;
B4[206]<=640'd17822033661549321552528373423306018220851615944340928236791407795079861046679348418358668186406792586127810692045600783513122754148355379320392905922386451156147226409552537350686246215221111;
B4[207]<=640'd1140401302448306149112230677346321941219708768955471595559393673040500842529040290892572912017779516460157723923326287421333200960073004404733457860998232681989534192599366165185517624835571711;
B4[208]<=640'd4561988105048670240582095848341502584815527532567938444435906780136956397487203296050752095754278805182948013209206046629145765872288767491889248011419211964258417962068364343043682831985311743;
B4[209]<=640'd4562022913708220222726812385220166561245640391782822934812977880289007476232802597517719518259359446464651648778359452489517514647437749235896836610548032946819876547347694088247705603489460223;
B4[210]<=640'd4562440617614932033067062161215574647993940309360858009722711930709033722111364176501281191831516863485201625389372932358374664288548081400761638702478330318701546135067289303170019504372369407;
B4[211]<=640'd4562437354163059548797503556190533139557018468604861664193678684218780292578275683302402188421874403852998410032608236060244738222070079712621856873722592484640277179292784044368889805948092415;
B4[212]<=640'd4562437350069562439107074852255940796911614722139255546249625008235284369489567090290027209274807511436552000589040726260879128235372006844731167233783878985339914058797284300431878520612945919;
B4[213]<=640'd4562366593986689238059818898174521560835516801198579754969750579051318431084980708829613766455754037698734134897406113799649398100752194907211512060233538747533443534351056248164721129738600447;
B4[214]<=640'd4551858377221130848796974560515536637789479908588968643600820149410431937852691012648905361525429186135993154870598393480574272493163516998348526720339249288816395851735251138760291026201735167;
B4[215]<=640'd3999331822889952162852407846251890503563901243291207840310325054760413821917895664589132326310301182390705772206034163295790933584453355151964495041558055385852891230428616822311727975955636223;
B4[216]<=640'd4063458212035591612236467987432676324080670242495793126555670161478228462127610742352625913608693635813497519947823051481431195675875700105663491734153907027566920174154861769656541088365215503;
B4[217]<=640'd4535724427692057720426159394819251106617056876395651994684148320756491030427181228688105432258159182934053830958130695601380669391910827471957009347366147400128359122608172061334726547667124199;
B4[218]<=640'd4482344807651451899248842315091933863071196602149507189959193474798846498041470170724377582114702552711367816842000964777173681605818776676666895274754226520916242584021867394029594211340876597;
B4[219]<=640'd4417201487592013273536698955089736505837514564669737718002550492555228613864252054445418520231711238353961903149161660512132796538322609729370843263845261440797257325097485022143503288460934079;
B4[220]<=640'd4562439530648164767351158252955007701883070029157493596722745222132152334899891315292124042057455933462231877699301035575269093603291417942192373124889931014302481958669486580337991531474403235;
B4[221]<=640'd2254225106662591650320414612161196685933507852398008634335084486971523307639194661871458550722653475506476446402386382892556235428265180153687559787669154930479371132007103471838795114755065735;
B4[222]<=640'd1391824251059388905831116046403755377427841923271696372613100196728776032066302697372301696737531772347744620084964884211538598845548563916724914913426714873284069194144662309144066106212274009;
B4[223]<=640'd3537677086617993666666878374160392567357685339460292124752768291793314066254804418629665980586911126157701987996677111837065989520673297316790460665384550205031043889016364077782228911661608855;
B4[224]<=640'd2441619353243003218866733133082784314824443818395459428011588390429115782800596477604734901027748420899165429199822970105927304011956416897114789941070864413853032621765453850333232048681583726;
B4[225]<=640'd2708950204483786686742371918770322434015983094527555455295331605465621389436807421483938843162210293720010263014956743894684288043345468044715070130602356709768232187540637518340750150205582433;
B4[226]<=640'd70637103939674424694565641872237752537323930599296791259364199929348022215492767550017222923482576862208307492937431176330173761548014295891977958051553591684522369193274379481511305654080;
B4[227]<=640'd106971361717453777861911930180045306978589452757546420045561874992283538469579124624731405520566251290428506668828376885215368072999917666488178125895047063454169074926625753387766955070314101;
B4[228]<=640'd37645565246264640366107618352750004169224138535201304123619965862848301112290605675519694214867900943415551429148580524371038675569828716093441132446961044656109450638581158574710467229990913;
B4[229]<=640'd144682193200276599205675463444422023225517017564345258745617530545419796900479304145891814585163043005614215477935757291433484582196291594795648719254642982787438344735601178408984734479840369;
B4[230]<=640'd714987270403051001647892102291279148167208642217448946003709767005643277408904132952944212848311659726968778864044565430967012545489553824887115605964743782056802566669008272929589452529602273;
B4[231]<=640'd1832275605949033218358826034985411171021710975540360251002302115271152769167511109889882652305269566383674658250938012233802105476046151931982858821377120569946143177618704215585201286829467744;
B4[232]<=640'd842091090557221515122092287171432695139388475875583591249257653862082176482490992526430905337416386644432760551417755364009893082576655601516056005159855458722241205470427825835219647909603667;
B4[233]<=640'd4562440617622195163237229639632792002663865942452588902826440228892389427576682172792367692207822175961815955665223797715635399489525534511206598545450823190689666850657640641517097658092838884;
B4[234]<=640'd4562440617622193384249552030980678150504512404500397187383435318322848409013775575502163018302333210555543679246806557064503789451212269549405794953459720138947378388075222978258636531774384356;
B4[235]<=640'd4562440617622191237394615422804488645339726985266712925782083845119613311773364002889214796384116593524817433901055975604632955429128375373333408905690273233855596810027226445778480627793256485;
B4[236]<=640'd4562440617622195218393841322163400094083270889935261238185768312596468773184955779483679462809613781795828715449224344061063897269681463041857450281437388740680776160078223991091392474018081854;
B4[237]<=640'd4562440345679542895498072272257916184664984077823954294557719194529889837355680696767127822087332478925794824083878959317415482049545928424333742394545785855919019882557100028635353320086281080;
B4[238]<=640'd4562431092459000845241493385790140418707546854472770112327256698525612108847923576532599233697863404967324396486964683629802526228225832644161312663466555207692093796722082218731234640724603177;
B4[239]<=640'd4562336191710095685480952865415124459086943649392737791685747168960974547098330249629060109463613346373287455079899358832708131991798235600999924773592476053970313825594287722426349776474526192;
B4[240]<=640'd4562301382984450852006150908306827928498969135548731489201801192511377891641179021412549250140991628027646734327866548683923043592701036429017430832389651647186147130372540116267910682581850621;
B4[241]<=640'd3564128263241362097375683301112771246705390702620500942692842410089396181745647834785440692602866931462761776305755159716124753986686537266813357889253292699453964485810021455082667398018193162;
B4[242]<=640'd61832600368275254834432781453882113745280144130707190103831347776558760253113094843324132693037028803733255670741505374425116601371136623341818564835925489975239989108563798;
B4[243]<=640'd47796600084677451179739625287104916423894858976988372145320849628679891798895535847614105591282920365589409977381118336890933162979627044570002950510729691799293923079737613810;
B4[244]<=640'd47518353383020208578921560002454148459583541716647948791173549670394127632311178961379872522722549157503580665177904803833577464849748929821125871111259947154439896557458978228;
B4[245]<=640'd14847553163414028542287364639171581933831033526673680490712418636827643066568601967472955572149147980153540440233172607186836290002825215595361625987999816246036568797169283602;
B4[246]<=640'd15550898878343355561604772082841374761723238512867948811496506084885646323780408076196157506164865761208282803620950818330912756805155972190525197123622261677827308900363974902;
B4[247]<=640'd1978612551075948679424103873665105236601691376036389197379318003309897576850434466120082681485993505132968543941852222401474545090058086954361581101556324527962594568551075689;
B4[248]<=640'd15595146276120956070095622991017242525510989592664599699491252008187924736087258778066400476804035016413344578189552371088174814271563147196540311215991812256517320925747137422746318723605885;
B4[249]<=640'd3674682605374503597385173194856681717232534965918080024919417020936008829415948359629933893966641224416535105662780263901369949910281001155599808069881899145363992242449559351203666557654574328;
B4[250]<=640'd4549039250785210313869938134971426798672933190631320625563772936535473434164480038726078023908291492211781269824852730376496212251134397782495658827491892238312630359862345059478703830223814741;
B4[251]<=640'd4562440600625779511820211606286059321752304898623407315312971227743891719912851223169405332266042905888259212182133970833454186378028356020288920366203037836133362299427901340248633587760367660;
B4[252]<=640'd4562440617091057447432442104058529794361423387658430079453731953909078857357071745034737258965716785264147405407538665301482879772238994884264404613590499372122907003518940099996380481706899063;
B4[253]<=640'd4562440481567878762000316284375401874561277949038944820254426808759521947797824641830497809180626600948079798872333605590283998800024206785664199479261586755356996056704165228895369040970449464;
B4[254]<=640'd4562440617090797944417919013197069938659364945842002571529222146872087849571908270567274794311707981387068989598433120905898129494956088319919701664744390207868793442645854701064804981352469734;
B4[255]<=640'd4544061645391054621915539927788501684657940820794381129842422732395672970576252674543805252008208915514979864514894958622923107171595212025903727154664301285102043520043001540401813430314682807;
B4[256]<=640'd4561360461108471216017484231163548362774481519761457203377777419037571583335607516480605933810055886652171877276237259452811477389009934843066865355374427100151264688462056991990617277280091891;
B4[257]<=640'd2281460702501943795323195900104134615962189844460646700859487341659911987665175462868617063823540818153976563253933894492706444288807484084078911198712514479455955025404042328158220323068705939;
B4[258]<=640'd3422052774745663427808377016420805346359721941436702333416976657081616106189440449227913159800212271173501814097619974161088848182697149945572120755018909659354017507146120383742750175468373191;
B4[259]<=640'd3421863436232122896270900386606161016697099929784854539319211082508889759986663148731203970422186886267214185971017975793703397018087016971979636034656141463050388963918898760117615801040111899;
B4[260]<=640'd3421900080519042863634910552042809834718679057896994881596971554391528042429715195420418289857256273950393782598490961655878275577799794564394137640680158434108661275612840721691437107606765572;
B4[261]<=640'd3992170349062336203216313018167755200095242232888171265039173662711246896614542497121290066765721756647762255210323859178988208706622301800375390829974290615202943462356867232173135474735773004;
B4[262]<=640'd4419866013829228200476577910378277395375631639717369464453026386885037112995265915639392897198853093936120966434408227718075628095619313467523728304467978332301684834978068865642459100243493055;
B4[263]<=640'd4419865571663268159999655514107877442387684525242232020671608262119054068850722197030531444611605631947793454002768111772126153371936384217690468180229757995012514079700724039676704583114564150;
B4[264]<=640'd4553529872733067919317853229424219245593154486545482263668767342526234243590484461664548822204346690331953294436477761691373091308928340264474539956513036086990123336446112206168718558924030238;
B4[265]<=640'd4557985381149140081766522903477920012501602285725179367353512949308184336729121768240859779555513759722470492911173431301631309849828731236287515391076372364824082320622945442900090802603450635;
B4[266]<=640'd1140105700785487149145665570994228643776481502928353348459423811169446814514766425375896208137832841181028459054227443225764208600139651133539995411209207930885231960914249173374441166563549674;
B4[267]<=640'd4455507888657691237656418227936724996354457708631456793423290157273475287337741256710607262384548978149190949828726886760187840957960120380358900066510501957296199208959588627780853911109120;
B4[268]<=640'd4420978224363655986918704839811547779278451230530072454669200360721242984981927028017372827277209922972009361961001473655275806331004896537253258131557201955005549407139411032339758561779261749;
B4[269]<=640'd4553538301893758651174243564497502118665800623288839009889853683071460785670460304101073016309687113475990115158295915805018090367187897864852701816406040359456673145545126539846593217533133044;
B4[270]<=640'd4560213950135380673406015230503404063773274759637005139471540653412198158982642475132229101261552127627913973482506552681541605293747924468422761858808767559784699256482656851144555169837491464;
B4[271]<=640'd4561884766839000872520116639079748355379645039146805923161396075976616727682967122057291605458394323750455057327294413576744159389823514047524866852518661346872770237853691873045640201085464644;
B4[272]<=640'd4561344144847902500564662991110801860805830626811550404850700794705843254477509623808176778640159691862994848287353636071484894011568952649577276464000592149058718113265688577775594373477487628;
B4[273]<=640'd4561335442679916050818545255723343253893719330061404955746109170909014022827738904891782500729599810311879183857520396141074942793027213407016266469374311285803555854518031544957971692529060513;
B4[274]<=640'd4561888030144377508105393776384684176141042689778107310569309092664219976031951751454845012885968649941896673314250244193901519544119864218750291723210795899975181763437706380556898515433042006;
B4[275]<=640'd4561892381202825276155685775811768845933920777398497334713348975912334488305813171606348427706311105406779894361833877457716547173481810366753752951012797968217862078681539699278498397217227448;
B4[276]<=640'd3546654316173618121426230151044041567434571298310134901296010318069622754679292580018423171942892361514089817042110468398664037280437264043685521848978042883009095877135725544763795574464514030;
B4[277]<=640'd556938551696489654220471583366936279263935628019901329606670782672663999476797320922681413849281923520408862793994282989424359567026962562500245060013061784349723163300759208756412041246670;
B4[278]<=640'd2281220253601792965358974489842559036035715139403688239866096762190229950163507920238414886543609907343187246615452630369861047784593752111061320944960240443309015101029225621403987456364327849;
B4[279]<=640'd4562440073736890574271662547561967815165354121745208908344040379512478215308113775384556072529436470846218721038623887114766474029612577575459353545490877957525085765480139568659467356708252704;
B4[280]<=640'd4562440073736890574271662547561967815165354121745228721153613101080235892440570072566427463454441265195060741206497958275367736885016286304438195349578814882069321691717746471528644775948474307;
B4[281]<=640'd4277843929802154563114355797710650058975023709971845766001352926764130781746956069762966066743759191756461359041376505522907487141115145914878794498685753027835459560367915358273912829082929749;
B4[282]<=640'd68529548385190558141325428762225712172573422421614055413580087032456367504114587864593766250650919065421623375774187622520276156797378437797888776364327005604039065591035159618815492294157;
B4[283]<=640'd16452530465492177649008684286169268200161476414712726912549252998499837625743546054820624260723530801697313493034104117751489073738279901230856845992326760475025829943552335525610986318084;
B4[284]<=640'd135971326161092377264534580877431968596375838138306220494080066340304878421400613835518357232865111412876370868603672805721270325651913443681139504636792123515697646516212772150184264057;
B4[285]<=640'd186069449125617808859688659243373913175598978053566751715008255495528512404834297123139000610173531284587116768257938586993069527888058812;
B4[286]<=640'd47634102081552798814437079140779119159192034510077115879117020125123022875062809131482095039722589682190789981666321327987731087936773480695;
B4[287]<=640'd47633557485555325801728790073357577301341424589379305209820019721197927327772692450251350253871912829431460605555053907503117671525584870507;
B4[288]<=640'd21491165836327522650258880588454432049238849361585747432482010378419741359631975547577789713154181804750143173747774276021559202147148783535;
B4[289]<=640'd21119025884754307311700141973551098510794348817494187895384539298018505654843210923634094059177488523400766241799139316746850398116863437320;
B4[290]<=640'd585351670212852551696399994379075394784198192113186678809393323700995576032801558066832448541177886831435204402843394738312518040671623972942941;
B4[291]<=640'd1463390339751158144466060652010579106461099653362207532123113012766665385485898613717376902396031867568234026939094090784092701277699033049075065;
B4[292]<=640'd1524291284157938237510175454456317313318760162678981221185790309579122352554817365083092018130094917948062786910828632507674871442916790176325962;
B4[293]<=640'd1560874275078498130220965975747493922838190600145057796438127705486296624155608764996409867798518188561952979003981088720306165190623140139503852;
B4[294]<=640'd1560874275067318726014270842670874235483907999878782340428701960537073182403934094674274605376183980064499736144160046884431090396231538260322226;
B4[295]<=640'd390218568052546991917786455459628729990705453789769336221491693334934907258994838452697943519533388128162166869105720996548551722641657706956897;
B4[296]<=640'd1560874275067175240357598377259642646083829452559232209095331834541497315934290351832021222240251132138053634761273157129748648829464762844188194;
B4[297]<=640'd3121748550043816403403488909375914132415617322301255658237047657429130199867563989934497696292466037292172114274346785114774936112775123003073628;
B4[298]<=640'd1560874274794577215880250522122580016918767026538746661442027386899602601074549988499594407835721205839752293792123707322340234136039371106459238;
B4[299]<=640'd3902185686441323931483788523407145540180945672466616009788678539954313994346652634441948035649432183027869668442991545768968742012625207223217744;
B4[300]<=640'd4682622639403313744941978763360960227321749694824820420578040559960613119237648181930224136593592074830938435691438188500672196899211976074921749;
B4[301]<=640'd1560874134876558541100413983627194494314814599718076106674906665854362754885813771838354827055866335507732766341393385378835193286645194050611740;
B4[302]<=640'd3121743165531336559583506989511300938011921612718724347880949800727828954172422759635202318649123152645445208223546005336895329957155500852517156;
B4[303]<=640'd3121743162740744350242532214408953620245648265150064031259641696580162652042865173553443328595962215488984886490095754701717744133766973141375340;
B4[304]<=640'd331961245510479436680992629095292892082556572668845654056567745971887523593600568791181490335835095181308547109293313330226181366456641527296812832668608636191977261163544397364866334;
B4[305]<=640'd497941868265719155021488943642939338123054421958906549419472544479865638624727363978252912195761076313941151040549205352023386221483459239291030395852213970265743147569291818661197146;
B4[306]<=640'd500016626050159651500745147574784918697389989508939144561283282280607734109341686055719948109968729745500456767599496310133504589405716467221960489621321043110691817884922183123576645;
B4[307]<=640'd1032710687205257122549775507076137731458612774607223399008275644317183744856363543287528986170773353705221118519426710076605542108556150533202713702405648586099806078161770409481071159;
B4[308]<=640'd8771783255577084613319442293183890853466839185954005616973975748509292558687574879804432469409616843045987092765559863271205030357035958381198765380010287189693032876227168475465370379520626;
B4[309]<=640'd8771784317836861201662698293616114865186550247089207987332290485994736687292327333956634449977430432436872662357446268244264450360794843367831939854354380415861570868263786315095726921651210;
B4[310]<=640'd4562438714023382535207721371567438791044496720188106822526074865883055864540364436439169991984813159684081683216294898051231769225823943601015817015824154104255195703793817947174393417884503224;
B4[311]<=640'd4562438714022604501038556185387717714576758531440385035963038276706760549113560361878738870184875431927252215405031961244181435421462002139510485386598607591541842399294163890157865065047404769;
B4[312]<=640'd4562440617621806201553690594726127120951747822147946408178155998549377204455959468531116215761270881952462688239101242600847836917525272117432777784613140275408464434434114665029262251205613096;
B4[313]<=640'd4562440617622195162991831288993590462663401926858690048302512955585678928193998834882881757874409560118188478986326149164130100775199547536030312521898630116684247214686620021287188144316232832;
B4[314]<=640'd4562440617620104251811540153147250671799046200663876536159418354164813558306479035487907045771817610807646823190958072625153725330677803743923917312238195991161650275493990703178093144567746638;
B4[315]<=640'd4562440617622195155309187302671873738411130906688905361495755109883673118517636469624751328981881289205157535456723984526746430710700780503797255811516875977375913428349358048451477977740100709;
B4[316]<=640'd4562440617621182153316737769528782197554825989621942860132789662308654542328420659153680192872443632509584891231803645882577272205278546371591782480912807012908125604609709010629597345321485620;
B4[317]<=640'd1069322087738660654769245199844311446999975908888357443536620352655761998462478441484653206981362652712468664577424795996469241289934269224921207235066625241463920575955409536731194483819818177;
B4[318]<=640'd141671244153911251110724192824446099527621653959669228805902976379509170427546209086066121978097360960917590462209780399139943154329278063096459346225658963445711958876704795103689805828605530;
B4[319]<=640'd3444036212965752045716604688918567637519146315145272819463865694361085153164457172086234413450769037816399687253279502873459438233380045112442766139492631953881284836569785545050106863039155482;
B4[320]<=640'd71288134650331097778739567136367896808256292871080406050830584170029710482089630615045138031077504229134920402751277691697699917316492502878295029283643166530970533021467223301092585644238929;
B4[321]<=640'd3368356137025913597528277319896209500079384106113434957107655084625126203212567613697676467918082690182479371944980606504033835090882004877294522244469071634244990605577395038877688321452277788;
B4[322]<=640'd4561326740518514528780587914740730656657544198401455847902489144945932799903596836161262479779923367337676447157912898969526769496751057815036673414593131952486929446811179962705171626451949185;
B4[323]<=640'd4562440617618550209603009992894221296220544873586074111633296111373888249118500011943400223629951038012813386665454524029674689053078591067929859640901346779654046831005400913747010772820978272;
B4[324]<=640'd4562440616560162875094528736768037616255978299327385547932354898752581706206034190867733858844547327064860977355747860263846356353422400553108381649876166367743231405957791182026856408518498388;
B4[325]<=640'd4562371000303200992363016644712900858880126752673190035665699369525514369863360871605158490307246756933500183382117570783721648611969294315270642898825930615244542809251784167820249954569441429;
B4[326]<=640'd4562439665822920195269795823174492743355554583397168844886907822331266247173260934276940703940176494880247525154949380140637968770090192974323232668313540647874588343393182812979020390677230084;
B4[327]<=640'd16847391196663989665254491235932796576462830829018451798370095296447476231980979441703268745117178607531727124975966830863935476146814106954948807321361643315275761864845047817518420809362570;
B4[328]<=640'd463372535302828970008247527563683315800029219359033032148572321508108344444882208307705002320296723003454147474837285013431038289498320758915078583444492996697894289326764275696754234043014540;
B4[329]<=640'd891101412248956640989051788971427699800134421337458842713862569991218018676620091321794809038317009008846357213594218599223176539129991035629994697162525898476085187241640363978898010667234176;
B4[330]<=640'd1782168565035104730353545116296875586022677105081474224309013472111252759141163733051937684230910965897602959876255850820006924817329237046558325867449926693960719274985288053599374009653401159;
B4[331]<=640'd3158398528143611572652897030650422047352128376405298948086465016320512892432887175008556294413453170880774461244849088480425365930386021449032024747318607099501030402462028887751313560979918596;
B4[332]<=640'd2321257337210757809266864235710212014491828235969953456616484144858131302347368095193102482457791977368551431285609595208699477434402147771149009484050126814816799953260021710230766011173334028;
B4[333]<=640'd10585367741641041569983633751304861072768947693836203516186636237205795624145327706017973182349685565804474901591872725777270985966894062971733710503338769270486514639319986424719225294553165;
B4[334]<=640'd1069443850063456557464557607613141339874227658644190320281245435632012621209051128950642652598515196470359839778131219337860755189344494705306805708632698287822446763191587826590535711929796120;
B4[335]<=640'd2270360211004948096184605458308771597958048806358013558338982289459219196450489843710827290912429641806722168045542487139160243354702227567485929137170473793080320230683695765835356127454058212;
B4[336]<=640'd356413211288820096713831933094520373182113468193057268307318709720349386234101414581360705775011057889804620849057788540481472835945866965717697880643804729889892822516559189619891681095985232;
B4[337]<=640'd3773823839446102687638361707858035254008454767520948390906808115827408050913595422238614929918405790675852028112481856595255198389815178809091032115261475909147574069900386132766907849455440496;
B4[338]<=640'd54545687822855518489110897226233177410955973773056369977595853577262158797692152933310444333254801437881478294779152486303700961719401913949342189876078931042237444840149877567670647423248920;
B4[339]<=640'd3453153959857670537695271541910834293585192098283846427523161332958913199268964679147249213701356188339736844010152323872963941025217394117924670572451617147687324764377830908591526372404636386;
B4[340]<=640'd2530728478400899072325930936593290644239494075659302591535751774251469782272275579011793675474707686948269676316456972213779814725121776939698892149224469661647744806016953358691508113524937752;
B4[341]<=640'd1425831502996181403636535560312676324444532624128123029771681016707484044520168027666755179194247273539980155943648255311885669861404007548495016307601243225714432024912964939472784273308916333;
B4[342]<=640'd2388186898784824738526525821057591273402607123939707811514003827922863264310399324404718197918610260324965626865482099825764633878032734751313558944744503221794488038947608465522817334588479578;
B4[343]<=640'd3813943273374198196090485936497627164264950319615178705151620989655240950015825424992700264070139943401212556082387013535708331659274988816046753722769396371025986947487026976181262469432411917;
B4[344]<=640'd2811495318177613817138084339880166485785000961536962822718762029857482683908146584764886328787351880602551117946969252985591772438651311897021921191754846428645992864953032984811343892240335136;
B4[345]<=640'd1995579913585486569160089072113843936620053007938236689482217558651238893746820478591465460352777263451639834112014013769082082487895881159710523823870404130772128764090398800981989643675006985;
B4[346]<=640'd2297997827742530567887803882851434602730717142839122380618851316583240913448614673356751715899307554924797285533531384704644702539456297243918404826851472458051996693906973245165022229572355622;
B4[347]<=640'd975790879741649307258525832707830939228569922149611245278617839223636067323233306905450961376376395118686526314508832024746588543049944505794648153885590159682796578441871456438050129902186848;
B4[348]<=640'd206632904674976092598486725436278682972635861613067550648822081062263102018206808080206160312713306562493027684103166356239178752126729854153071175238831836468400138154663276550772159629631783;
B4[349]<=640'd1372305267876122015098956698599410860338158064058826621988128116852862783780160506210377980348240905532194673828531514987991351921979474600150890327930394228192104384272866497217769531947352192;
B4[350]<=640'd160402517273535796854412076750395568136203668091796185939877321749132974012801164607292334683820393761548629310174759230561317430919098869218575330112711087135986059500753238085477611127048232;
B4[351]<=640'd320798779340108976623922291781973222539002716486820492923944539781170490606050367470901863714837351190494129545816450572511605160286622242365712954452167926810130848812627216304276141468816240;
B4[352]<=640'd231686570398113148330350868593127984708662232101372884917445994147095733191816224182802665005329879597486119180179581367049619356793955600953358990478359437696544182516104954302035923025673607;
B4[353]<=640'd71288168643170307272681477854234248488892042818580530828185251534882867221434801739314265660944415448480231000178444220222071661789680023102082397096779619381847294749986274608395317989364924;
B4[354]<=640'd298519072346527007533922623953449355785262876327791049788622772626434787053506195503351780115763648694218917053383810127978548459874633633148471033641232790975013225899216131168179375444076035;
B4[355]<=640'd316480335435315401602191494680916263411242885466257287206035014700457118917148462042879988533974010755944350572016612595727094460231691683352298286318442269690829373544682405169763083307983650;
B4[356]<=640'd388708300605837246022911229121431126556706947545669512658323305985008414495205585385632057693708784314491299028782984130942586746084891178712709340474434868801403686535876284881252562531591462;
B4[357]<=640'd748494956251590424088422045979670042950460008215785736511601921234582736294366732585364433111595534945707525605508663223712604070702222791158042477535687295588469158511891931195835133680296492;
B4[358]<=640'd1888802710427747908734228107530603436483590695792807970001980929693168207757389235552164678037216441970284148379178224113474996264991094348058102293729991919469343825890003196034815671822195889;
B4[359]<=640'd177112986145611097795407968315964271952119885068841562412182727150290969632399156528474394262652058072067673963621531256072627534017682493451001401530777883925078029179912742524754368608085143;
B4[360]<=640'd2130899233871746760052128724614515820856753321118633570695943217263637430113043664180089062849636222953623393271796116881701954913584190098417450558860526009833958210939296324787162975679293839;
B4[361]<=640'd1873476729358902984970477294101679153220421740177576899293898501570097181818881161480711214730696343636489665493850756614835116148221345418302549183130259912581642154197025041069656555865244992;
B4[362]<=640'd2630125469111758465064794148471825444608848914930968277932729124110483482936634026019460997812285721523407611252633520915407047710925897758424358305814610650123943388925706242465292437726189577;
B4[363]<=640'd954972204564050318933978987667962028824556973744596874267711827691205550875182513943394862383855731074021103350631745645026959854966412878968784394751863153522442716658851245841800789360382600;
B4[364]<=640'd3536580536831350523619588758477537987708384541637203334777565716732961836833001356775517692114076864527261053115976234958698772908035509203387005677933272903883961067093002299482845507905274436;
B4[365]<=640'd1084047057032988091679847227432031004534817134504264863623785765407266365760266278236331754900836222419967972244765052106415704179951252046851914269553331618070123871704552500967985146753089647;
B4[366]<=640'd1596345520221384256813297196627279019787730971510556671826359467733338665347963871477886969213913092954995151319938424915706958214558623438120057774233270546200233433027518391306218973643674177;
B4[367]<=640'd993580001296521906616075942150473161014385865402492984058982614070245241235258206210119361437487570896904972700780328947162669382163950823420685546043661915679514578841979781478815101400516833;
B4[368]<=640'd130168244341920154278825296349849145685053364900654770005111213440012919022363436376789265614328503981442805976215175118882302267570997506363091126017435812251420032085509830317572892801;
B4[369]<=640'd10854789161462376867984870093156600538006090695165055438329397163156825726276694300516836441697070185609803432442231346017166617352198410038638109680552641913527355381589569938504421448;
B4[370]<=640'd7385654283257674810057161503751759548864468969041095361080874237699475807937413657216452661446932727442825592400512854722943481452890256335659132792392854856416109898903913664035881408;
B4[371]<=640'd69599245045362990834814426422999394377985859986127719376306307702545651439425311152275849220866859315460154852008025649438407732270218540619450612085601524023568506841218565158782369924;
B4[372]<=640'd9605049495317229662367787998898344630489389523405973935107149989548091385472606418238163743090713596705479160323976002039128431076008542723349259266005614090823641163059610746037997702;
B4[373]<=640'd9009996168588770494088592882763107671360514075206910152929785206844495516749691828525834189474963172055494377628553621803369868496272808778531293003809132323463271105664113990162579856;
B4[374]<=640'd29808114990934627521379049220189094321882085403934721909710273327134570612777832974577988512037382845008317210085169359712632035440638224557800078233701541394119665283208341205616264;
B4[375]<=640'd16266607781030191282098465559417010614260902772201890147858938369588755649026959766727772853405495031875610072848234243387770477078937069528692656731918181225892316654335105111704136;
B4[376]<=640'd7556513026811736555819941521986199928076083924366493121589582252870042026694130383944243012931764245670802587171178961282615715883081147508935056860618525827589897633567856784245706;
B4[377]<=640'd3959174022859731068220547697020117138825450902950342845597277550212599058022039533642208349404574669567916726256032340344189851923356082534305302030294052522053820569564726399280109;
B4[378]<=640'd16216987096703906538728031205829168979814835622600640314368782725279775579119873069371165015023860465367836638546637081872849818364061389894750647654146893077142074557440081281064;
B4[379]<=640'd96233300311925119131003675189061638103799005585240762269746366827218503412671794869828081296219842604096772420050559989617981558627761623516354915042194972780415424737143368453154;
B4[380]<=640'd25674613000958570096700802931751216301790357134310291007938373515764575189841414148789412120042396843558823237677117362163816156707889911361508564264744105057169656942824379190946;
B4[381]<=640'd15525671114281793549346254738296985807362649137031384920716644531009083690640805802440388857211696065884256659483961665678627607700813643130131558231397450446720133159082222783530;
B4[382]<=640'd356155297859651416718751925423078712062146030525341716188525435640458993933687647188768210800945312390178029000756380415375672864808472789712885653889788456587300623585982349354;
B4[383]<=640'd161073899137157954563031808996044099635000851909057003237953476705405038853619578250141141789171829261992745410982416027489033400378928407164599858863910035541676473450621829161;
B4[384]<=640'd45755399207384291697226885512831274120304169603703336419933773257249444236287531838564368265181300408609622937507345967154008780432152346743545720827017959978308717947316600832;
B4[385]<=640'd7187934121633874809555012310468119129438749047398775793377774809054203571410819902738896893029323845651932544670709887171214101148165466586870898445338364829034995204745068544;
B4[386]<=640'd10619801950395256909066038918980435474620628334826615734215839230981345285511122126820276002659401659974549993024114553777670680315425221282018643331660663435622230883926278144;
B4[387]<=640'd28010168083844894103433488966952496366974905400220617105323853692540680125918780961624195653443854910947534641555933426091624117353415644498139193259853096762174622769593974784;
B4[388]<=640'd14979792806826755568901820660736321290645753394993491237280068171655753021143257438031704930896863874552742936502992475235792759086767829982332585525785162449770213366229368832;
B4[389]<=640'd243660616480681350005216378361605409704997255808898302284296474484965187334733395790154484973438968817122154993922930260487637024979593213391292244732140430469217957994429265825624745836544;
B4[390]<=640'd17404329748651702712688522588498579769648240808015136771784476561304629109026339006601591488880300260219345484263980723002983094077564836588071655948931711400587832348775673995372510838784;
B4[391]<=640'd78319483868789332198032752574198361021587936633049335705976063344864888476581846493550668981234861945646124446719147417637555807711601432116827476446615803327247413708261364147755553914880;
B4[392]<=640'd635258035824623637286877603798517909761850687751972578259491425389794173420637410284586510916576219121272954652279477367976634822768330581194046669445763275858610740903231012678335341789184;
B4[393]<=640'd844109992808061480058430770835258613020399203658702521216291742043837072404293137994047921778399040232996248278658117956762793068065002630071326876949272092392737037271733954338335286624256;
B4[394]<=640'd469916903212735257679254749816873215868651322690266189799481024677945325987130695824654046584483169533183407954555383815566811577367968299151838307567108236528362057001973974877320454864896;
B4[395]<=640'd69617318994479298044022656201128736741725230211896620133995751848111058188248758114945407410538197787766761277528085507944464933200050571807383098514572592393106440252229542596219739570176;
B4[396]<=640'd220721504014641988886083180374762156165222098002170998814269314743078757291563796878091811577322217132057609929386313763388835600553335413949107363150744378848377432965120;
B4[397]<=640'd1903598566255293382200036919057058091164267239391201422680031783231609737316406482233074563900120414848116043982332221447192542793798954215823002318960204191732277064263167561118380982272;
B4[398]<=640'd558026322565123116295356311184427176856947384848239952116310202339900416160880333361939057262890710752762611010169861932668075370335046097726283989880336010417080135518850156415214591934464;
B4[399]<=640'd142576269300693600582542494293493291460984429201482179071860519456602524459386366967785710116210709690904910260856818611000406576099509233370095030162382231806151541017947751832882719557156864;
B4[400]<=640'd424402333459955913533284916288401215142230584976900030028078799598264141884851593214187359981336863065889810536712639272843445132709466898394677002215227792637233725440;
B4[401]<=640'd42440164983597486435432820437370815442834064965889408539532523660388297066532997647912429277625891845635413365908371374194338346714889102883232517457356658009681428480;
B4[402]<=640'd16588169970896061554170342722253618393458063359462544251877762923935900676261619264719186508758071560782928860612287534105818304246689719105683888076110814428123889664;
B4[403]<=640'd25751782559965259157620949305923225237653352715466252403264985564897336147781554528274409152818939516526168616500540147744922950883995103580759518503456811681880997888;
B4[404]<=640'd5641665138075400576712865232719079647126934472480331501105229341773013587407635395076145690451642859151092645756063867330166154752906435598671944760926977862787923968;
B4[405]<=640'd7041646271629720889124426574280003411721906262079098827449211521341782216576525618138346342570474701323366567522892085675352856314110137917264461245146194629093228544;
B4[406]<=640'd874192523200916682867405252402651458533648310032937110900937319156462542721691142526848587322942971536565837279072545899588990576951920686482004848750817128176680960;
B4[407]<=640'd73330536624836054247347676855462185459754476615971518604121410640526276349990590856177367678226749209417445733936537402833949634018940009232268495829749770819207168;
B4[408]<=640'd18564149666434562113938406815169093236853328380909744121654010549110522933869953781626002733777698811575132383825772218744295553844676645152629440044106802329026816;
B4[409]<=640'd12379042490951777847601265858002582951771389945724396133510311001345781167085567721137686607927921542519160420228032659187567856577376692638796993243230050078162944;
B4[410]<=640'd3135180553819494241351050825039645524610585609721931814353108874619721074635337964120733344345348206864602186025381906135224563269825746090586817114572505806274560;
B4[411]<=640'd463504367918535729965943733928941932243844360891681286320452855691687794932180762225156410332343781497617660375946243323793918615082697855645821358562730752081920;
B4[412]<=640'd397145706449281543897048924720439474983131802669594706144193051512503729197913192536501482880188146426870757724450594399991794340509879501387576446166777141919744;
B4[413]<=640'd43852327451252088237003379734242931776618460889481424054854330729812303262302198881481916861657695677714914201721553915383945879195835207803696513208893241819136;
B4[414]<=640'd55907768960660915302804513961145021084127783999974341193085515702151138282258992136223749930825636453709259824021759039563435894385796855385987734858430997856256;
B4[415]<=640'd12363996309626570326560370365762275102660266327192654353635667893473055956591874562703977324345808547067425748087191619562707210172107941528303747906006748758016;
B4[416]<=640'd798419944116753091208179236927823763319506707772650681870908465202918974535238068681044293043513218128281301745667792063301707172698213978527465569667690529024;
B4[417]<=640'd1381835658397991530716868442479450531407002497854034463881322867259962470178467937157297362050518550287881249420570425524305309823799906525130177689539313920;
B4[418]<=640'd107678101575644286662839100363707113057811002591100549802782228111270244215553448389681708972173654450891214219261450720118729593153188866153506927519790530816;
B4[419]<=640'd206613901228894105273419785789015488985263780735192617145239391379840346380672011100714538229739736856350929366122138601661872760005425295025580077536946159616;
B4[420]<=640'd6541536991488976400186847861037956801507456286791664726354557847465204727603517053332293534960581316190340880404609268723218570504498662712864535231042945024;
B4[421]<=640'd1033707293458154211399811573280001671495498008505239438264162006797631549601646633854945819594487361207234195666886891217267094101030620909521926614371270656;
B4[422]<=640'd431144822948073351524261989259837253816871148874791605103214237656985366139816277861653003119181160734734476505091580308109928275510714248488389428383842304;
B4[423]<=640'd1538349556524049030095674562518499123302802973746338496002377452424845599270904824659990571374727342922654967087682490057544606947244091614613591978160422912;
B4[424]<=640'd416867470290344719900144920282130657787639294927531399444051579528901259569108676499158157930485432894888009108949346010816887936992449500608565863595902977;
B4[425]<=640'd9086113979867721568978315794758309138193250530417240728025328018539221203551350430515991992100049007633771252893021868140847594981348502669761517040175104;
B4[426]<=640'd1584411362517373355211448929839865629278931812003462763001654423338607154937861273901144598081158854694717635212617193601701059794340949971506135033708544;
B4[427]<=640'd705735293104467845024315246005276154755480649726612508810968775817116877512281696908170770650945800606006927817700822600077066921633407546150773451653376;
B4[428]<=640'd632992905420093488391696057073674337665863625860484181279508457454222652324594642494840470765120815511747578609207952823771949413502564500583897871941632;
B4[429]<=640'd83934954117879133896064008301203933821776360212773139867630383098532842088221994611966582533340017128741701588327095677264727292946573624750457657229312;
B4[430]<=640'd25147004273953452054188129431895132378408273249151284714376823540641199856841134253237047159262868563010452792681446418409774598855167992371260550692208640;
B4[431]<=640'd51966125214084022540735404862830196360201056981843608027424762280877342034392227617867164344315908878006278702038077908864901739228006851690596926832510976;
B4[432]<=640'd3036381208361885243647897015431245357216455620748869932040299440989735905069754448990913168875320561837469102335857726575240352651560852934514817630208;
B4[433]<=640'd247364233366533865124049451887231460567673965231720766012967856336962926651172299317695641833379311739166316168688960265852590991411034843798480879616;
B4[434]<=640'd122278866327216869216761925999438780348091779101130226741790767971330339627791987917755544484135841379279180931104516469901373944040415876402833784832;
B4[435]<=640'd195995092739627383243910230724565328029782914749606874745353792552532288422917031133490532100949804220055689400505493180796362555732561480347400798208;
B4[436]<=640'd49123844334084890695960790352582806007601883646048972146663269590920255576775414743635983088785090355564003550193905419728747893004084768564838400000;
B4[437]<=640'd1873049223969234831052243045423166675104611933156164553660469704644653826066480362568061187512253093877634686206585397596683343546550464929251459072;
B4[438]<=640'd680588794486969309785680747753092004406589204884537491838486221809090606052421464929274234707599275576756803579799764694060878010266455159345250304;
B4[439]<=640'd180963819422539785316272279930177016741161969653533557625927386680883324499578229840992926722624470049582007108677694397713099770394761081674268672;
B4[440]<=640'd45173849098273419819064010086709197755524426379973743178470673138051474065920310815310705980602895026746839560408393011877016027706472473213034496;
B4[441]<=640'd11877651534597851153875389214694375135888760871043919565809155817525368683514974351325554302076626167469757842787452390743573943478772891056660480;
B4[442]<=640'd2771113332077174581249098874252422932309962451926485759564773830405933295592176193304565035908027443529161404387136061460569930430881828654047232;
B4[443]<=640'd3097234850247230520229343324681496462627770925854140844747885127754803971116504246572461008180818200298232443751168488777363852277772286768971776;
B4[444]<=640'd756119928190705558294449717062406880001614412844569614621308552039352365268634655146899567970205778893917035320458355808212445154602438608551936;
B4[445]<=640'd9145748430003394019202953128671782233523571564237815326118948881165595172344475569937999475282145070491794712190949028112317612193124355964928;
B4[446]<=640'd21340077980675728144210141213837833172393450079953920295192280833493609680174058941120235972551347846382391746769520177803697514532899297165312;
B4[447]<=640'd63461376944064480661949369323403322418965060190312881422631351254143936986256081052634967911879700520266560053480071008124928;
B4[448]<=640'd1433169506199070937416054733497569661664514865569756412299956053838075647843372010358393944650382188034705335279365308563873792;
B4[449]<=640'd2778071843986401967350916717854421189544710780419041507505527224793601637089196488975485690897427643449842875519897756692335566849;
B4[450]<=640'd18599470984391163389068285940328043756880855267820277587241357207387271919939562641524247786569635883506894913107680247668539392;
B4[451]<=640'd1439017929896646059452398950779675294703095657031066324495215640232144841608422191827350890944722918646257345631185560537658923417600;
B4[452]<=640'd311927857889967328693739708242717828153496164822539776230951337976737341776194417215413416551913911622203100814308528550926285275136;
B4[453]<=640'd9400738459450477398542128289209592222706647551052575838740088012754275169164351864793151677786016569075908605411464940356482587688960;
B4[454]<=640'd7426942359414614285766222261449348198006648146952036457202922756172553147760572139211857392951045318838254829153260136707560837221888;
B4[455]<=640'd2391432180398305676964493456037456100396876092152634492784201929902039549095263024931679384886522174238605739122828397998500112244480;
B4[456]<=640'd13729595320261219429963804361128136626016483894956128967640935165207170703548405563221930583956121093597052410113861213673215063076346152849620721418717562368;
B4[457]<=640'd11334500417711627463778961997672469119961813084468375877712386177820355410774420222689947042570540497043967254527995937683360072139264;
B4[458]<=640'd536312317197703883982982382583623049984688389610591475692022508150141225478466622454466375062338439064078091465523313672536220314574850456529594877027037952;
B4[459]<=640'd858099707516326236701224406653698534105757209291839660601982489345235113478138337559794251140208422719840896244595969034504741165109260839050446039919114176;
B4[460]<=640'd6757535196691069584129790246589451285612350794134047403199990309197268053764798179475309029467593726881099042636755413954526068319295398208857009640598672064;
B4[461]<=640'd12442445758986730842407141960599417272958798606126448022554490798068002516538317020585699956519557139898265203840651706232186133821619796984025097765025226496;
B4[462]<=640'd1429991446876967046611433097146182140594935629902213563743851357944953209238949570556940984065381821905529688766781485123823522678141743206116490523018824341068680272992;
B4[463]<=640'd3767512106834170683423211829750186426898005779007262223366524783820091324601432129542731642672144943395230949276041414049930628688961248761807174206377677862747504509584;
B4[464]<=640'd427728807902080801748452825641764221519091987796597189874803206302014582816771739410963642734008366221365172690046042217531733475776849780005627508506580592377352761683361489482193011269833696;
B4[465]<=640'd552761513065136683925810526204851591910947958605238587801160958827241904629124987990715020282797967238416713461604677812745956957976974994446819234712351852278903779322935918158412199705318368;
B4[466]<=640'd3119691298780600189870494525170057932126291226929289155832061376527495322757157203763185751934906605758242924782601731742307902891254514605917572623785483217045979776393594826209316470033682432;
B4[467]<=640'd499604746595324742223732088454207106886962087233581110045829594448672536538384925547882757175563843118951130836861993805424623752972205667200380829880322665843964401429365688709144189599875072;
B4[468]<=640'd251728610060641460560311669037765595234810362373347436714564658970879996997015811944045795309439635976774250720619798288949568235681750782475780457974693755433853892801204207046510679223702272;
B4[469]<=640'd134778719551359281508278224155318655921461662574807524470097534259388715891165575928335544048077580121354104721151303254400829052646815096943795072481914680491062049002155512969565770182820352;
B4[470]<=640'd258967724508091625482031910153045640993760182866477665051351425011565601745372083280301843129339073345344199655520754505798531081622586684785750230046974242172015457404657111978758811780419072;
B4[471]<=640'd657170087786786812527778355030881350252997541237916660397617118076379587397056929039258466002586428027253408452029102909242861074543740440520021884788184777727548971011854483730912543438705536;
B4[472]<=640'd3220690656873082106607826585446616407160777542272079545636067879246165274019684162376751201016145281168784127100947868412037453984187563081516671518567378982279292212664386784548915686644613520;
B4[473]<=640'd4442159292452226240828013477563585478780755024068117988037138892701991256915007504095369484443538678700357862438289877688977849789637905790320276925346256833716827684234439859455491016329569158;
B4[474]<=640'd1207371207062020936108193944298796276402676368087080111628308573040768839790704217862684426654423441432801764935321533849585413930020123473382526853826689860579595583071208764435817498678919298;
B4[475]<=640'd4219368644564264591799258215819450675317301044808556321845936219055705936666675431726524391185241520450206537956785283824720208323369647800764002975770177679103091182129013844497325782150024831;
B4[476]<=640'd214351588938240199285597267214695884665063971084871378892177485006383556632631127587531159194017753602435695305951462278915782882209126137983120336500703837586903133901212860717709018831887871;
B4[477]<=640'd1978314381191351639665156243797796629024807476116115287024189872683404155378422132394526867859635532699438351078000717667595952270402310191310173967704847039149531236979106719535257549912539614;
B4[478]<=640'd1942598322963964503080436861769047984926347773075976468184944368058717675575886546457988066070492255913611486575721400641047970889910987473052665440229542151559342909204591076244387032989664875;
B4[479]<=640'd1710637158363456532459975082879842637784614442408524722711639649430191046664744387319151112925410394847596649358565025718024967580878589415898609211745877122423444093871854506163567398893159018;
end

//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)   pixel_data <= 12'd0;
    else begin
        pixel_data <= {R1[pixel_y][pixel_x], R2[pixel_y][pixel_x], R3[pixel_y][pixel_x], R4[pixel_y][pixel_x],
                       G1[pixel_y][pixel_x], G2[pixel_y][pixel_x], G3[pixel_y][pixel_x], G4[pixel_y][pixel_x],
                       B1[pixel_y][pixel_x], B2[pixel_y][pixel_x], B3[pixel_y][pixel_x], B4[pixel_y][pixel_x]};
    end
    
end  
endmodule


// The whole VGA 
module VGA_out_color(
    input sys_clk,
    input sys_rst_n,
    input [1:0] choise,
    //VGA
    output vga_hs,
    output vga_vs,
    output [11:0] vga_rgb);

//Wire define
wire vga_clk_w;
wire [11:0] pixel_data;
wire [9:0] pixel_x;
wire [9:0] pixel_y;

//****************************Main Code**************************
// 这样的话每个VGA输出都有个时钟分频
//优化的时候可以将时钟分频拿出来
clockDiv clkdiv1(
     .sys_clk(sys_clk),         
     .sys_rst_n(sys_rst_n),
     .clk_25M(vga_clk_w));

vga_driver_color VGAdriver1(
    .vga_clk(vga_clk_w),   
    .sys_rst_n(sys_rst_n),
  
    .vga_hs(vga_hs),      // 行同步
    .vga_vs(vga_vs),      // 场同步
    .vga_rgb(vga_rgb),      //4+4+4
    
    .pixel_data(pixel_data),    //像素点RGB data
    .pixel_x(pixel_x),       //像素点横坐标
    .pixel_y(pixel_y)        //像素点纵坐标
);
 
vga_display_color vgadisplay1(
    .vga_clk(vga_clk_w),
    .sys_rst_n(sys_rst_n),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .choise(choise),
    .pixel_data(pixel_data));

endmodule