`timescale 1ns / 1ps


// VGA Driver
module vga_driver(
    input vga_clk,      // VGA驱动时钟
    input sys_rst_n,    // 复位信号
    //VGA
    output vga_hs,      // 行同步
    output vga_vs,      // 场同步
    output [11:0] vga_rgb, //4+4+4
    
    input [11:0] pixel_data,    //像素点RGB data
    output [9:0] pixel_x,       //像素点横坐标
    output [9:0] pixel_y        //像素点纵坐标
);

// some parameters for sure in the reference Table 
parameter H_SYNC = 10'd96;
parameter H_BACK = 10'd48;
parameter H_DISP = 10'd640;
parameter H_FRONT = 10'd16;
parameter H_TOTAL = 10'd800;

parameter V_SYNC = 10'd2;
parameter V_BACK = 10'd33;
parameter V_DISP = 10'd480;
parameter V_FRONT = 10'd10;
parameter V_TOTAL = 10'd525;

// counters for H and V
reg [9:0] cnt_h;
reg [9:0] cnt_v;

wire vga_en; // 使能控制rgb数据输出
wire data_req;

//*******************************Main Code************************************
//VGA 行场同步信号
assign vga_hs = (cnt_h <= H_SYNC - 1'b1) ? 1'b0 : 1'b1;
assign vga_vs = (cnt_v <= V_SYNC - 1'b1) ? 1'b0 : 1'b1;

// 使能使RGB输出 // 范围内输出
assign vga_en = (((cnt_h >= H_SYNC + H_BACK) && (cnt_h < H_SYNC + H_BACK +H_DISP))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;

//在范围内RGB赋值
assign vga_rgb = vga_en ? pixel_data : 12'b0;

// 请求像素点颜色数据输入
assign data_req = (((cnt_h >= H_SYNC + H_BACK -1'b1) && (cnt_h < H_SYNC + H_BACK +H_DISP -1'b1))
                &&((cnt_v >= V_SYNC + V_BACK) && (cnt_v < V_SYNC + V_BACK + V_DISP)))
                ? 1'b1 : 1'b0;
// 像素点坐标
assign pixel_x = data_req ? (cnt_h - (H_SYNC + H_BACK -1'b1)) : 10'd0;
assign pixel_y = data_req ? (cnt_v - (V_SYNC + V_BACK -1'b1)) : 10'd0;

// H counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_h <= 10'd0;
    else begin
        if(cnt_h < H_TOTAL - 1'b1)  cnt_h <= cnt_h + 1'b1;
        else cnt_h <= 10'd0;
    end
end
// V counter
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)  cnt_v <= 10'd0;
    else if(cnt_h == H_TOTAL - 1'b1) begin
        if(cnt_v < V_TOTAL - 1'b1)  cnt_v <= cnt_v + 1'b1;
        else cnt_v <= 10'd0;
    end
end
endmodule 


module vga_display(
    input vga_clk,
    input sys_rst_n,
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input [1:0] choise,
    output reg [11:0] pixel_data);

parameter H_DISP = 10'd640;
parameter V_DISP = 10'd480;

// some frequently-used colors define
localparam WHITE = 12'b1111_1111_1111;
localparam BLACK = 12'b0000_0000_0000;
localparam RED = 12'b1111_0000_0000;
localparam GREEN = 12'b0000_1111_0000;
localparam BLUE = 12'b0000_00000_1111;

reg [0:639] R0 [479:0];
reg [0:639] R1 [479:0];
reg [0:639] R2 [479:0];
reg [0:639] R3 [479:0];
reg [0:639] G0 [479:0];
reg [0:639] G1 [479:0];
reg [0:639] G2 [479:0];
reg [0:639] G3 [479:0];
reg [0:639] B0 [479:0];
reg [0:639] B1 [479:0];
reg [0:639] B2 [479:0];
reg [0:639] B3 [479:0];

always @(posedge vga_clk) begin
B0[0] <= 640'h0
B0[1] <= 640'h0
B0[2] <= 640'h0
B0[3] <= 640'h0
B0[4] <= 640'h0
B0[5] <= 640'h0
B0[6] <= 640'h0
B0[7] <= 640'h0
B0[8] <= 640'h0
B0[9] <= 640'h0
B0[10] <= 640'h0
B0[11] <= 640'h0
B0[12] <= 640'h0
B0[13] <= 640'h0
B0[14] <= 640'h0
B0[15] <= 640'h0
B0[16] <= 640'h0
B0[17] <= 640'h0
B0[18] <= 640'h0
B0[19] <= 640'h0
B0[20] <= 640'h0
B0[21] <= 640'h0
B0[22] <= 640'h0
B0[23] <= 640'h0
B0[24] <= 640'h0
B0[25] <= 640'h0
B0[26] <= 640'h0
B0[27] <= 640'h0
B0[28] <= 640'h0
B0[29] <= 640'h0
B0[30] <= 640'h0
B0[31] <= 640'h0
B0[32] <= 640'h1840000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[33] <= 640'h0
B0[34] <= 640'hc000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[35] <= 640'h800000000000000003600000c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[36] <= 640'h80000000000000000060000004000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[37] <= 640'h1800000000000000001c0080000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[38] <= 640'hfc00000000000000001e990000c0400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[39] <= 640'he700000000000000001f99100104000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[40] <= 640'hc400040000000000007fe644c066100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[41] <= 640'hc400000000000000807f6744f8f6700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[42] <= 640'hc40000000000016080ffff63fcf9800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[43] <= 640'hc40000000000010007ffff63cf99040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[44] <= 640'hc400000000c0000003fffff33f99d80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[45] <= 640'hc400000040000019e3ffffff7cfffc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[46] <= 640'hc400000077010099f3ffffdffcff7f8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[47] <= 640'h3c001993fffffdfc37ff1c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[48] <= 640'h3b0173077fffffff7bff0080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[49] <= 640'h800000003fc078c1efffffffffff0090000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[50] <= 640'h80810000000f00f8e0effffffffffec000000000000000000000000000000000000000000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[51] <= 640'hc1980000000e06c70f7fffffbfffff6100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[52] <= 640'hc118000000ce06ce0f7fffffffffff7142000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[53] <= 640'hc018000000ecc63e1ffffffffffffffcc0000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[54] <= 640'h8000000030667e3cffffffffffffced0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[55] <= 640'h10810000003067e31f7fffffff7ffeceb8009800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[56] <= 640'h3c87200000c091ff9fffffff3fffff796000010000000000000000000000000000000000c020000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[57] <= 640'hc31c0000000091ffdffffffffffffffc76000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[58] <= 640'hc3180000000067fefffffffcffffffdf7e008000000000000000000000000000000000180000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[59] <= 640'hc3308000000067fe7ffffffffffffffffe180800000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[60] <= 640'hffe08000000067ff67fffffffefffff8ff981800000000000000000000000000000000012000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[61] <= 640'h7ec38000000002ffe7ffffffffffffffffe01800100000000000000000000000000000182000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[62] <= 640'hffc30000000011feeffffffffffffffffd668c88000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[63] <= 640'he30000000000183effffffffffffffffff67ce8c810000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[64] <= 640'h200100000000803fffffffffe7fffffffffffe1110000000000000000000000000000000b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[65] <= 640'h3f0ffffffffffffffffffffff9000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[66] <= 640'h1bffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[67] <= 640'h119fffffffffffffffffffffff9000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[68] <= 640'h897fffffffffffffffffffffd8c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[69] <= 640'h100000000003889ffffffffffffffffffffffddc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[70] <= 640'h3089ffffffffffffffffffffffdd000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[71] <= 640'h100000000c18dffffffffffffffffffffff89000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[72] <= 640'h2008000000000f3fffffffffffffffffefff9f10c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[73] <= 640'h33f3fffffffffffffffdffffffc800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[74] <= 640'h833fffffffffffffffffffffffec800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[75] <= 640'h7e3fffffffffffffffffffffefc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[76] <= 640'h3fe7ffffffffffffffff3ffffef8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[77] <= 640'h800000003e3ffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[78] <= 640'h1f3ffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[79] <= 640'h7ffffffffffffffffff7fffffc80c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[80] <= 640'h80000008c37fffffffffffffffffffffffb9380080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[81] <= 640'hff7fffffffffffffffffffffffbf90000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[82] <= 640'h3fe7ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[83] <= 640'h3fffffffffffffffffff7ffffffeff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[84] <= 640'h8037ffffffffffffffffffffffffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[85] <= 640'h8c3fffffffffffffffffffffffffffff040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[86] <= 640'hc3ff3ffffffffffffffffffffffffff9e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[87] <= 640'h401ff7fffffffffffffffffffffffffffffe0800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[88] <= 640'h8000000033407effffffffffffffffffffffffff710100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000
B0[89] <= 640'h234c7ffffffffffffffffffffffffffffb80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[90] <= 640'h16dffffffffffffffffffffffffffffff00000000000000000000000000000000000080000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[91] <= 640'h1017dfffffffffffffffffffffffffffffe00000000000000000000000000000000000c60000000000000000000000000000000000000000000000000000001000000000000000000000000
B0[92] <= 640'h11f4187ffffffffffffffffffffffffff9c80000000000000000000000000000000008e00000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[93] <= 640'h81f410ffffffffffffffffffffffffffb0800000000000000000000000000000000008600000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[94] <= 640'h1e483ffffffffffffffffffffffffff90000000000000000000000000000000000001fc0000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[95] <= 640'h40000000010c481f7ffffffffffffffffffffffffb8000000000000000000000000000000000001f80800000000000000000000000000000000000000000000000000004100000000000000000000000
B0[96] <= 640'h180000019300103ffffffffffffffffffffffffffc0000000000000000000000000000000000024e0000000000000000000000000000000000000000000000000000008ce0008000000000000000000
B0[97] <= 640'h8100000ffffffffffffffffffffffffff4000000000000000000000000000000000001fe080000000000000000000000000000000000000000000000000000ff70000000000000000000000
B0[98] <= 640'h300c7fffffffffffffffffffffffee0000000000000000000000000000000000013ee0c0000000000e00000000000000000000000000000000000000000f738000000000000000000000
B0[99] <= 640'h6600100cffffffffffffffffffffffffe000000000000000000000000000000000000020e0f810000000ff8f000000000000000000000000000000000000010f7fc002000000000000000000
B0[100] <= 640'h60060004fffffffffffffffffffffffef000000000000000000000000000000000000007f83c10000003ffcffc0000000000000000000000000000000000000fffc206800000000000000000
B0[101] <= 640'h40060081ffffffffffffffffffffffff3000000000000000000000000000000000000067f8ef10180007fffff80000000000000000000000000000000000003fffc78e800000000000000000
B0[102] <= 640'h10060185ffffffffffffffffffffffff00000000000000000000000000000000000000e6f9ff123c003ffffff0000000000000000000000000000000000002ffffff9f800000000000000000
B0[103] <= 640'h3904710cfffffffffffffffffffffffb000000000000000000000000000000000000200699fc1fff663ffffffb00000000000000000000000000000000000fffffff9b800000000000000000
B0[104] <= 640'h668f7fffffffffffffffffffffe600000000000000000000000000010e000000183e9cfffe7f937fffffff0000000000000000000000000000000000ff7fffff0f300000000000000000
B0[105] <= 640'h3800076df7fffffffffffffffffffffe60000000000000000000000000000f80000001800f8fffeffbeffffffff8000000000000000000000000000000003ffffffff0e000000000000000000
B0[106] <= 640'h800019dfffffffffffffffffffffffe000000000000000000000000080203b0000008023f9ffffffbeffffffffc0000000000000000000000000000001fffffffefea0000000000000000000
B0[107] <= 640'h380019fffffffffffffffffffffffff0000000000000000000000000813f3f8000008033ffffffffbfffffffffc0000000000000000000000000000003ffffffff3c30000000000000000000
B0[108] <= 640'h101180091fffffffffffffffffffffffff80000000000000000000000021f7fffe0800cce3fffffffffbfffffffffe000000000000000000000000000008fffffffff0030000000000000000000
B0[109] <= 640'h1318000f3fffffffffffffffffffffffff80000000000000000000000033ffffff0820eff7ffffffffffffffffffff000000000000000000000000000049fffffffff3800000000000000000000
B0[110] <= 640'he1007f7ffffffffffffffffffffffff8000000000000000000000000fffffff1befefefffffffffffffffffffff00000000000000000000000000001fffffffbff0000000000000000000000
B0[111] <= 640'h3fc007fffffffffffffffffffffffffd8010000000000000000000032fffffffffefbfeffffffffffbffffffffff800000000000000000008000002417ffffffbfe0000000000000000000000
B0[112] <= 640'h8f66003fffeffffffffffffffffffffffc060000000000000000000083fffffffffffffffffffffffedffffffffffc00000000000000000004000100017ffffffeffe000000000000000000000
B0[113] <= 640'h3ee003ffff7fffffffffffffffffffffe82000000000000000000009ffffffffffffffffffffffffffffffffffff80000000000000000000000c901037ffffffefc0000000000000000000000
B0[114] <= 640'h31cc00fffffbfffffffffffffffffffffe83000000000000000000009ffffffffffffffffffffffffffffffffffff80000000000000000004000cc83c7ffffffe00c0000000000000000000000
B0[115] <= 640'h339c00fffff9ffffffffffcbffffffffff830000000000000000000017fffffffffffffffffffffffffffffffffff8000000000000000000001fecfc8fffffffe0040000000000000000000000
B0[116] <= 640'he000000778007ffffbffffffffffc3ffffffffff90c000000000000000000003fffffffffffffffffffffffffffffffffffc000000000000000000000f7ffc0fffffffc0000000000000000000000000
B0[117] <= 640'h810000cff1007fffffffffffffff1cffffffffff90c0000000000000000000b3fffffffffffffffffffffffffffffffffffe000000000000000000013fffe79fffffffc0000000000000000000000000
B0[118] <= 640'h30000fff9007fffffffffffffee047ffffffffff34000000000000000000087fffffffffffffffffffffffffffffffffffe000000000000000000103fffeffffffffed0000000000000000000000000
B0[119] <= 640'h306027fff800ffffffffffffff9e0106fffffffff6440000000000000000008effffffffffffffffffffffffffffffffffffc700000000000000000003effefffffffff0000000000000000000000000
B0[120] <= 640'h30103fffd807fffffffffffff8f811fffffffffff3f00000000000000000077fffffffffffffffffffffffffffffffffffd8d00000000000000000000397fffffffffc0000000000000000000000000
B0[121] <= 640'he300c1ffff007fffffffffffffdf1c0cffffe8ffffff80000000000000000007fffffffffffffffffffffffffffffffffffffd0000000000000000000001ff7ffffffcc0000000000000000000000000
B0[122] <= 640'he1f0c3ffff006feff3fefffffffffc0fffff40207fff80000000000000000007fffffffffffffffffffffffffffffffffffffc0000000000000000000001fc3ffffffc00000000000000000000000000
B0[123] <= 640'h39ff3ffffe002ffff3dffffffffffffffffe04000300000000000000000000c7fffffffffffffffffffffffffffffffffffffc80000000000000000000000cfffffffc00000000000000000000000000
B0[124] <= 640'h7ffffcfffe00367f88e3ffffffe3fff0ffdf40000000000000000000000000ffffffffffffffffffffffffffffffffffffffe9800000000000000000000004e7fffffc00000000000000000000000000
B0[125] <= 640'hffffffffff00007f8c3ff7ffffff7fffffef800000000000000000000000003fffffffffffffffffffffffffffffffffffffef0300000000000000000000000ffffffc00000000000000000000000000
B0[126] <= 640'hffffffffff0003cf803ce3fffffffeff4ffe8980000000000000000000000006ffffffffffffffffffffffffffffffffffffff1fc80000000000000000000003ffff7000000000000000000000000000
B0[127] <= 640'hfffffefffe000180c10cfffef9700701c77e88c00000000000000000000000041fffffffffffffffffffffffffffffffffffff7fdc0000000000000000000003fffdc000000000000000000000000000
B0[128] <= 640'hfffffffffee002a10020009ffc800804231f06000000000000000000000000000fffffffffffffffffffffffffffffffffffffffff80000000000000000000017ff0c000000000000000000000000000
B0[129] <= 640'hffffffffffc00200000081fffc000800029e0e000000000000000000000000000fffffffffffffffffffffffffffffffffffffffff80000000000000000000017ff00000000000000000000000000000
B0[130] <= 640'hfffffffffe9802040007c07fde000160860e01800000000000000000000000009fffffffffffffffffffffffffffffffffffffffffc4400000000000000000007f000000000000000000000000000000
B0[131] <= 640'hfffffffffe9000060007cc7b8f0003efccc600008000000000000000000000089fffffffffffffffffffffffffffffffffffffffffe4f0000000000000000000ff000000000000000000000000000000
B0[132] <= 640'hffffffffff8000631031fc3f800067fffff6810000000000000000000000000c1fffffffffffffffffffffffffffffffffffffffffffff80000000000000000038800000000000000000000000000000
B0[133] <= 640'hffffffffff8000633f30ff1f20006fffff7e013800000000000000000000000cffffffffffffffffffffffffffffffffffffffffffffffc0000000000000000000000000000000000000000000000000
B0[134] <= 640'hffffffffff60029bff3061df01000fffffff06ff8000000000000000000000cfffffffffffffffffffffffffffffffffffffffffffffffffc80000000000000000000000000000000000000000000000
B0[135] <= 640'hffffffffff700099ff8030ff00000fffffff7effe380000000000000000000effffffffffffffffffffffffffffffffffffffffffffffffffc0000000000000000000000000000000000000000000000
B0[136] <= 640'hffffffffffd903dfeee67cc7800007ffffff7fffffc0000000000000000003fffffffffffffffffffffffffffffffffffffffffffffffffffe0000000000000000000000000000000000000000000000
B0[137] <= 640'hfffffffffff8003ffee7f83e8000e7ffffffffffffc00000000000000000003fffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000000
B0[138] <= 640'hfffffffffff93e7f7ffff37c260003fffffffffffff8000000000000000001ffffffffffffffffffffffffffffffffffffffffffffffffffffff0c000000000000000000000000000000000000000000
B0[139] <= 640'hffffffffffffffffffff7fff660013ffffffffffffe8000000000000000001ffffffffffffffffffffffffffffffffffffffffffffffffffffffcc000000000000000000000000000000000000000000
B0[140] <= 640'hfffffffffffd7fffffff7fff6600f9ffffffffffffe9180000000000000009fffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000
B0[141] <= 640'hffffffffffffffffffffffffe40013fffffffffffffc00000000000000000cfffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000000000000000000000000000000000
B0[142] <= 640'hfffffffffffffffffffffefffc8007fffffffffffff960000000000000000cfffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000000000000000000000000000000000
B0[143] <= 640'hfffffffffffeffffffffffffffc0e6fffffffffffff96040000000000000017fffffffffffffffffffffffffffffffffffffffffffffffffffffe7000000000000000000000000000000000000000000
B0[144] <= 640'hfffffffffffffffffffffffffffffdfffffffffffefbd97c80000000000000fffffffffffffffffffffffffdbfffffffffffffffffffffffffffff000000000000000000000000000000000000000000
B0[145] <= 640'hffffffffffffffffffffffffffffff7fffffffffff7fffff800000000000003ffffffffffffffffeffffffffffffffffffffffffffffffffdffff0000000000000000000000000000000000000000000
B0[146] <= 640'hfffffffffffffffffffffffffffeff7fffffffffffffffffd00000000000003fffffffffffffffffffffffffe7fffffffffffffffffffffffffff0000000000000000000000000000000000000000000
B0[147] <= 640'hfffffffffffffffffffffffffffeffffffffffffffffffff980000000000007fffff7fffffffff3ffec36e7f47ffffffffffffffffffffffbffe80000000000000000000000000000000000000000000
B0[148] <= 640'hfffffffffffffffffffffffffffff7fffffffffffffffffe08000000000002ffffff60fffffffff001ee067deeffffffffffffffffffffff337c1f000000000000000000000000000000000000000000
B0[149] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffe00000000000012ffffff203cfffffff000000648fefffffffffff7fffffffffc001c0f000000000000000000000000000000000000000000
B0[150] <= 640'hfffffffffffffffffffffffffffffefffffffffffffffffec0000001000032fffefa1b3fffffffa0000000000f737effdffff277fffffffe00000600000000000000000000000000e6f0000000000000
B0[151] <= 640'hfffffffffffffffffffffffffffffeffffffffffffffffee1c0000008000367efff79be7ffffffb0000000010170e40f39fff666ffffffffc0000000000000000000000000000033c6fe800000000000
B0[152] <= 640'hffffffffffffffeffeffffffffffffffffffffffffffff7b2100000000003effff7c927ffffffef00000000018f81c00ff37c4703fffffff800000000000000000000000000000fffefe800000000000
B0[153] <= 640'hffffffffffffffeffffffffffffffffffffffffffffffff001000000000007f9ffff837fffffff800000000018f00120f0bf020fc13fffffc00000000000000000000000000000fffefe000000000000
B0[154] <= 640'hfeffffffffffffefffe7fffffffffffffffffffffffffff803000000000003f8ffff83ffffffff8000000000000001000096018c997ffe3ffe6000000000000000000000000001ffffff000000000000
B0[155] <= 640'hf77ffffffffffffdfffffffffffffffffffffffffffffffc00000000000003f9fefe97ffffffff8000000000812100000002008c1dc3ff03fff000000000000000000000000001bfffff200000000000
B0[156] <= 640'he73ffffffffffffdfcfffffffffffffffffffffffffffffe84000000000000013fffbffffffffd8000000000877bf0000000800e1803ffe1feffa0000000000000000000000000bfff7e000000000000
B0[157] <= 640'hf67efffffffffffc7c3ffffeffffffffffffffffffffffff84000000000000801ff3bfff7ffffc80000000017efffe0000000000801bfffc3e9fe0000000000000000000000000ffff7e000000000000
B0[158] <= 640'h64d8fffffffffffc0003fffefffffffffffffffffffffff98c8000000000008000c3bfff3efffc80000000017fffff8000000000020cfef8ff9fc00000000000000000000000017ffffe800000000000
B0[159] <= 640'he70f7ffffffffffc0003ffe77efffffffffffffffffffffd1e80000100000080010cb3e78c8bf8800000001bfffffff80000000020007ec1c289e00000000000000000000000037ffffe800000000000
B0[160] <= 640'hf307bfdffffffffc0001ffffff7fffffffffffffffffffff7002000000000000001f0747c000e00000000037ffffffc03000000110003f00303ce7010000000000000000000027ffffff000000000000
B0[161] <= 640'h7807bffffefffffc00007fffffffffffffffffffffffffffff80000000800000000218c60000e00000000007ffffffc0c000000001003f200103fe680000000000000000000007ffffffc00000000000
B0[162] <= 640'h3847b3fffefffffc00003ffffffffffffffffffffffffffffe0000000000000000000006000080000000000fffffffc08000000080003e000707fef80000000000000000000007ffffff600000000000
B0[163] <= 640'h91e493ffeffffffe00001eff9ffffffffffffffffffffffffc0200000000000000000000000000000000000ffffffe000c0000068000fec10c1ffffc84000000000000000000037fffff700000000000
B0[164] <= 640'h817c02ffffffffff00001fff9fffffffffffffffffffffffff92800001000000000000200000000000000003fffffe10000000040001b780103ff7fc0600000000000000000003ffffff700000000000
B0[165] <= 640'h987e327f7effffff800067ffffffffffffffffffffffffffffb60000c0800000000000200000000000000001b3cffef000000000001ff37ce1ffffee000000000000000000000bffffffe00000000000
B0[166] <= 640'h1c6e027ffeffffd8800071ff7fffffffffffffffffffffffffff0000808200000000000000000000000000009007fe400000000082fffffcc7ffffef000000000000000000061befffffc40000000000
B0[167] <= 640'h9d4002e3e77ffff800007bff67fffffffffffffffffffffffffe0000190600000000000400000000000000001001e600000000001effffffde3fffefe2000000000000000000f9ffffff3c0000000000
B0[168] <= 640'h6390003fff9bcff80000009f3ffffffffffffffffffffffffffe00003300000000001000000000000000000000000000000000119fffffffdf7ffffe6000000000000000000009fffffffe0000000000
B0[169] <= 640'h7c02003fff01f7f1000003dcf9ffffffffffffffffffffffffff8000003f00000080020000800000000000000000000000000011ffffffffffffffffe000000000000000000009fffffff80000000000
B0[170] <= 640'h5c320033e1077121000003ddfdfffffffffffffffffffffffff90000101f80000000020000000000000000000000000000000003fffffffffffffffff480000000000000000000fffffff80000000000
B0[171] <= 640'h88f00011e10671000000000f1ffffffbfffffffffffffffffff8000010030000000002000000000000000000000000000000003fffffffffffffffffffa0000000000000000000ffffffff0000000000
B0[172] <= 640'h89b0000dfc00000000000001cbfffffffffffffffffffffffffc000002030000000026000100000000000000000000000000003fffffffffffffffffffa1000000000000000000ffffffff0000000000
B0[173] <= 640'hd02009cfc00008000000001c3fffffffffffffffffffffffff800000203c000000006c00000000000000000000000000000007ffffffffffffffffffff30000000000000000027fffffff8000000000
B0[174] <= 640'h7d86008ffc000080000000018fffffffffffffffffffffffffe000008213e000000003e04000000000000000000000000000007ffffffffffffffffffffb0000000000000000003ffffffc8000000000
B0[175] <= 640'h659e0081cc000000000000039c7ffbffffffffffffffffffffe0000080100001061018800000000000000000000000000000066ffffffffffffffffffffb0000000000000000000fffdff80000000000
B0[176] <= 640'h68c0080c9000000000000008ce3ffffffffffffffffffffffe0000080008000000006000000000000000000000000000000003ffffffffffffffffffffe00000000000000007800fffff80000000000
B0[177] <= 640'h4086038098000000000000008c33fffffffffffffffffffffff0000000120000000000e0000000000000000000000000000000fffffffffffffffffffffe00000000000000000001ffed300000000000
B0[178] <= 640'he2c7c3111800000000000000183bfffffffffffffffffffffff0000000140000001000000000000000000000000000000000001fffffffffffffffffffff00000000000000000003fffd300000000000
B0[179] <= 640'h677ffe31d80000000000000000386fffffffffffffffffffffc00000001200000001000000000000000000000000000000000007ffffffffffffffffffff00000000000000000003ffed000000000000
B0[180] <= 640'h7e7f7f70980000000000000001010e1ffffffffff9ffffffffc000000013000000010000000000000000000000000000000000033fffffffffffffffffffc0000000000000000007ff40000000000000
B0[181] <= 640'h7eff87601c000000000000000101e40ffffffffff97fffffff8000000003000104200000000000000000000000000000000000021fbfffffffffffffffffc0c0000000040000003fffe9000000000000
B0[182] <= 640'h3effef6618000000000000000001648fffffffffff6fffffffc0000000020001002001000000000000000000000000000000000093bfffffffffffffffffc000060189ff0000001ffefd000000000000
B0[183] <= 640'h7cffc46c3000000000000000001040ffffffffffee9ffffffc00000008400002000010000000000000000000000000000000000829fffffff7fffffffffc0007efe9fff30600003fe40000000000000
B0[184] <= 640'h1ffeff79390000000000000000060803fffffffffb07fffffd060000003080c0108000000000000000000000000000000000000001e3ff7ffffffffffeffc07cfffffffecfc3003f6789000000000000
B0[185] <= 640'hffffffe3f90000000000000000001007fffffffffa071c67ff848000023f8007010000000000000000000000000000000000000000e0fee7ffcffffffffc806dfffffffffeee003f6618000000000000
B0[186] <= 640'hffffffe3ff0000000000000000000013fffffffff0001c7fffb00000061f0001013000400000000000000000000000000000000000787ee1838ffffffffc004fffffffffffffc003e020000000000000
B0[187] <= 640'hffffff7eff0000000000000000000031fffffffff0000006ff90000006feb00000200160000000000000000000000000000000000001001901ffffffff00006ffffffffffffff8076402000000000000
B0[188] <= 640'hffffff7eff0000000000000000000001ffffffffb00000006f90000007ff308300010100000000000000000000000000000000000000c0190000fffffe00007ffffffffffffffcc40402000000000000
B0[189] <= 640'hffffffffffc000000000000000000001ffffffffb00000076f8000001fff18860000000410000000000000000000000000000000000080000700fffffcc0007ffffffffffffffffc4620000000000000
B0[190] <= 640'hffffffffffc000000000000000000000ffffffff208000006f8000001f3f19f8000000001800000000000000000000000000000000000000c300f9fffe00007fffffffffffffffccc618000000000000
B0[191] <= 640'hffffffffffc0000000000000000000009fffffff0000000c6ea20004dffffd3f010800318000000000000000000000000000000000000026c100f9f8e700004fffffffffffffff8ec681000000000000
B0[192] <= 640'hfffffffffff8000000000000000000007efffffe0000000083c080035f7fe33ef803c7dff00000000000000000000000000008000000000006801c012c000037ffffffffffffff77d1f0300000000000
B0[193] <= 640'hfffffffffff0000000000000000000007e3ffffe00000000180000067cffce0f900007c778000000000000000000000000000000000000000000000000000037ffffffffffffffff3fe0010000000000
B0[194] <= 640'hfffffffffffc000000000000000000009c3ffffc000080001800008ec88e8c03100001e37c00000000000000000000000000000000000000000000000000000233ffffffffffffffffe0000000000000
B0[195] <= 640'hfffffffffffe0080000000000000000089ff8ffc0000000000000007c1868c01310119fff800000000000000000000000000200000000000000000000000000003ffffffffffffffff60800000000000
B0[196] <= 640'hfffffffffffe0003c000000000000000897f3c1c0000010000000003cd6080000001197fe000000000000000000000000000200000000000000000000000000000ff7fffffffffdffff8000000000000
B0[197] <= 640'hffffffffffffd813e000000000000000013e388000000000000000604c7000000001193ffc000000000000000240000000000000000000000000000000000000003e0dfffffffffffff8000000000000
B0[198] <= 640'hffffffffffffffbff00000000000000003000080000000000000000048080000000106fffc000000000000000000000000000000000000000000000000000000000009fffffffffffff8000000000000
B0[199] <= 640'hffffffffffffdffff00000000000000020e000000000000000000100c10c008000106effec8000000000000000000000000000000000000000000000000000000000003fffffffffffe0000000000000
B0[200] <= 640'hfffffffffffffffff80000000000000009808000000000000000000304830000000081f3dc20000000000084000000000000000000000000000000000000000000000021dfffffffffe0000000000000
B0[201] <= 640'hfffffffffffffffffc000000000000000100000000000000000000010000000000001cfb8800000000000004000000000000000000000000000000000000000000000000ffffbffffff0000000000000
B0[202] <= 640'hfffffffffffffffffc000000000000000380000000000000000000000000000000011cff000000000000240c80000000000000000000000000000000000000000000000007ffb7ffffc0000000000000
B0[203] <= 640'hfffffffffffffffffe000000000000000cc0000000000000000000000000000000019f7f0000000000017efe80000000000000000000000000000000000000000000000001f082ffff81000000000000
B0[204] <= 640'hffffffffffffffffff000000000000000ec000000000000000000000008000000000897f01040000000127ff8200000000000000000000000000000000000000000000000007020fff80000000000000
B0[205] <= 640'hffffffffffffffffff4000000000000003c0000000000000000000000000000001001cff031e0000000367e783c0000000000000000000000000000000000000000000000000006ccf10000000000000
B0[206] <= 640'hffffffffffffffffff0000000000000003c000000000000880000000000000000063ffff033f800000867f7fffc000000000000000000000000000000000000000000000010000048400000000000000
B0[207] <= 640'hffffffffffffffffff8000000000000003c0000000000000800000000000000000e3ffffe3fb9901011e7effff8800000000000000000000000000000000000000000000000000060000000000000000
B0[208] <= 640'hffffffffffffffffff000000000000000080000000000080000000000000000003ffffffbd6fc20f00fffbffff8000000000000000000000000000000000000000000000000004100300000000000000
B0[209] <= 640'hfffffffffffffffffff000000000000007c00000000000000000000000000003007fffffbfffec0683ffffffffe000000000000000000000000000000000000000000000000000300000000000000000
B0[210] <= 640'hffffffffffffffffffe0000000001cc0018000000000000000000000000c0001007effffc7fffcc787fffffffffc80000400000000000000000000000000000000000000000000000000000000000000
B0[211] <= 640'hfffffffffffffffffffc00000000ffffe300000000000030000000000008008003fffffe67ffffc7c7ffffffffffc0007efff80000000000000000000000000000000000000000000000000000000000
B0[212] <= 640'hfffffffffffffffffffe00000000ffffc70000000000000f000000000000001983fffff867ffdfc7ffffffffffffef01fffffe0000000000000000000000000000000000000000000000000000000000
B0[213] <= 640'hfffffffffffffffffffe80000001ffffc7000000000001cf800000000048001bf8fffffc67ffffcf7ffffffffffffcc3ffffffc000000000000000000000000000000000000000000080000000000000
B0[214] <= 640'hfffffffffffffffffffff4801fe7ffffff000000000003fcf8000000000801f0fcfffffe81fffeff7ffffffffffffff7fffffffe00000000000000000000000000000000000000000000000000000000
B0[215] <= 640'hffffffffffffffffffffffc33fffffffffe00000000007fff800000000000167fffffffe81fff7ffffffffffffffffffffffffffc0000000000000000000000000000000000000000000000000000000
B0[216] <= 640'hfffffffffffffffffffffffb9fffffffff8000000000137fff00000000000079fffffffff0fffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000
B0[217] <= 640'hffffffffffffffffffffffffffffffffffc000000000bfffff000000000001f8fffffffff0fffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000000000000000
B0[218] <= 640'hffffffffffffffffffffffffffffffffffc000000000ffffff800000000081fffffffffff8ffffffffffffffffffffffffffffffff100000000000000000000000000000000000000000000000000000
B0[219] <= 640'hffffffffffffffffffffffffffffffffff00000000037fffffc000000000007ffffffffffc3fffffffffffffffffffffffffffffffb00000000000000000000000000000000000000000000000000000
B0[220] <= 640'hffffffffffffffffffffffffffffffffff80000000037ffffee1f0000001007fffffffff3c1ffffffffffffffffffffffffffffffff20000000000000000000000000000000000000000000000000000
B0[221] <= 640'hffffffffffffffffffffffffffffffffffe000100047ffffff73fc46200003ffffffffff1e3ffffffffffffffffffffffffffffffffe8000000000000000000000000000000000000000000000000000
B0[222] <= 640'hffffffffffffffffffffffffffffffffffc00010007ffffffffeffeef100c7ffffffffffdffffffffffffffffffffffffffffffffffe8000000000000000000000000000000000000000000000000000
B0[223] <= 640'hffffffffffffffffffffffffffffffffff000083007ffffffffeffff23817fffffffffffdfe7fffffffffffffffffffffffffffffffe0000000000000000000000000000000000000000000000000000
B0[224] <= 640'hfffffffffffffffffffffffffffffffffe00000fe7ffffffffffffffa39067fffffeffffff3fffffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000000000000
B0[225] <= 640'hffffffffffffffffffffffffffffffffff00003ffffffffffffffffff7c167fffffffffff8cfffffffffffffffffffffffffffffffffc000000000000000000000000000000000000100000000000000
B0[226] <= 640'hffffffffffffffffffffffffffffffffff0000ffffffffffffffffffffc39fffffffffff9fe7fffffffffffffffffffffffffffffffff000000000000000000000000000000000104000000000000000
B0[227] <= 640'hfffffffffffffffffffffffffffffffffe0003ffffffffffffffffffffff9fffffffffff1ffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000
B0[228] <= 640'hfffffffffffffffffffffffffffffffffe000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000400000000000000000
B0[229] <= 640'hfffffffffffffffffffffffffffffffffe001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000480000000002040000
B0[230] <= 640'hffffffffffffffffffffffffffffffffff80fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000248000000000000000
B0[231] <= 640'hffffffffffffffffffffffffffffffffff81fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000040000000400000
B0[232] <= 640'hffffffffffffffffffffffffffffffffff83fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000000000000000000080000000000010000
B0[233] <= 640'hffffffffffffffffffffffffffffffffffc7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000000000000000000282008001000000008
B0[234] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000000000000000000040040040801000000
B0[235] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000000000000000000808010000800000000
B0[236] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000000000000000000448000000000000000
B0[237] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000044200000000000000
B0[238] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000020048000000008200
B0[239] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000620044101080020808
B0[240] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000226000400000000000
B0[241] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000021104008000000000004
B0[242] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000000000000000090100008000000201200
B0[243] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00080000000000000000000000000000000411000400000000
B0[244] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00100000000000000000000000000000200000002000000000
B0[245] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff100000000000000000000000000041330004001000040200
B0[246] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000004000080000062190004000000040000
B0[247] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff030000000000000004000090000201180000080000000020
B0[248] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000400409000028008000100b120000000
B0[249] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000020011000804602000001980040800
B0[250] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc0000000ffbf82a6040900008208480101013100080548800
B0[251] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000ffffffffff88401441a202000080020100040400000
B0[252] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00003ffffffffffc24d04021002000c00004001000010080
B0[253] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00fffffffffffe80100420010000001001008c02600000
B0[254] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff01fffffffffffe82040482002000101002094602400000
B0[255] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2a0004008001001000044004106440840
B0[256] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa00401088008801001008021090440800
B0[257] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffba40480849000003089103000400010000
B0[258] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffffffffffffff9f7400104410001200001006004002001000
B0[259] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff10ffffffffffffffffc80103400000800019040060600101380
B0[260] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec000fffffffffffffff646015208008000608982440210050000
B0[261] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000ffffffffffffffd322225008491000008910490248088400
B0[262] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef3ffffffffffffffe109347630491090888001068808204008
B0[263] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe9885264204998208284000040009012100
B0[264] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6d03410cb25924188104090102001000000
B0[265] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe539c4cd8b702e088012190905200024000
B0[266] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6cbcb44a1b0d2c0c6a183b01251c0100030
B0[267] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff663cb2528b4c6643218c320320ce0000200
B0[268] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe25e7307091641b22484300380210090400
B0[269] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe61f734200d4d9b64442020094010193810
B0[270] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa79d9302018cca09206a0280c4040104008
B0[271] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4deb8718d3887c0b634ba0319840424200
B0[272] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcce1a298d2900519006192183018124230
B0[273] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb36fc94b019b280c4086320060008049108
B0[274] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb36f031c40b225446a22064826400199906
B0[275] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcf326625848a2c60301192180c0900008900
B0[276] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa7337a8cc8081860761c8202413000828820
B0[277] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3bd3ecce0093008031e40f0032170c23100
B0[278] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddb3344084813821011961fa04805045180c
B0[279] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9ebe2948c2012824dcc9a3c2649209010000
B0[280] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefb607ec404124c22cc64661a604c8432000
B0[281] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe798174d20c8258804c26591098101860e01
B0[282] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff719d63650c0121041a7221c48164f0404800
B0[283] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcd98ce1042961423b03200e648490404400
B0[284] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe96e64f20448141a27c0127c824d309a01220
B0[285] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcf8826782148093309e4ca4c02409b0e25184
B0[286] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7e6993c31c8d35b1b324f205250922604100
B0[287] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee7f349bc2460c676497386613830004001010
B0[288] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff76ece0de246cccb4e969c0723987010000070
B0[289] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff33ec31e61b0048e0e4f962240848881e06400
B0[290] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7a33bb8e4998408e9304da0486844a24310708
B0[291] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcc9bd898364088230a940011010000e11006c
B0[292] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffce74c4c301a4481d641fe080b0230316c03224
B0[293] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2484024cda0413c8b0fc8c321904196003210
B0[294] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd2620f2481e2017989678b070643008b004242
B0[295] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff231c326110219e14c7329840e19d3600818c0
B0[296] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff91061a2811a0801c0e965c198314321782048
B0[297] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbc02189000819040ec09e582f05cc666184b2c
B0[298] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe448000088091904684e403998c1242501914
B0[299] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3ffffffffffed300405a40601291662750331264588401900
B0[300] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbe13fbfff3fefa689018202c0804c02e93020660e1004480180
B0[301] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0213ff7a00baac0702cb008c088482203922104200038784190
B0[302] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00211bf3000000201084b2246189821823882068990071383024
B0[303] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3fff3fffffffffffffffffffffffffffffffffffffffff00211161008000104214099410a804c0212020988b1211981204
B0[304] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1ff807fffffffffffffffffffffffffffffffffffffff8800008917d80009202220014022021e629b2619c233209d82048
B0[305] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc01f8023ffffffffffffffffffffffffffffffffffffdfe300100043fff80012002131c82363214c08116120f89007485802
B0[306] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe003f003fffffffffffffffffffffffffffffffffffffffe3b09014000000000060991080202433110c106169e8856320980a
B0[307] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800ff003fffffffffffffffffffffffffffffffffffffffffe000000000000061080024009040a699912820d9850060709804
B0[308] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe003e0001ffffffffffffffffffffffffffffffffffff0010000108000000003200990023198602209892120e6198840d8c802
B0[309] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7801f00000fffffffffffffffffffffffffffe17fff600001c0f6988e10000007319612182c420008e194518109f78588b86060
B0[310] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3203e040007fffffffffffffffffffffffff00000fffc3fffffff180e400001829014195894c64201d8d83080b2db84984c2031
B0[311] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbf00000007ff9fffffffffffff830ffffffffffffffc187fffff108640eccfc2020006c84c464267e1931281ce0752188c9830
B0[312] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7e00600003ff8fffffff06fd0381ffffffffffffff0000ffffff108c40efff9221e30e486602e627e49560819e825202600800
B0[313] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff03e000008003ff7cfffffffffbfffffffffffff80000ffffff9809b1cfffd88b8045a0c330a027338922c06eccc8013c2086
B0[314] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000007ff9fffffffffffffffffffffffe00009fffffdc8c521dfffcc89d836c01138e326298b38e0c641c9073c00c6
B0[315] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000080181f000f8787fffffffffffffff3ffffffe0003ffffcfe009a31bfffec01c822430088a18d65924cea4e722c23044040
B0[316] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000008380fffffffffffffffbffffffe07ffffffcfe4408113fffd8109248304c48a0c08610e0480467281cd46200
B0[317] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbf8000000000000003ff0ffff1ffffffffffffff7fffffffefe50b2332fffe812c12930662402001039f809c848c622444000
B0[318] <= 640'hf80cffffffffffffffffffffffffffffffffffffffffffffffffffffffff07000000000000000f0071f007ffffffffffff9efc5ffff64809b20261ffe400408e8883306080208bdea94c080511844040
B0[319] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2000000000000000001060003fffffffffff9ffffffff648a4108021fff204206fc2219a089b809316c165002132c40200
B0[320] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7ffff3000000000000000000000000e9ffffffffffffff70f924024101203fff00230150011c2089b1422660111018191901230
B0[321] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0e0fc0000000000000000000000000005ffffffffffffef07904232340213ff900490858444b020918808e7011a1c3085883011
B0[322] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff800f800000000000000000000000000001fffffffffffe784490132244c83ff9e01c261c500986000023092803876d4440c2049
B0[323] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffe07fc000000000000000000000000000007fe707fffffb38408181a4001a124440002402000080004022222812139454e141680
B0[324] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1ffc000000000000000000000000000001ff0effffff9384841c08000601040021001c000a0e6c0c2023248962080024c04810
B0[325] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000000000000000007ffffff9200020008044008040021114f841380048c3e32404148624104842026
B0[326] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000000000000000000000000001fe6800002130248000005802001ac0c14c82480170420c118105906041602
B0[327] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000000000000000000000001006001040001224c89018000a12411a50462344012408808124c802058460c
B0[328] <= 640'he7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1000000000000000000000000000000000000620000011130040271820020002021800312221060020102501911e80808
B0[329] <= 640'hffffffffffffffffe0e0fff810ffffffffffffffffffff7fff0000000000000000000000000000000000000000000000007ffe0900089388200031920040018201a01c1232006440c025251259c82880
B0[330] <= 640'hffffffffffffffffffffffff3e7fffffffffff0b1fc0ffffffffffffffffff00078f6000000000000000000000000000007ffc831000110400002144004291c800111e081202156808216000600062d0
B0[331] <= 640'h7fffffffff7ffffffffffffffffffffffffffffffffffffffffffff0c0000100000000000000000000000000000000000001e6010002089200400100020002060901c9008102010c4838006000005298
B0[332] <= 640'hffffffffffffff0007ff7fff01fffffffffffe00000080c00003ffe000ffffffffffffffff00030000000000000000000000ae000001001108801080020046010084411299a2041008200e7008486220
B0[333] <= 640'hff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff07f800008000000000000000000000200000010001018011000122400058c411904802103401b122125a346400
B0[334] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1ff800000000000000000000000000b0000902012400002100082000120c0840000c20013c00d3001822242210
B0[335] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc081f80000000000000000000001040c00201000c240040004804118880310c0620c00080400c10090c6830
B0[336] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecf1e00000000000000000000480820e040000138000040a0200004c0253884200244988044161801344800
B0[337] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000e000000003800000e001240909000400000040000024200620002490880404c10006080a
B0[338] <= 640'hfffffe1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3c0000000000000006000000801e000208082240900900140004001800100020001082100c018821251
B0[339] <= 640'hffffffcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0c2000000000000000010080124080000920848809000104c28010041000820400861203009002021
B0[340] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fffeff000000000000000000c00000000000000210040010040883010c0130060004829247020842224
B0[341] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0ffffee7ff000000000000000c0000000800882321082020001048101000010000804024810060a42810
B0[342] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0ffffc6000c0001000000000400800000c0082430000004040002000000210100084042080008022080c
B0[343] <= 640'hfffffcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0ffffc600000001fc00000004081000200400a0400040048002000330181088000208208001100021800
B0[344] <= 640'h3ffffe7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff07ffdce000000000000010000006000100400a000100180000300000c000808001008010101000003040
B0[345] <= 640'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3fffffffff0dfffc3a000000000000000000200018200c0c400000092004801280c049100010069604901010000000
B0[346] <= 640'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff03fffffffe0df99ff00000000000000000000010180204088100000000208000404860880018100204080082000020
B0[347] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff201bff1fffd8e0000000000000000000000000000040810810005000008000020000600806010200010000020000004
B0[348] <= 640'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff8861fff80900e07ff98000000000000000000000000000000030c0004004220048460106c20020080000000010000000060800
B0[349] <= 640'h3fffffffffffffffffffffffffffffffffffffffffffffffffffffc0400000ff00180000710000000000000000000000000001000000042402000120048120202015010480800100000800000000020
B0[350] <= 640'h7fffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000180000000000000000000000000000000000000000720012400400000022022082408020800800000000000001028
B0[351] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000000120008008400000400000060100000000c02000000000041008
B0[352] <= 640'hfffffffffffffffffffffffffffffffe7fffffffffffffffffffffc00c00000000000000000000000000000000000000000000000200080001000040031086301011140000120400000000400000800
B0[353] <= 640'hffffffffffffffffffffffffffffffffcfffffffffffe3ffd7feff800000000000000000080000000000000000000000000000000000010080000840408000900019008000005004000000000000800
B0[354] <= 640'hffffffffffffffcfffffffffffffffffffffcfffffffc0fffff800000000000004000000000000804000000000000000000000012000001008008000048201800004820000000802000000000000000
B0[355] <= 640'hffffffffffffffc03bfffe07fffffffffffffff13c0fc000ff0800000000000418080000000000000010000000000000000000000200000080024000000000200002000010000241000000000000000
B0[356] <= 640'hffffffffffffffffbfff007fffff8001ffffffff000f8000000000000000000000024000000400000000000000000000000000480124010004020008001000002101000000008080000000400100000
B0[357] <= 640'hffffffffffffffffffffbfffffe0fffc3ffc0818c00f0000000000000000000008800000000400000000000000000000000002400124002000000800400000000020000000000042000000000900200
B0[358] <= 640'hffffffffffffffffffffffffffcfffff8ffc0000000e000c1c0000000000000008000080000200000000000000000000000000404002060210084000009000000000000000004000000000000000000
B0[359] <= 640'hffffffffffffffffffff99f9f7fffffff00ff000007e0000000000000000000000000080004000000000000000000000000008004240010100000000000800002000000000000001000000000000000
B0[360] <= 640'hfffffffffffffffffffffffffffffffffe0fffe3ffee0000000000000000000000400080000000000000000000000000000004000000008001200001001800000000000000000009000000000000000
B0[361] <= 640'hfffffffffffffffffffffffffffffffffffffffff8000000000000000000000400408080000000000000000000000000000000800102204001004800800000000000000000000008000000000000000
B0[362] <= 640'hfe00fffffffffffffffffffffffffffffffffff80000000000000000000000000000218000000000000000000000000000000000000000010008c042000000000000000000000000000000000400000
B0[363] <= 640'hfc003fffffffffffffffffffffffff03ffffffe000001000000000000000000018100100000000000000000000000000000004004000400208804200001000000000000000000000000000000000000
B0[364] <= 640'hf8001ffffffffffffffffffffffffe03bffff7cffffe1c00000000000000000008004010000000000000000000000000000000004000402204204000130000000000000000000000000000000200000
B0[365] <= 640'hf00000fffffffffffffffffffffffe03fffffc3ffffc0000000000000000001000040000000300000000000000000000000000000400000008400000900000400000000000000000000000000000000
B0[366] <= 640'hc000003fffffffffffffffffffffff02ffffffb7fc300000000000000000000000000000200200000000000000000000000000000026000000000000980000000000000201000000000000000000000
B0[367] <= 640'h80000008fffffffffffffffffffffe03ffffffffe6040000000000000000000000826000000000004040000000000000000000000009000008000000890000000000000000000000000000000000000
B0[368] <= 640'h3dffffffffffffffffffff02efffffffef9e0000000000008000000000844000000000000040000000000000000000000100020000000000104000000000000800000000000000000000000
B0[369] <= 640'h3bfffffffffffffffffb027fffffffff973000000000000000000800920100000000000080000000000000000000080020800000004000040000000000000000000000000000000100000
B0[370] <= 640'h7ffffffffffffffff703fffa3ffe1dff8800000000000000000800120100000000000000000000000000000000000010800000004000000000000000000200000000000000000000000
B0[371] <= 640'h800033ffffffffffffffff01c1ff80c3fffb080000200000000000400090c400000000000000000000000000000000000000000000000800804000000001900000000000000000000000000
B0[372] <= 640'hcffffffffffffffe00700077f00f000000000000000000000000909020000000000000000000000000000010000000000802000000800002000000101000000000000000000020000
B0[373] <= 640'h80000031ffffffffffff8001fc00e0ff7f00000000004000000000020968020000000000000000000000000000000000000000100004002800000000000000000000000000000000000000
B0[374] <= 640'h1f00000003fffffffff00000fffc00007f00000000004000000000000060240900000000000000000000000000000000000440000000001000000000000000000000000000000000000000
B0[375] <= 640'h7f0000001fffffffff00000ffffff000000030000002042080000000000000000000000000000000000000000000000000000104000000800000000000000000000000000000000000000
B0[376] <= 640'h1cf000000007ffffff00000ffffffff0008000000000080040000000110800000000000000000000000000000000000010000010000000804000000000000000000000000000000000000
B0[377] <= 640'hfe0000000007fffff00000ffff7ffc03ff800000000080000040000080000000000000000000000000000000000000000000002000000004000000000001000000000000000000000000
B0[378] <= 640'hffc0ff80000067ffec0001fffeffff0f0000002000000000002000009c000000000000000000000000000000000000000000088000080000000000000000000000000000000000000000
B0[379] <= 640'h1ffff69e0000003ff800013fcec1fff80000001f0000800000000000b0400000000000400000000000000000000000000040000000000024000000000000000000000000000000000000
B0[380] <= 640'h3fffe011f00001f7c00013f000027f00000009b8020002000800220b1000000000000000000000000000000000000000000010000000120000000000000000000000000000000000000
B0[381] <= 640'hfbffe000fe000018000176000effe000023077006000300000102022000000000000080000000000000000000000000000000000004000000000000200000000000000000000000000
B0[382] <= 640'h7f007f41000000000001ffc0000000031f1002000040000000000040000000000000000000000020000000000000000000003000001000000000000000000000000000000000000000
B0[383] <= 640'h1fc006ffc00000000001ffe000000400f9e000000050000000000410080000000000000000000020000000000000000000011000000000000000000000000000000000000000000000
B0[384] <= 640'h7ffc01f7fa000000000f8780001f8003efc09000000000000000000000000000000000000000000000000000000000000008800000000000000000000000000000000000000000000
B0[385] <= 640'h3fffc0003fff00f0000000e0407f800a00131800040000008000000000000000000000000000000000000000000000000000400400000000000000000000000000000000000000000
B0[386] <= 640'h1ffffffe30000f80000000302000000120001800000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000
B0[387] <= 640'h3ffffffffc303f80000000e8c000000000e8200000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000
B0[388] <= 640'hfffffffffff63fc80880032800000001f80070000000000000204000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000
B0[389] <= 640'hffff0f310fff3f6000800c00000000f000000000000020000204000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[390] <= 640'h3ffffff0801ff8e7f34c07000200ffc000000000000000000200000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000
B0[391] <= 640'hcfffffffffe7ffffffb201c00703000000000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[392] <= 640'h3fffffffffffeeeffc1980714003000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[393] <= 640'hfffffde3f0fff001fc10012cf9f000000000000000000000048000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[394] <= 640'hfffa801e801ff8040ff000000400000000000000000000c010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[395] <= 640'h1fffffffc00a07fe0fff400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[396] <= 640'h3ffffffffff010ffd05900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[397] <= 640'h1efffffffe9ff9801ff8600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[398] <= 640'hffffffffc00ffff807fd88010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[399] <= 640'h1fff7ff9f0303fffe03777800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[400] <= 640'h3ffffffffffc03fff6018000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[401] <= 640'h1ffffffffffff8000ff90000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[402] <= 640'h1ffffffffffffff807ffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[403] <= 640'h7cfffffffffffffff03ff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[404] <= 640'h3ffe0fff10000fffffc0180000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[405] <= 640'hfffcffc7fff1800bffffc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[406] <= 640'h1ffffffffffff80007fffe000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[407] <= 640'h3fffffffffffffffe3fff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[408] <= 640'h17ffffffffffffffffeff400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[409] <= 640'hf7ffffc3c7801fffffffc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[410] <= 640'h3fffffc1ffff0671ffffff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[411] <= 640'h1ffffffffffffff1331fffe000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[412] <= 640'h7ffffffffffffffffff3f0000000000003000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[413] <= 640'hfffffffffffffffffffffe00000000001c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[414] <= 640'h7fffffffe86f8fffffffff80000000000380000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[415] <= 640'h3ffb06f8dfffc7fbf807ffe00000000000e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[416] <= 640'hfff1ffefffffffffffffff000000000001c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[417] <= 640'h3fffffffffffffffffffffe78000000000f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[418] <= 640'hfffffffffffffffffffffff80000000001e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[419] <= 640'hfffffffe007c7ffffff99e800000000007c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[420] <= 640'hffc013c03fffffffffffff800000000001f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[421] <= 640'h7ff0ffffffffffffffffff8000000000007e000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[422] <= 640'h3ffffffffffffffffffffff000000000001f800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[423] <= 640'h7fffffffffffffff3fffffc000000000007e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[424] <= 640'hffffffffe3ffffffffffff000000000000fc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[425] <= 640'h3fffffffffffffffffffff8000000000003f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[426] <= 640'h1ffffffffffffffffffffff0000000000007c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[427] <= 640'hffffffffffffffffffffffff80000000000e000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[428] <= 640'h3fffffffffffffffffffffffffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[429] <= 640'h7ffff8ffffffffffffffffffffffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[430] <= 640'h1ffffc77fffffffffffffffffffffc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[431] <= 640'hffffffffffffffff7ff1ffffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[432] <= 640'h3ffffffffffffffffffffff86000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[433] <= 640'hffffffffffffffffffffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[434] <= 640'h3fffffffffffffffffffc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[435] <= 640'h7fff00033ffffffffe00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[436] <= 640'h7ff3fffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[437] <= 640'h7fffffffffffe000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[438] <= 640'h1ffffffffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[439] <= 640'hffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[440] <= 640'h3ffffec00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[441] <= 640'h7ff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[442] <= 640'hc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B0[443] <= 640'h0
B0[444] <= 640'h0
B0[445] <= 640'h0
B0[446] <= 640'hc000000000000000000000000000000000
B0[447] <= 640'h0
B0[448] <= 640'h7fc780000000000000000000000000000000000
B0[449] <= 640'h7f7e00000000000000000000000000000000000
B0[450] <= 640'h183c00000000000000000000000000000000000
B0[451] <= 640'h0
B0[452] <= 640'h100000000000000000000000000000000000000000000000000000000000000
B0[453] <= 640'h0
B0[454] <= 640'h3ce000000000000000000000000000000000000000000000000
B0[455] <= 640'h43fffcf000000000000000000000000000000000000000000000000
B0[456] <= 640'h1c000000ffe7f601c3000000000000000000000000000000000000000000000000
B0[457] <= 640'h1ffffc00117700600c7000000000000000000000000000000000000000000000000
B0[458] <= 640'h19fc0000000180000c7000000000000000000000000000000000000000000000000
B0[459] <= 640'h7f301c7800000000000000000000000000000000000000000000000
B0[460] <= 640'h3ffffe7800000000000000000000000000000000000000000000000
B0[461] <= 640'h1fffff7800000000000000000000000000000000000000000000000
B0[462] <= 640'hff0001fffff7e80000000000000000000000000000000000000000000000
B0[463] <= 640'h1cc0001fffff3ef3c00000000000000000000000000000000000000000000
B0[464] <= 640'h7ffff3ef3fc0000000000000000000000000000000000000000000
B0[465] <= 640'h7fff3ef3fe0000000000000000000000000000000000000000000
B0[466] <= 640'hfff3cf3ffc000000000000000000000000000000000000000000
B0[467] <= 640'h0
B0[468] <= 640'h802800000000000000000000000000000000000000000000000000000000000000000000000000000000000001f9cf1ff7000000000000000000000000000000000000000000
B0[469] <= 640'h1c03c0480000000000000000000000000000000000000000000000000000000000000000000000000000000000009cfbffff00000000000000000000000000000000000000000
B0[470] <= 640'h7ffe23c00000000000000000000000000000000000000000000048000000000000000000000000000000000000000004f9ffffc000000000000000000000007f800000000000000
B0[471] <= 640'hfffffe6300000000000000000000000000000000000000000000007700000000000000000000000000000000000000000001fffff00000000000000000000003ff0c0100000000000
B0[472] <= 640'h7bfffffffe600000000000000000000000000000000000000000000000fc0000000000000000000000000000000000000000000003fff000000000000000000000ffff0f1280006000000
B0[473] <= 640'h1ffffffffffe600000000000000000000000000000000000000000000000fe00000000000000000000000ff0000000000000000000001ff800000000000000007f08ffff000000000000000
B0[474] <= 640'hfc00000083ffffffffffe600000000000000000000000000000000000000000000000fe00000000000000000000000e000000000000000000000000180000000000000000ff007fff000000000000000
B0[475] <= 640'hff00000083ffffffffffee00000000000000000000000000000000000000000000000f700000000000000000000000000000000000000000000000000000000000001f3ffff007ffe000180000000000
B0[476] <= 640'hfff9000003e3ffffffffc000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001ffbffffe0ff80004000000000000
B0[477] <= 640'h383f3ffffffff8000000000000000000000000000000000000000000000000000080001f0000000000000000000000000000000000000000000000000403fffbf9ffe8000e000000000000000
B0[478] <= 640'h4fc3fffffffff90000000000000000000000000000000000000000000000000000000001f0000000000000000000000000000000000000000000000000003fff8bfff400380000000006000000
B0[479] <= 640'hfe3fffffffff00000000000000000000000000000000000000000000000000000000001f000000000000000000000000000000000000000000000000000001f0ff800000000000000000e0000
end
always @(posedge vga_clk) begin
B1[0] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[1] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[2] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[3] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[4] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[5] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[6] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[7] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[8] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[9] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[10] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[11] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[12] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[13] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[14] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[15] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[16] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[17] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[18] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[19] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[20] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[21] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[22] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[23] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[24] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[25] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[26] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[27] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[28] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[29] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[30] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[31] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[32] <= 640'he7bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[33] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[34] <= 640'h3ffffffffffffffffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[35] <= 640'hff7ffffffffffffffffc9fffff3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[36] <= 640'hff7fffffffffffffffff9ffffffbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[37] <= 640'he7ffffffffffffffffe3ff7ffff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[38] <= 640'h3ffffffffffffffffe166ffff3fbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[39] <= 640'h18ffffffffffffffffe066effefbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[40] <= 640'h3bfffbffffffffffff8019bb3f99efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[41] <= 640'h3bffffffffffffff7f8098bb07098fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[42] <= 640'h3bfffffffffffe9f7f00009c03067fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[43] <= 640'h3bfffffffffffefff800009c3066fbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[44] <= 640'h3bffffffff3ffffffc00000cc06627ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[45] <= 640'h3bffffffbfffffe61c000000830003ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[46] <= 640'h3bffffff88feff660c0000200300807fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[47] <= 640'hfffffffffc3ffe66c00000203c800e3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[48] <= 640'hffffffffffc4fe8cf8800000008400ff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[49] <= 640'hff7fffffffc03f873e100000000000ff6fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[50] <= 640'h7f7efffffff0ff071f1000000000013fffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[51] <= 640'h3e67fffffff1f938f08000004000009effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[52] <= 640'h3ee7ffffff31f931f08000000000008ebdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[53] <= 640'h3fe7ffffff1339c1e0000000000000033fffffffffffffffffffffffffffffffffffffffffdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[54] <= 640'hff7fffffffcf9981c3000000000000312fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[55] <= 640'hef7effffffcf981ce08000000080013147ff67ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[56] <= 640'hc378dfffff3f6e0060000000c00000869ffffeffffffffffffffffffffffffffffffffff3fdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[57] <= 640'h3ce3ffffffff6e00200000000000000389ffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[58] <= 640'h3ce7ffffffff9801000000030000002081ff7fffffffffffffffffffffffffffffffffe7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[59] <= 640'h3ccf7fffffff9801800000000000000001e7f7fffffffffffffffffffffffffffffffffefeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[60] <= 640'h1f7fffffff980098000000010000070067e7fffffffffffffffffffffffffffffffffedfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[61] <= 640'h813c7ffffffffd001800000000000000001fe7ffefffffffffffffffffffffffffffffe7dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[62] <= 640'h3cffffffffee01100000000000000002997377ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[63] <= 640'h1cffffffffffe7c10000000000000000009831737efffffffffffffffffffffffffffffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[64] <= 640'hdffeffffffff7fc00000000018000000000001eeefffffffffffffffffffffffffffffff4fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[65] <= 640'hffffffffffffffc0f00000000000000000000006fffffffffffffffffffffffffffffffffdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[66] <= 640'hffffffffffffffe4000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[67] <= 640'hfffffffffffffee6000000000000000000000006ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[68] <= 640'hffffffffffffff768000000000000000000000273fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[69] <= 640'hfeffffffffffc7760000000000000000000000223fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[70] <= 640'hffffffffffffcf76000000000000000000000022ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[71] <= 640'hfffeffffffff3e72000000000000000000000076ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[72] <= 640'hfdff7fffffffff0c00000000000000000100060ef3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[73] <= 640'hfffffffffffffcc0c000000000000000200000037fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[74] <= 640'hffffffffffff7cc00000000000000000000000137fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[75] <= 640'hfffffffffffff81c000000000000000000000103ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[76] <= 640'hffffffffffffc0180000000000000000c0000107ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[77] <= 640'hffff7fffffffc1c000000000000000000000000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[78] <= 640'hffffffffffffe0c000000000000000000000000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[79] <= 640'hfffffffffffff800000000000000000080000037f3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[80] <= 640'hffff7ffffff73c80000000000000000000000046c7ff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[81] <= 640'hfffffffffffff00800000000000000000000000406ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[82] <= 640'hffffffffffffc01800000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[83] <= 640'hffffffffffffc00000000000000000008000000100ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[84] <= 640'hfffffffffff7fc8000000000000000000000000001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[85] <= 640'hfffffffffff73c00000000000000000000000000000fbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[86] <= 640'hffffffffffff3c00c0000000000000000000000000061fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[87] <= 640'hfffffffffbfe008000000000000000000000000000001f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[88] <= 640'hff7fffffffccbf81000000000000000000000000008efefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3ffffffffffffffffffffffff
B1[89] <= 640'hffffffffffdcb38000000000000000000000000000047fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[90] <= 640'hfffffffffffe92000000000000000000000000000000ffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[91] <= 640'hfffffffffefe82000000000000000000000000000001fffffffffffffffffffffffffffffffffff39ffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffffffffffffffffffff
B1[92] <= 640'hfffffffffee0be7800000000000000000000000000637fffffffffffffffffffffffffffffffff71ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[93] <= 640'hfffffffff7e0bef000000000000000000000000004f7ffffffffffffffffffffffffffffffffff79ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[94] <= 640'hffffffffffe1b7c000000000000000000000000006ffffffffffffffffffffffffffffffffffffe03fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[95] <= 640'hbffffffffef3b7e0800000000000000000000000047fffffffffffffffffffffffffffffffffffe07f7ffffffffffffffffffffffffffffffffffffffffffffffffffffbefffffffffffffffffffffff
B1[96] <= 640'hfe7fffffe6cffefc000000000000000000000000003fffffffffffffffffffffffffffffffffffdb1ffffffffffffffffffffffffffffffffffffffffffffffffffffff731fff7ffffffffffffffffff
B1[97] <= 640'hfffffffff7efffff00000000000000000000000000bfffffffffffffffffffffffffffffffffffe01f7ffffffffffffffffffffffffffffffffffffffffffffffffffff008ffffffffffffffffffffff
B1[98] <= 640'hffffffffffffcff380000000000000000000000011fffffffffffffffffffffffffffffffffffec11f3ffffffffff1fffffffffffffffffffffffffffffffffffffffff08c7fffffffffffffffffffff
B1[99] <= 640'hffffffff99ffeff30000000000000000000000001fffffffffffffffffffffffffffffffffffffdf1f07efffffff0070fffffffffffffffffffffffffffffffffffffef0803ffdffffffffffffffffff
B1[100] <= 640'hffffffff9ff9fffb0000000000000000000000010ffffffffffffffffffffffffffffffffffffff807c3effffffc003003fffffffffffffffffffffffffffffffffffff0003df97fffffffffffffffff
B1[101] <= 640'hffffffffbff9ff7e000000000000000000000000cfffffffffffffffffffffffffffffffffffff980710efe7fff8000007ffffffffffffffffffffffffffffffffffffc00038717fffffffffffffffff
B1[102] <= 640'hffffffffeff9fe7a000000000000000000000000ffffffffffffffffffffffffffffffffffffff190600edc3ffc000000ffffffffffffffffffffffffffffffffffffd000000607fffffffffffffffff
B1[103] <= 640'hffffffffc6fb8ef3000000000000000000000004ffffffffffffffffffffffffffffffffffffdff96603e00099c0000004fffffffffffffffffffffffffffffffffff0000000647fffffffffffffffff
B1[104] <= 640'hffffffffffff9970800000000000000000000019fffffffffffffffffffffffffffef1ffffffe7c1630001806c80000000ffffffffffffffffffffffffffffffffff00800000f0cfffffffffffffffff
B1[105] <= 640'hfffffffc7fff8920800000000000000000000019ffffffffffffffffffffffffffff07ffffffe7ff0700010041000000007ffffffffffffffffffffffffffffffffc00000000f1ffffffffffffffffff
B1[106] <= 640'hffffffff7fffe62000000000000000000000001fffffffffffffffffffffffff7fdfc4ffffff7fdc0600000041000000003ffffffffffffffffffffffffffffffe00000001015fffffffffffffffffff
B1[107] <= 640'hffffffffc7ffe60000000000000000000000000fffffffffffffffffffffffff7ec0c07fffff7fcc0000000040000000003ffffffffffffffffffffffffffffffc00000000c3cfffffffffffffffffff
B1[108] <= 640'hfffffefee7ff6e00000000000000000000000007fffffffffffffffffffffffde080001f7ff331c00000000040000000001fffffffffffffffffffffffffffff7000000000ffcfffffffffffffffffff
B1[109] <= 640'hfffffece7fff0c00000000000000000000000007fffffffffffffffffffffffcc000000f7df100800000000000000000000ffffffffffffffffffffffffffffb6000000000c7ffffffffffffffffffff
B1[110] <= 640'hffffffff1eff8080000000000000000000000007ffffffffffffffffffffffff0000000e410101000000000000000000000ffffffffffffffffffffffffffffe0000000400ffffffffffffffffffffff
B1[111] <= 640'hfffffffc03ff8000000000000000000000000027feffffffffffffffffffffcd000000000104010000000000400000000007fffffffffffffffffff7fffffdbe8000000401ffffffffffffffffffffff
B1[112] <= 640'hffffff7099ffc000100000000000000000000003f9ffffffffffffffffffff7c000000000000000000000001200000000003fffffffffffffffffffbfffefffe80000001001fffffffffffffffffffff
B1[113] <= 640'hfffffffc11ffc0000800000000000000000000017dffffffffffffffffffff60000000000000000000000000000000000007ffffffffffffffffffffff36fefc8000000103ffffffffffffffffffffff
B1[114] <= 640'hffffffce33ff00000400000000000000000000017cffffffffffffffffffff60000000000000000000000000000000000007ffffffffffffffffffbfff337c380000001ff3ffffffffffffffffffffff
B1[115] <= 640'hffffffcc63ff00000600000000003400000000007cffffffffffffffffffffe8000000000000000000000000000000000007ffffffffffffffffffffe01303700000001ffbffffffffffffffffffffff
B1[116] <= 640'h1ffffff887ff80000400000000003c00000000006f3ffffffffffffffffffffc000000000000000000000000000000000003fffffffffffffffffffff08003f00000003fffffffffffffffffffffffff
B1[117] <= 640'h7effff300eff8000000000000000e300000000006f3fffffffffffffffffff4c000000000000000000000000000000000001fffffffffffffffffffec00018600000003fffffffffffffffffffffffff
B1[118] <= 640'hfcffff0006ff8000000000000011fb80000000000cbfffffffffffffffffff78000000000000000000000000000000000001ffffffffffffffffffefc00010000000012fffffffffffffffffffffffff
B1[119] <= 640'hcf9fd80007ff0000000000000061fef90000000009bbffffffffffffffffff7100000000000000000000000000000000000038fffffffffffffffffffc1001000000000fffffffffffffffffffffffff
B1[120] <= 640'hfcfefc00027f80000000000000707ee00000000000c0ffffffffffffffffff8800000000000000000000000000000000000272ffffffffffffffffffffc680000000003fffffffffffffffffffffffff
B1[121] <= 640'h1cff3e0000ff8000000000000020e3f30000170000007ffffffffffffffffff800000000000000000000000000000000000002fffffffffffffffffffffe00800000033fffffffffffffffffffffffff
B1[122] <= 640'h1e0f3c0000ff90100c010000000003f00000bfdf80007ffffffffffffffffff800000000000000000000000000000000000003fffffffffffffffffffffe03c0000003ffffffffffffffffffffffffff
B1[123] <= 640'hc600c00001ffd0000c200000000000000001fbfffcffffffffffffffffffff38000000000000000000000000000000000000037ffffffffffffffffffffff300000003ffffffffffffffffffffffffff
B1[124] <= 640'h8000030001ffc980771c0000001c000f0020bfffffffffffffffffffffffff00000000000000000000000000000000000000167ffffffffffffffffffffffb18000003ffffffffffffffffffffffffff
B1[125] <= 640'hffff8073c008000000800000107fffffffffffffffffffffffffc000000000000000000000000000000000000010fcfffffffffffffffffffffff0000003ffffffffffffffffffffffffff
B1[126] <= 640'hfffc307fc31c0000000100b001767ffffffffffffffffffffffff900000000001860000000000000000000000000e037fffffffffffffffffffffc00008fffffffffffffffffffffffffff
B1[127] <= 640'h10001fffe7f3ef30001068ff8fe3881773ffffffffffffffffffffffffbe0000000011fe00000000000000000000000008023fffffffffffffffffffffc00023fffffffffffffffffffffffffff
B1[128] <= 640'h11ffd5effdfff60037ff7fbdce0f9fffffffffffffffffffffffffff000000003ffc000000000000000000000000000007ffffffffffffffffffffe800f3fffffffffffffffffffffffffff
B1[129] <= 640'h3ffdffffff7e0003fff7fffd61f1fffffffffffffffffffffffffff000000007fff000000000000000000000000000007ffffffffffffffffffffe800fffffffffffffffffffffffffffff
B1[130] <= 640'h167fdfbfff83f8021fffe9f79f1fe7fffffffffffffffffffffffff6000000007fff000000000000000000000000000003bbfffffffffffffffffff80ffffffffffffffffffffffffffffff
B1[131] <= 640'h16ffff9fff8338470fffc103339ffff7ffffffffffffffffffffff76000000003fff800000000000000000000000000001b0fffffffffffffffffff00ffffffffffffffffffffffffffffff
B1[132] <= 640'h7fff9cefce03c07fff980000097efffffffffffffffffffffffff3e000000003fff8000000000000000000000000000000007fffffffffffffffffc77fffffffffffffffffffffffffffff
B1[133] <= 640'h7fff9cc0cf00e0dfff90000081fec7fffffffffffffffffffffff30000000001ffe0000000000000000000000000000000003fffffffffffffffffffffffffffffffffffffffffffffffff
B1[134] <= 640'h9ffd6400cf9e20fefff0000000f9007fffffffffffffffffffff300000000000ffc0000000000000000000000000000000000037ffffffffffffffffffffffffffffffffffffffffffffff
B1[135] <= 640'h8fff66007fcf00fffff000000081001c7fffffffffffffffffff100000000000ff00000000000000000000000000000000000003ffffffffffffffffffffffffffffffffffffffffffffff
B1[136] <= 640'h26fc20111983387ffff80000008000003ffffffffffffffffffc0000000000000000000000000000000000000000000000000001ffffffffffffffffffffffffffffffffffffffffffffff
B1[137] <= 640'h7ffc0011807c17fff180000000000003fffffffffffffffffffc0000000000000000000000000000000000000000000000000007fffffffffffffffffffffffffffffffffffffffffffff
B1[138] <= 640'h6c18080000c83d9fffc00000000000007fffffffffffffffffe000000000000600000000000000000000000000000000000000000f3ffffffffffffffffffffffffffffffffffffffffff
B1[139] <= 640'h800099ffec00000000000017fffffffffffffffffe00000000000060000000000000000000000000000000000000000033ffffffffffffffffffffffffffffffffffffffffff
B1[140] <= 640'h280000000800099ff0600000000000016e7fffffffffffffff600000000000000000000000000000000000000000000000000000007ffffffffffffffffffffffffffffffffffffffffff
B1[141] <= 640'h1bffec00000000000003fffffffffffffffff300000000000000000000000000000000000000000000000000000003ffffffffffffffffffffffffffffffffffffffffff
B1[142] <= 640'h100037ff8000000000000069ffffffffffffffff300000000000000000000000000000000000000000000000000000001ffffffffffffffffffffffffffffffffffffffffff
B1[143] <= 640'h1000000000000003f19000000000000069fbffffffffffffffe80000000000000000000000000000000000000000000000000000018ffffffffffffffffffffffffffffffffffffffffff
B1[144] <= 640'h20000000000010426837fffffffffffff00000000000000000000000002400000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffff
B1[145] <= 640'h8000000000008000007fffffffffffffc000000000000000010000000000000000000000000000000020000fffffffffffffffffffffffffffffffffffffffffff
B1[146] <= 640'h1008000000000000000002fffffffffffffc000000000000000000000000018000000000000000000000000000fffffffffffffffffffffffffffffffffffffffffff
B1[147] <= 640'h10000000000000000000067ffffffffffff8000008000000000c0013c9180b8000000000000000000000040017fffffffffffffffffffffffffffffffffffffffffff
B1[148] <= 640'h8000000000000000001f7fffffffffffd0000009f000000000ffe11f982110000000000000000000000cc83e0ffffffffffffffffffffffffffffffffffffffffff
B1[149] <= 640'h1ffffffffffffed000000dfc30000000ffffff9b7010000000000080000000003ffe3f0ffffffffffffffffffffffffffffffffffffffffff
B1[150] <= 640'h10000000000000000013ffffffeffffcd000105e4c00000005ffffffffff08c810020000d8800000001fffff9ffffffffffffffffffffffffff190fffffffffffff
B1[151] <= 640'h1000000000000000011e3ffffff7fffc981000864180000004ffffffffefe8f1bf0c6000999000000003fffffffffffffffffffffffffffffcc39017fffffffffff
B1[152] <= 640'h1001000000000000000000000000000084deffffffffffc10000836d800000010fffffffffe707e3ff00c83b8fc00000007fffffffffffffffffffffffffffff0001017fffffffffff
B1[153] <= 640'h100000000000000000000000000000000ffefffffffffff80600007c800000007fffffffffe70ffedf0f40fdf03ec000003fffffffffffffffffffffffffffff000101ffffffffffff
B1[154] <= 640'h10000000000001000180000000000000000000000000007fcfffffffffffc0700007c000000007ffffffffffffffeffff69fe73668001c0019ffffffffffffffffffffffffffe000000ffffffffffff
B1[155] <= 640'h88000000000000200000000000000000000000000000003fffffffffffffc06010168000000007fffffffff7edefffffffdff73e23c00fc000ffffffffffffffffffffffffffe400000dfffffffffff
B1[156] <= 640'h18c0000000000002030000000000000000000000000000017bfffffffffffffec00040000000027fffffffff78840fffffff7ff1e7fc001e01005fffffffffffffffffffffffff400081ffffffffffff
B1[157] <= 640'h98100000000000383c000010000000000000000000000007bffffffffffff7fe00c40008000037ffffffffe810001ffffffffff7fe40003c1601fffffffffffffffffffffffff000081ffffffffffff
B1[158] <= 640'h9b27000000000003fffc0001000000000000000000000006737fffffffffff7fff3c4000c100037ffffffffe8000007ffffffffffdf3010700603ffffffffffffffffffffffffe8000017fffffffffff
B1[159] <= 640'h18f0800000000003fffc0018810000000000000000000002e17ffffeffffff7ffef34c187374077fffffffe400000007ffffffffdfff813e3d761ffffffffffffffffffffffffc8000017fffffffffff
B1[160] <= 640'hcf8402000000003fffe00000080000000000000000000008ffdffffffffffffffe0f8b83fff1fffffffffc80000003fcffffffeefffc0ffcfc318feffffffffffffffffffffd8000000ffffffffffff
B1[161] <= 640'h87f8400001000003ffff8000000000000000000000000000007fffffff7ffffffffde739ffff1ffffffffff80000003f3ffffffffeffc0dffefc0197fffffffffffffffffffff80000003fffffffffff
B1[162] <= 640'hc7b84c0001000003ffffc00000000000000000000000000001fffffffffffffffffffff9ffff7ffffffffff00000003f7fffffff7fffc1fff8f80107fffffffffffffffffffff80000009fffffffffff
B1[163] <= 640'h6e1b6c0010000001ffffe10060000000000000000000000003fdfffffffffffffffffffffffffffffffffff0000001fff3fffff97fff013ef3e000037bfffffffffffffffffffc8000008fffffffffff
B1[164] <= 640'h7e83fd0000000000ffffe000600000000000000000000000006d7ffffeffffffffffffdffffffffffffffffc000001effffffffbfffe487fefc00803f9fffffffffffffffffffc0000008fffffffffff
B1[165] <= 640'h6781cd80810000007fff98000000000000000000000000000049ffff3f7fffffffffffdffffffffffffffffe4c30010fffffffffffe00c831e000011fffffffffffffffffffff40000001fffffffffff
B1[166] <= 640'he391fd80010000277fff8e008000000000000000000000000000ffff7f7dffffffffffffffffffffffffffff6ff801bfffffffff7d00000338000010fffffffffffffffffff9e41000003bffffffffff
B1[167] <= 640'h62bffd1c18800007ffff84009800000000000000000000000001ffffe6f9fffffffffffbffffffffffffffffeffe19ffffffffffe100000021c000101dffffffffffffffffff06000000c3ffffffffff
B1[168] <= 640'h9c6fffc000643007ffffff60c000000000000000000000000001ffffccffffffffffefffffffffffffffffffffffffffffffffee60000000208000019ffffffffffffffffffff600000001ffffffffff
B1[169] <= 640'h83fdffc000fe080efffffc2306000000000000000000000000007fffffc0ffffff7ffdffff7fffffffffffffffffffffffffffee00000000000000001ffffffffffffffffffff600000007ffffffffff
B1[170] <= 640'ha3cdffcc1ef88edefffffc220200000000000000000000000006ffffefe07ffffffffdfffffffffffffffffffffffffffffffffc00000000000000000b7fffffffffffffffffff00000007ffffffffff
B1[171] <= 640'h770fffee1ef98efffffffff0e000000400000000000000000007ffffeffcfffffffffdffffffffffffffffffffffffffffffffc00000000000000000005fffffffffffffffffff00000000ffffffffff
B1[172] <= 640'h764ffff203fffffffffffffe3400000000000000000000000003fffffdfcffffffffd9fffeffffffffffffffffffffffffffffc00000000000000000005effffffffffffffffff00000000ffffffffff
B1[173] <= 640'hf2fdff6303ffff7ffffffffe3c00000000000000000000000007fffffdfc3ffffffff93fffffffffffffffffffffffffffffff800000000000000000000cfffffffffffffffffd800000007fffffffff
B1[174] <= 640'h8279ff7003ffff7ffffffffe700000000000000000000000001fffff7dec1ffffffffc1fbfffffffffffffffffffffffffffff8000000000000000000004ffffffffffffffffffc00000037fffffffff
B1[175] <= 640'h9a61ff7e33fffffffffffffc638004000000000000000000001fffff7feffffef9efe77ffffffffffffffffffffffffffffff99000000000000000000004fffffffffffffffffff0002007ffffffffff
B1[176] <= 640'hf973ff7f36ffffffffffffff731c00000000000000000000001fffff7fff7ffffffff9ffffffffffffffffffffffffffffffffc000000000000000000001ffffffffffffffff87ff000007ffffffffff
B1[177] <= 640'hbf79fc7f67ffffffffffffff73cc00000000000000000000000fffffffedffffffffff1fffffffffffffffffffffffffffffff0000000000000000000001fffffffffffffffffffe0012cfffffffffff
B1[178] <= 640'h1d383ceee7ffffffffffffffe7c400000000000000000000000fffffffebffffffefffffffffffffffffffffffffffffffffffe000000000000000000000fffffffffffffffffffc0002cfffffffffff
B1[179] <= 640'h988001ce27ffffffffffffffffc790000000000000000000003fffffffedfffffffefffffffffffffffffffffffffffffffffff800000000000000000000fffffffffffffffffffc0012ffffffffffff
B1[180] <= 640'h8180808f67fffffffffffffffefef1e00000000006000000003fffffffecfffffffefffffffffffffffffffffffffffffffffffcc00000000000000000003ffffffffffffffffff800bfffffffffffff
B1[181] <= 640'h8100789fe3fffffffffffffffefe1bf00000000006800000007ffffffffcfffefbdffffffffffffffffffffffffffffffffffffde04000000000000000003f3ffffffffbffffffc00016ffffffffffff
B1[182] <= 640'hc1001099e7fffffffffffffffffe9b700000000000900000003ffffffffdfffeffdffeffffffffffffffffffffffffffffffffff6c4000000000000000003ffff9fe7600ffffffe00102ffffffffffff
B1[183] <= 640'hf83003b93cfffffffffffffffffefbf00000000001160000003fffffff7bffffdffffeffffffffffffffffffffffffffffffffff7d6000000080000000003fff81016000cf9ffffc01bfffffffffffff
B1[184] <= 640'he0010086c6fffffffffffffffff9f7fc0000000004f8000002f9ffffffcf7f3fef7ffffffffffffffffffffffffffffffffffffffe1c00800000000001003f8300000001303cffc09876ffffffffffff
B1[185] <= 640'h1c06ffffffffffffffffffeff80000000005f8e398007b7ffffdc07ff8feffffffffffffffffffffffffffffffffffffffff1f01180030000000037f92000000000111ffc099e7ffffffffffff
B1[186] <= 640'h1c00ffffffffffffffffffffec000000000fffe380004ffffff9e0fffefecfffbfffffffffffffffffffffffffffffffffff87811e7c7000000003ffb00000000000003ffc1fdfffffffffffff
B1[187] <= 640'h8100ffffffffffffffffffffce000000000ffffff9006ffffff9014fffffdffe9ffffffffffffffffffffffffffffffffffffeffe6fe00000000ffff9000000000000007f89bfdffffffffffff
B1[188] <= 640'h8100fffffffffffffffffffffe000000004fffffff906ffffff800cf7cfffefeffffffffffffffffffffffffffffffffffffff3fe6ffff000001ffff80000000000000033bfbfdffffffffffff
B1[189] <= 640'h3ffffffffffffffffffffe000000004ffffff8907fffffe000e779fffffffbefffffffffffffffffffffffffffffffffff7ffff8ff0000033fff800000000000000003b9dfffffffffffff
B1[190] <= 640'h3fffffffffffffffffffff00000000df7fffff907fffffe0c0e607ffffffffe7ffffffffffffffffffffffffffffffffffffff3cff060001ffff80000000000000003339e7ffffffffffff
B1[191] <= 640'h3fffffffffffffffffffff60000000fffffff3915dfffb200002c0fef7ffce7fffffffffffffffffffffffffffffffffffffd93eff060718ffffb00000000000000071397effffffffffff
B1[192] <= 640'h7ffffffffffffffffffff81000001ffffffff7c3f7ffca0801cc107fc38200ffffffffffffffffffffffffffff7fffffffffff97fe3fed3ffffc800000000000000882e0fcfffffffffff
B1[193] <= 640'hfffffffffffffffffffff81c00001ffffffffe7fffff9830031f06ffff83887ffffffffffffffffffffffffffffffffffffffffffffffffffffc80000000000000000c01ffeffffffffff
B1[194] <= 640'h3ffffffffffffffffffff63c00003ffff7fffe7ffff71377173fceffffe1c83fffffffffffffffffffffffffffffffffffffffffffffffffffffdcc00000000000000001fffffffffffff
B1[195] <= 640'h1ff7fffffffffffffffff76007003fffffffffffffff83e7973fecefee60007ffffffffffffffffffffffffffdffffffffffffffffffffffffffffc00000000000000009f7fffffffffff
B1[196] <= 640'h1fffc3fffffffffffffff7680c3e3fffffefffffffffc329f7ffffffee6801fffffffffffffffffffffffffffdfffffffffffffffffffffffffffff008000000000200007ffffffffffff
B1[197] <= 640'h27ec1ffffffffffffffffec1c77fffffffffffffff9fb38ffffffffee6c003fffffffffffffffdbfffffffffffffffffffffffffffffffffffffffc1f200000000000007ffffffffffff
B1[198] <= 640'h400ffffffffffffffffcffff7fffffffffffffffffb7f7fffffffef90003fffffffffffffffffffffffffffffffffffffffffffffffffffffffffff600000000000007ffffffffffff
B1[199] <= 640'h20000fffffffffffffffdf1ffffffffffffffffffeff3ef3ff7fffef9100137fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000001fffffffffffff
B1[200] <= 640'h7fffffffffffffff67f7ffffffffffffffffffcfb7cffffffff7e0c23dfffffffffff7bffffffffffffffffffffffffffffffffffffffffffffffde20000000001fffffffffffff
B1[201] <= 640'h3fffffffffffffffefffffffffffffffffffffeffffffffffffe30477fffffffffffffbffffffffffffffffffffffffffffffffffffffffffffffff00004000000fffffffffffff
B1[202] <= 640'h3fffffffffffffffc7ffffffffffffffffffffffffffffffffee300ffffffffffffdbf37ffffffffffffffffffffffffffffffffffffffffffffffff8004800003fffffffffffff
B1[203] <= 640'h1fffffffffffffff33ffffffffffffffffffffffffffffffffe6080fffffffffffe81017ffffffffffffffffffffffffffffffffffffffffffffffffe0f7d00007effffffffffff
B1[204] <= 640'hfffffffffffffff13fffffffffffffffffffffff7fffffffff7680fefbfffffffed8007dfffffffffffffffffffffffffffffffffffffffffffffffff8fdf0007fffffffffffff
B1[205] <= 640'hbffffffffffffffc3ffffffffffffffffffffffffffffffeffe300fce1fffffffc98187c3fffffffffffffffffffffffffffffffffffffffffffffffffff9330efffffffffffff
B1[206] <= 640'hfffffffffffffffc3ffffffffffff77fffffffffffffffff9c0000fcc07fffff798080003ffffffffffffffffffffffffffffffffffffffffffffffefffffb7bffffffffffffff
B1[207] <= 640'h3000000000000007ffffffffffffffc3fffffffffffff7fffffffffffffffff1c00001c0466fefee181000077fffffffffffffffffffffffffffffffffffffffffffffffffff9ffffffffffffffff
B1[208] <= 640'h680000000000000ffffffffffffffff7fffffffffff7ffffffffffffffffffc00000042903df0ff000400007ffffffffffffffffffffffffffffffffffffffffffffffffffbeffcffffffffffffff
B1[209] <= 640'h6000000000000000ffffffffffffff83ffffffffffffffffffffffffffffcff800000400013f97c000000001fffffffffffffffffffffffffffffffffffffffffffffffffffcfffffffffffffffff
B1[210] <= 640'h1c00000001fffffffffe33ffe7ffffffffffffffffffffffff3fffeff810000380003387800000000037ffffbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
B1[211] <= 640'hc00238000000003ffffffff00001cffffffffffffcffffffffffff7ff7ffc000001980000383800000000003fff810007ffffffffffffffffffffffffffffffffffffffffffffffffffefffffff
B1[212] <= 640'hc03fe0000000001ffffffff000038fffffffffffff0ffffffffffffffe67c0000079800203800000000000010fe000001ffffffffffffffffffffffffffffffffffffffffffffffffffafffffff
B1[213] <= 640'h10033fef8240000017ffffffe000038fffffffffffe307fffffffffb7ffe40700000398000030800000000000033c0000003fffffffffffffffffffffffffffffffffffffffffff7fffff8fffffff
B1[214] <= 640'h17ffffb600000000b7fe018000000fffffffffffc0307fffffffff7fe0f030000017e000100800000000000000800000001ffffffffffffffffffffffffffffffffffffffffffffffffc7ffffff
B1[215] <= 640'h217fffefff000000003cc0000000001ffffffffff80007fffffffffffe98000000017e0008000000000000000000000000003fffffffffffffffffffffffffffffffffffffffffffffff87ffffff
B1[216] <= 640'hffffffff600000000460000000007fffffffffec8000ffffffffffff86000000000f0000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffec4ffffff
B1[217] <= 640'h1fffffffff00000000000000000003fffffffff400000fffffffffffe07000000000f00000000000000000000000000000007fffffffffffffffffffffffffffffffffffffffffffffec5ffffff
B1[218] <= 640'h40003ffffffffe00000000000000000003fffffffff0000007fffffffff7e00000000000700000000000000000000000000000000effffffffffffffffffffffffffffffffffffffffffffa64ffffef
B1[219] <= 640'h8003fffffffffe0000000000000000000fffffffffc8000003fffffffffff800000000003c00000000000000000000000000000004fffffffffffffffffffffffffffffffffffffffffffff46fffff7
B1[220] <= 640'h3fffffffffc0000000000000000007ffffffffc8000011e0ffffffeff8000000000c3e00000000000000000000000000000000dffffffffffffffffffffffffffffffffffffffffffffc6ffffff
B1[221] <= 640'h8183c3ffffffffdf0000000000000000001fffefffb80000008c03b9dffffc0000000000e1c0000000000000000000000000000000017fffffffffffffffffffffffffffffffffffffffffff347ffffb
B1[222] <= 640'hb1e7ffffffffffdffc00000000000000003fffefff800000000100110eff3800000000002000000000000000000000000000000000017fffffffffffffffffffffffffffffffffffffffffff303ffffb
B1[223] <= 640'h397ffffffffffffffe0000000000000000ffff7cff80000000010000dc7e800000000000201800000000000000000000000000000001fffffffffffffffffffffffffffffffffffffffffff5a27fffe9
B1[224] <= 640'h76ffffffffffffffff8000000000000001fffff018000000000000005c6f98000001000000c0000000000000000000000000000000007fffffffffffffffffffffffffffffffffffffffffff9277fff9
B1[225] <= 640'h67ffffffffffffffff8000000000000000ffffc00000000000000000083e9800000000000730000000000000000000000000000000003ffffffffffffffffffffffffffffffffff7defffff7166dfffd
B1[226] <= 640'hfffffffffffffffffff800000000000000ffff000000000000000000003c6000000000006018000000000000000000000000000000000fffffffffffffffffffffffffffffffffed9ffffff7926cfffc
B1[227] <= 640'hf9ffffffffffffffffff00000000000001fffc0000000000000000000000600000000000e0000000000000000000000000000000000007fffffffffffffffffffffffffffffffffeddfffee3484c3df8
B1[228] <= 640'hfdffffffffffffffffff00000000000001fff0000000000000000000000000000000000000000000000000000000000000000000000007ffffffffffffffffffffffffffffffffbedbfffee96a247ff8
B1[229] <= 640'hffffffffffffffffffff80000000000001ffe0000000000000000000000000000000000000000000000000000000000000000000000007ffffffffffffffffffffffffffffffffb4f3fffff89820efd8
B1[230] <= 640'hffffffffffffffffffffe00000000000007f00000000000000000000000000000000000000000000000000000000000000000000000007ffffffffffffffffffffffffffffffffc911fffff0ca64ffd8
B1[231] <= 640'hffffffffffffffffffffe00000000000007e00000000000000000000000000000000000000000000000000000000000000000000000007fffffffffffffffffffffffffffffffff39a3ffff0c009bf5c
B1[232] <= 640'hffffffffffffffffffffe00000000000007c00000000000000000000000000000000000000000000000000000000000000000000000003fffffffffffffffffffffffffffffffff1867ffff0c0089ed8
B1[233] <= 640'hfffffffffffffffffffff00000000000003800000000000000000000000000000000000000000000000000000000000000000000000003ffffffffffffffffffffffffffffffff044467ffc811206e44
B1[234] <= 640'hfffffffffffffffffffffa0000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ffffffffffffffffffffffffffffffffa8449ffb705a30cf2c
B1[235] <= 640'hfffffffffffffffffffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ffffffffffffffffffffffffffffffff3b116fff2468218f26
B1[236] <= 640'hfffffffffffffffffffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ffffffffffffffffffffffffffffffff92133ffe252c232602
B1[237] <= 640'hffffffffffffffffffeff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffffffffffffffffffffffefda155fff340121cd03
B1[238] <= 640'hffffffffffffffffffdff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffffffffffffffffffffffefe4c4d7ff38890f4d0c
B1[239] <= 640'hfffffffffffffffffffe10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffffffffffffffffffffffef90ce39ee0c0905c544
B1[240] <= 640'hfffffffffffffffffff800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffffffffffffffffffffffaf500e5fbb18b005dd2e
B1[241] <= 640'hffffffffffffffffff1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffffffffffffffffffffff96280e01fb1a400ed820
B1[242] <= 640'hffffffffffffffffc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fffffffffffffffffffffffffffffc238c4c75f98e111ec005
B1[243] <= 640'hffffffffffffff3ec000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fff7ffffffffffffffffffffffffffdfc4102afda8317be706
B1[244] <= 640'hffffffffffffff3fe000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffefffffffffffffffffffffffffffc7c22461f81798472623
B1[245] <= 640'hffffffffffffffc3f80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000efffffffffffffffffffffbffffe3a001461f88bcc0230b2
B1[246] <= 640'hffffffffffffffc1200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffffffff9ffff3ffffe018015a0fd4bcc42713b
B1[247] <= 640'hfffffffffffffff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fcfffffffffffffff9ffff2ffffc2a8010b1f7a3e40f598d
B1[248] <= 640'hff1ffccffeffc3f800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffbffbf2ffff81de43060fe00520e1831
B1[249] <= 640'h31cff87fffff03f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffffffffffffffffefdfeaefff3c3819047ff802c0ad212
B1[250] <= 640'hc0801effff8300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fffffff00407d59fbd2ffc77df3127610024efbc762a1452
B1[251] <= 640'hfffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffff0000000000779feb8a55f16f1941857aff68cc1a481
B1[252] <= 640'h7ffffc80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ffffc00000000003d223ae5e7f13740c926bbf48e81ab068
B1[253] <= 640'h8013ffffc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff0000000000017ae7fa47febb6265221a9d40b11ab0ec
B1[254] <= 640'hfff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fe00000000000168e9fb99ff912642a006148124319964
B1[255] <= 640'hd46edbad1ffcf0e791a8a2fa2b032c490
B1[256] <= 640'h5fe2fca54ff474a0b88c131e94f28c480
B1[257] <= 640'h45b3255212ffe56003209083f8476c2422
B1[258] <= 640'h400000000000000608bfd6f3b63ffc077cf910017bf04238040
B1[259] <= 640'hef000000000000000035fe0c3bbff9330c4408b90f9c2078010
B1[260] <= 640'hfc0000000000000000000000000000000000000000000000c0000000000000000000000000000000000000000013fff0000000000000009b9b2a117794f9a4944902bfc602ac320
B1[261] <= 640'h7e300000000000000000000000000000000000000000000180000000000000000000000000000000000000000007fff000000000000002c555daf14b0e5b31340a0867c11364258
B1[262] <= 640'h2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010c000000000000001eb20b800896ae40114111a13770112404
B1[263] <= 640'h60000000000000000000fee00000000000000000000000000000000000800000001800000000000000000000000000000000000000000000000001675b50a52c420d5c10a64d0bef023242bc
B1[264] <= 640'h7fffe8000000000000000000000000000000000000000000300000280000000000000000000000000000000000000000009afc3ee100c69ac55ac272e87c530326795
B1[265] <= 640'h7ffffe000000000000000000000000000000000000000000ff8ff1ff0000000000000000000000000000000000000000001ac1a5123007d1f6c9a686a4ba5813c2c11
B1[266] <= 640'h1fffffffffe0000000000000800000000000001c0000000000fffffffffe00000000000000000000000000000000000000000814142348052d3e2c5c184800a8002f7d80
B1[267] <= 640'h7f000000000000003ffffffffff8000000000001c00000000000003f8000000000fffffffffe000000000000000000000000000000000000000008dc24044189389206c985981b70043615b9
B1[268] <= 640'hffe00000000000007fffffffffff810000000011c00000000000007fe000000000ff807fffff000000000000000100000000000000000000000000fb3c4d88218ae4d3c0cce809fc2ab32281
B1[269] <= 640'hfff00e0000000007ffffffffffffff000000003bc0000000000000fff000000001ff007fffff0000000000000003e0000000000000000000000000be016bbc02a244f141c1f310a723a04828
B1[270] <= 640'hfcf1ffc0000000cfffffffffffffffff000000ffc0000000000000fffc00000003ff001fffff7ffc00000000001fffe000000000000000000000058626af3d85135d7c1b44f4011ab908b956
B1[271] <= 640'h71ff84000000ffffffffffffffffff800106ffc0000000000002fffc00000003ff070fffffffff00000000007ffffc0000000000000000000000a01138b5025582f18084118c25bc9804e4
B1[272] <= 640'h7fff30003ffffffffffffffffffff00000fffe00000000000003fe0000000000707fffffffffffc03c0020fffffff000000000000000000000466b75450026ef2e5722f29258ce6481040
B1[273] <= 640'hc7ffffc3ffffffffffffffffffffff80000fffc00000000000001fc0000000000707fffffffffffe00600fffffffffff000000000000000000164d1129cc00137f29b62196c07c84992e34
B1[274] <= 640'h1ffffffe7ffffffffffffffffffffffe00007f9000000000000001f870000000007007ffffffffffff07c0fffffffffff00000000000000000005374e842893042a200df70214999c050618
B1[275] <= 640'h7c7fffffffffffffffffffffffffffff000c0f8000000000003000007000000000703ffffffffffffffee0fffffffffff00000000000000000031e3d81888915417cee8254269b61d994626
B1[276] <= 640'h7fffffffffffffffffffffffffffffc00e000000000000001000000000000000107ffffffffffffffc61ffffffffffff000000000000000005bd8c50360d9800f8c612421280b709c1700
B1[277] <= 640'hffffffffffffffffffffffffffffffe04e00000000000000000000000000000010ffffffffffffffffc3ffffffffffffe00000000000000000d6a50910cd202f572202487c0188c85089a
B1[278] <= 640'h33f8ffffffffffffffffffffffffffffffff8ec0000000000000000000000000000081001ffffffffffffffeff87ffffffffff00000000000000003a4c7bce72480344fb862313093ba342a9e5
B1[279] <= 640'h1ffffffffffffffffffffffffffffffffffffdfe00000000000000000000000000000c0001fffffffffffffffff03ffffffffff000000000000000061437ea070cb52533b16123928144240782c
B1[280] <= 640'h1fffffffffffffffffffffffffffffffffffe3ff0000000000000000000000000000000001f1ffffffffffffffe007fffffff1f000000000000000004d9b806a412d83cc5ab8790514303844492
B1[281] <= 640'hff803fffffffffffffffffffffffffffffffffffefff8000000000000000000000000000000001f3fffffffffffa7f8007fffffffff000000000000000092f6c0a24ca5da1732a50248844efe417070
B1[282] <= 640'hffff03fffffffffffffffffffffffffffffffffffffff80000000000000000000000000000000000001fffff1ffe07e0003fffffffff00000000000000008efa8da8809c4bb3e431d622448209823718
B1[283] <= 640'hffffc37fffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000031e3fff0fe001000007ffffffff00000000000000008b679b0688154e81cc52d64201c168a13a1e
B1[284] <= 640'hffffff7fffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000071e001f07600000000380ff00000000000000000005e90590b3a668364983c850264a08f0426c45
B1[285] <= 640'hffffffffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000f1e000e06600000000300000000000000000000000685e81371aa9148df6039546f48d34b028208
B1[286] <= 640'hffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000001f1e0006000000000000000000020000000000000000ce467ca0860122584d6c06ba429cd090b886
B1[287] <= 640'hffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000a0a0002000000000000000000000000000000000017470f9973ac442088288311a064043230eb20
B1[288] <= 640'hffffffffffffffffffffffffffffffffffffffffffff8c80000000000000000000000000000000000000000000000000000000000000000000000000000c9592dc97a000e4a46924200d470aebd0600a
B1[289] <= 640'hffffffffffffffffffffffffffffffffffffffffffff8e800000000000000000000000000000000000000000000000000000000000000000000000000006c36dc7c84ac944b130db26bec8765210c34a
B1[290] <= 640'hffffffffffffffffffffffffffffffffffffffffcfff80000000000000000000000000000000000000000000000000000000000000000000000000000081cc511562441c100c2b0d0309328049538084
B1[291] <= 640'hffffffffffffffffffffffffffffffffffffffff87fe8400000000000000000000000000000000000000000000000000000000000000000000000000001036199c388c4c5f43168e02cfa0436103f702
B1[292] <= 640'hffffffffffffffffffffffffffffffffffffffff830000000000000000000000000000000000000000000000000000000000000000000000000000000035800a8c9f4200e21bc05d032fb06ca809451a
B1[293] <= 640'hffffffffffffffffffffffffffffffffffffffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000d30e6c1215700a67c801d84c523ba09f0416a
B1[294] <= 640'hffffffffffffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000000000000000000000000000000000000000000291954535e11c0c41aac64c46938df54f0a111
B1[295] <= 640'hffffffffffffffffffffffffffffffffffffffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000d220dd3c2b84810b386c6421066208bd00120
B1[296] <= 640'hffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000000000000000000000000000000000006aad918f0a419e62f128b066cccf66600dea4
B1[297] <= 640'hffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000000000000000000000000000043df25099dfd092f04f40c4506c1291320b444
B1[298] <= 640'hffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000000000000000000000000000000000000a97c5930580bc1ac6a8ea648f3ccb9a8ea22
B1[299] <= 640'hfffffffffffffffffffffffffffffffffffffffec0000000000000000000000000000000000000000000000000000000000000000000001c000000000012e3fb0e082cd396e18402a48ad2ba50998408
B1[300] <= 640'hfffffffffffffffffffffffffffffffffffffffe80000000000000000000000000000000000000000000000000000000000000000000041ec04000c0105946b640000f45bad312366084c13d38b44c3c
B1[301] <= 640'hffffffffffffffffffffffffffffffffffffffff80000000000000000000018000c000000000000000000000000000000000000000001fdec0085ff4553f83c544026105d75cec34e22f564c4640e400
B1[302] <= 640'hffffffffffffffffffffffffffffffffffffffff00000000000000000000000004000000000000000000000000000000000000000000ffdee40cffffffdf0d6c556a960d4d26d844620672088e29cf12
B1[303] <= 640'hffffffffffffffffffffffffffffffffffffffff000000000000000000000dc07cc00000000000000000000000000000000000000000ffd8ee9eff7fffefac8218806d82082642c2d147441bac35a06b
B1[304] <= 640'hffffffffafffffffffffffffffffffffffffffff80000000000000000000c3e007f800000000000000000000000000000000000000077ffdf76e827fff6dfc0d6d8871409c1846439333d61c82085810
B1[305] <= 640'hffffffff87ffffffffffffffffffffffffffffff800000000000000000033fe07fdc000000000000000000000000000000000000201cffa1ffbc0007ffe1c50a04330a249ace14a9a19f0125e8ac8450
B1[306] <= 640'hffffffff877fffffffffffffffffffffffffffffe0000000000000000019ffc0ffc0000000000000000000000000000000000000001c4f6febfbfffffedb9f08202db14244c8e22883144070a4c46044
B1[307] <= 640'hffffffff071fffffffffffffffffffffffffffffe0000000000000000027ff00ffc000000000000000000000000000000000000000001f921fa3ffffff0ef2c14a07302050026ac572324a8d8f90648b
B1[308] <= 640'hff81ffff000033fffffffffffffffffffffffffff000000000000000001bfc1fffe000000000000000000000000000000000000ffeffff885ff7fffffc4ff626ad4a16618014d64d21d32607be2048d5
B1[309] <= 640'hff81fffe000133ffffffffffffffffffffffffffe000000000000000187fe0fffff0000000000000000000000000001e80009ffffe3f090571e3fffff88869e104a18c23fc1c43ac20e0084a454408a1
B1[310] <= 640'h700000f33ffffffffffffffffff80ffffff00000000000000001cdfc1fbfff80000000000000000000000000fffff0003c000000085f19ffffe7d6febc0a4c022017a2319090145203301b03001
B1[311] <= 640'h700003f33ffffffffffffffffff00fffffe00000000000000000040fffffff800600000000000007cf00000000000000367800000ad79bf13303dddff08958242a002103ea5e1c0f82000700000
B1[312] <= 640'h180000030000ffffffffff00001ffc00000000000000000081ff9ffffc0070000000f902fc7e00000000000000fe3f000000ad33bb10006d9204e1282d5000481322c4d2217f18209cca54
B1[313] <= 640'he0ffffff0000fbfcfcffffff003f000000000000000000fc1fffff7ffc00830000000004000000000000070c3f00000046f64a300024307b1804313043488c56960291101bce40c058
B1[314] <= 640'h810000000000ff2f0f01ff0100003f00ffffc000000000fffffffffffffff8006300000000000000000000001c38760000023d3ad22000301201c113eb99c0e94a101881b99824a8848088
B1[315] <= 640'h1000ff0ff000000fffffffffffff30000000000003fffffff7fe7e0fff07878000000000000000c0000001fffc0000301fd654a400013bc37d0a27c9dd0e08a0ef84121c1c410fa9246
B1[316] <= 640'h3e7ffffffffffffffcf0000000000000000000000000000000007fffffffff7c7f00000000000000040000001f8000000301b9f72ac000278d6d9779924c414b518e1f2b199086e1ae8062
B1[317] <= 640'hffffffc000000000000000000000000000000000001fffff00000000000407ffffffffffffffc00f0000e0000000000000080000000101af4dc2d000174c3ad419936664c382850d0030c7295d9aa040
B1[318] <= 640'h7f3000000000000000000000000001fffffffff00000000000000000000f8fffffffffffffff0ff8e0ff80000000000006103a00009b7f441f09e00139cb7101074b402034b112c48e2d7ea2f4a8683
B1[319] <= 640'h33fffffff000000008000000000000000000000000000000000dfffffffffffffffffef9fffc000000000006000000008b74dcb77de0005639690343250c040498aea29c892760d024602
B1[320] <= 640'hfc000000000000000000000000000000000000000000000000000000180000cffffffffffffffffffffffff16000000000000008f06dbfc18925740009a50ba8a61800124028b192c06b6c240e689982
B1[321] <= 640'h1f1f03fffffffffffffffffffffffffffa00000000000010b86f9dc4c178c0006b8a4e605a8800014876160000626287587c0188
B1[322] <= 640'h7ff07ffffffffffffffffffffffffffffe00000000000180bb2fe8cca8050006140c812c9b17001118c0149610089298ac47200
B1[323] <= 640'h1f803fffffffffffffffffffffffffffff8018f800000444ae547a11ae612dbb9a201185598f46c081515134832468080202860
B1[324] <= 640'he003fffffffffffffffffffffffffffffe00f1000000047a3be29296617afbf602969319b514041a5f420240257563801c0024
B1[325] <= 640'h7ffffffffffffffffffffffffffffffff8000000018484b7c66a2e93fbff528bb07868082cd0080634804b118c27505852
B1[326] <= 640'h3fffffffffffffffffffffffffffff7fffffe0191384c060fc26ed89fa7edb7d53fe294074542212818001ee82810220e5
B1[327] <= 640'hff0e00000000000000000000000000000000000000000000000000000000001fffffffffffffffffffffffff0f00007ffeff9f92f2a91ad50112325fd71208404c8c07222e070d52c180135172a608e7
B1[328] <= 640'h180000000000000000000000000000000000000000000000000000000000003efffffffffffffffd0e7fffff0003ffffffff9d53f79c8e8f69180a59dcc1cd5b9c0d0900054b02d908b62fb30a145806
B1[329] <= 640'h1f1f0007ef000000000000000000008000ffffffffffffffffffffffffffffffffffff80a0807f8fff8001d2db110c555b4cca40fcabda1fc091800e15670623480eca88a8101056
B1[330] <= 640'h1c007ff8ffffff0000000000c1800000000000f4e03f000000000000000000fff8709ffffffffffffff00080ffffff03ff80034ceb0ecee26751c69364016204d80a80021a09000450499d09006c2409
B1[331] <= 640'h8000000000800000000000000000000000000000000000000000000f3ffffeffffffffffffffffffffffffffffffffff7ffe190af60967654987889f744db0610006162013260ee18041383110ec0402
B1[332] <= 640'hfff8008000fe000000000001ffffff7f3ffffc001fff0000000000000000fffcffffffffffffffffffffff5043e70a0bea45178933747b20f1c24a27a24060628dc11c300344d04505
B1[333] <= 640'h80000000000000000000000000000000000000000000000000000000000000000000f807ffff7fffffffffffffffffffffde53ef2c9b78aa47887bda111a48a00a000284b026080001c46d2442004b
B1[334] <= 640'h3e007ffffffffffffffffffffffffff4e8ec415029a35db087331075f0830258390002ca14081046ee4d9264c22
B1[335] <= 640'h3f7e07fffffffffffffffffffffe885294184bf21104a15e936438c15416280641811fd880b1269f01200c5
B1[336] <= 640'h130e1ffffffffffffffffffffb7d406039b6c8801684c260148609020c2048846182021c8232881fb0a7076
B1[337] <= 640'h7fffffffff1ffffffffc7ffe2710cc00c0a26a61aea0a989ac6827560840c20d2904673a0e32d06650
B1[338] <= 640'h1e0000000000000000000000000000000000000000000000000000000000000000000000c3fffffffffffffff9fffff77aa04859509390084b7007a849e2d04230e10690c5f0816ac24844408a8
B1[339] <= 640'h3000000000000000000000000000000000000000000000000000000000000000000000000f3dffffffffffffffffefd602c100b38600741502055a28821400a78213c80008401acdc1d0ca1252
B1[340] <= 640'h6000100fffffffffffffffff924a6dab4b519b7954c88b502a044581a301880c02c000508001c46a0319
B1[341] <= 640'h8000000000000000000000000000000000000000000000000000000000000000000000000000f000011800ffc7ffffffffffa33c49251191024018c34a134c23253029221b61550c8c1924110402002c
B1[342] <= 640'h3000000000000000000000000000000000000000000000000000000000000000000000000000f000039fff3fefefffffffffafc1335691f11c24196702388c13085335c119021148c21e5b510ed01400
B1[343] <= 640'h1c000030000000000000000000000000000000000000000000000000000000000000000000003000039fffffffe03bfffc3e980a29090cbc9c6acd00d04041140048884280c20994043408e09ef1036e
B1[344] <= 640'h600001800000000000000000000000000000000000000000000000000000000000000000000b800231fffffffffff7fef98002898e22c8d544cec9c44081183923a035004430836562d28662a100a3a
B1[345] <= 640'h30000000000000000000000000000000000000000000000000000000000000000c000000000b20003c5fefffff807347ffc0004d0c157708809e9949013880c9c0119b0982180004011036428183b69
B1[346] <= 640'h30000000000000000000000000000000000000000000000000000000000000000fc000000019206600ffe7303fe1c00003c0f3a4085992a8c18a52ce65b810c2041343118202808841281759d4c0946
B1[347] <= 640'h3000000000000000000000000000000000000000000000000000000000000000dfe400e000251ffc6ffff7fff7f0000000706093b3191470c59a029ecd16691d0800010448430500000084050240942
B1[348] <= 640'h300000000000000000000000000000000000000000000000000000000779e0007b68f1980040fcfc413fffffe0fc00000071255001e4806d22871118a30181ef8208100440c10723008820410201121
B1[349] <= 640'h1000000000000000000000000000000000000000000000000000003fbfffff00f8a03fff8e88dffe499fffffc03fe00000c08060002260813129761ceb42d09306a24a044400c0a1108304007321909
B1[350] <= 640'ha000000000000000000000000000000000000000000000000000007ffffffffeb92177f7ff00bfffc99ffc00e003ff80004050e105000015a4b32039ce5a04cc145521800000d180008100266340101
B1[351] <= 640'hc000000000000000000000000000000000000000000000000000007ffffffffe9b0b7fff9f4121fe499fc00000003fff0001884112892817b1f2491a4a9a024024816cc010040004401000400420923
B1[352] <= 640'h180000000000000000000003ff3fffff6470347681b2143c2490000000400180600000a0c04491113ba79db13c8a041008272a80800801302201002180265100
B1[353] <= 640'h3000000000001c002801007ffffffff486c29ffb07273bee40994000000000160782101b0690600d097904288616264e9100950000020060680c12026080100
B1[354] <= 640'h400000000000003000000000000000000000300000003f000007ffffffffff9ff3c93f67e694ff7e109ffc0808000387e790ca50009d34a1a12404e7481c4a60109848c0600002e164081060e800909
B1[355] <= 640'h400000000000003fc40001f8000000000000000ec3f03fff00f7ffffffffffb3e4d36ae7d184b4fa56efff8000000f87c2040a50380db2790b8412d18d9e8446349c52442000248020018004c94018d
B1[356] <= 640'h4000ff8000007ffe00000000fff07fffffffffffffffffd73c8018cf99e2b0fc92d6c000000fffdfcb0044824c48884fb1d45a30c60d120610221800102080000032000d0a00024
B1[357] <= 640'h400000000000000000004000001f0003c003f7e73ff0ffffffffffffffffffcb1010b8cf312360fc920c00000013ffffc90e612a6448610b181c8074949800001210842000348080203000068440100
B1[358] <= 640'h400000000000000000000000003000007003fffffff1fff3e3ffffffffffffdc1076b84e3194a0fa941c800c0111ffffc98142282c00211009c18d86d52644b02208488020022441300300262440980
B1[359] <= 640'h400000000000000000006606080000000ff00fffff81ffffffffffffffffffd93866f0106886f4790489903ff811ffffe98261449c08ca9a2db04d4911a423b400408000000260080f0100002401800
B1[360] <= 640'h7e000000000000000000000000000001f0001c0011ffffffffffffffffffcc1809f118a02e787c4317807fea12ffffec4081a25e8e400da813d810878160020841800000000004000000000521800
B1[361] <= 640'hc383c4000000000000000000000000000000000007ffffffffffffffffffffea6d01195c8087e23327278fffc270fffff6f30662509d1005b843808406b0600200a2400006000084800040000026c00
B1[362] <= 640'h8701000000000000000000000000010000000007fffffffffffffffffffffff53337801c4846e2703726dfffc840fffff1195802710a30682dd308a4930403082100000003000080400048403020000
B1[363] <= 640'h8c0006000000000000000000000000040000001fffffeffffffffffffffffff9a38f4ab8c1129079166c1fffc040fffff469a3a23a8418251414007917082498000004800100409e400000000240200
B1[364] <= 640'h98003180000000000000000000000000400008300001e3fffffffffffffffffcc11f0384c50182e903753fffc86147fffe0c86c611402405288603c1810c0c40042000080000200e000008000440000
B1[365] <= 640'h20000040000000000000000000000204000003c00003fffffffffffffffffe640d027f906140924c1f672fffc44987fffccef4c220442453a00a43630b2208800400004c01000003000000000000000
B1[366] <= 640'he000007fc000000000000000000000070000004803cffffffffffffffffffe98b46fff3300c982404b4c9fffc04980f9fa4b101226406401a4814739007261c00000000000020000020000040000200
B1[367] <= 640'h1000000177f00000000000000000001040000000019fbfffffffffb7fffffffc9d4441041080b04c40a148ffff26306e1fa4192404a52352084bd8cbd104c244c080000020402c000100000000860800
B1[368] <= 640'h42e600000000000000000005100000001061ffffffffff8d7dfffd596c5aa1816c4801624e8827ff613605017a0490420e35207a5a410ade810104040c00901404400014400000000001840
B1[369] <= 640'h5580000000000000000407800000000068cfffffffe705fdfbf9d02a5d00a4108c4120195877ff03202900700b1c810500174e0260004a104215100400004e00000000000000000823800
B1[370] <= 640'h78000bc0420000000000008060005c001e20077ffffffc323187b9c800d854680880c012019558fff8e024a602149810c220015810b6882a59a2424480001404100000000800000000002000
B1[371] <= 640'h760004df8000000000000023a3e007f3c0004f7ffffdfc212a84a9884dd1e0b8840140104494d3fff8311e24954201008209b1cd11e49c7441820041c2011ce8100000002a04000000060000
B1[372] <= 640'hf0000137f100000000000d00afff880ff0ffffffffffca05b048de44c88f2e48a0904402c94507ffc3b2320000000100408e0841140321071242003200108e0000000002210000000040000
B1[373] <= 640'h378000008c40000000000000203ff1f0080fffffffff8087f44d8d0040093240c0100920091c4fffc396600004720001082619081202243112dbc2800006480000000000406000000000000
B1[374] <= 640'he080000047460000000800000003ffff80ffffffffe809674c9000122d1a0214004882003347ffc19c0c4c14220010440021909866745389621e0180000000800000003007000000600000
B1[375] <= 640'h380f80000238800000000000000000fffffffcffffc84204448000000dfacc0013009604844400c016990008831000040c048109248400d1038c031000002040000010000002000000000d
B1[376] <= 640'he30fe00003088000010000000000000fff7ffffffec7257388040032ea44d8083020004826423e02a1a121800004e004898c8482508096023a8000000018c900000500000000000000000
B1[377] <= 640'h101ffff000003880008000100008003fc007fffff0cd9224c1020630116880300021046d26461002e32001040002220400c0809024c11f120000000000888800000000000000000000000
B1[378] <= 640'h3f007c00039b8018000300010000f0ffffffdf8489862c01406504206212050101224e0600801254000000080020c4f6400045b4f04020060da0008001c00000000000000000000000
B1[379] <= 640'h60000961fc0003c00c0001c0313e0007ffffffe08d99162486b0124404646424802330982400004966000000100080000200b9ef00881905d20020000000000000000000000000000000
B1[380] <= 640'h3c0001fee0fe0020880000c0ffffd80fffffff644cc1260400109950004864248030124c4c00004520009801000000000071008040005804200000001a08000000000000000000000000
B1[381] <= 640'h304001fff01c00114000089fff1001ffffdcf888481bb001084e010c11910c0884013105b00402c2400d001800000000000400070781225000002000400000000000000000000000000
B1[382] <= 640'h80ff80beffff80000000003ffffffffce0effd4cf1b810160418358f140c404066411806381900000000000000000000000002080000210c0000000000000000000000000000000000
B1[383] <= 640'h603ff9003ffffc000001001ffffffbff061fffc6f0a802209618308a14112042208010000112c30a070000000000000000008902005024020000000000000000000000000000000000
B1[384] <= 640'h18003fe0805fffff00019487fffe07ffc103f6f0c080620c0b1b861c8e13a002008010001800332e00000000000000000000518080100c000000000000000000000000000000000000
B1[385] <= 640'hc0003fffc000ff0f8000011fbf807ff5ffeca7c48a4e106444382242600e000204000001800180810000000000000000000204a908002020620000000000000000000000000000000
B1[386] <= 640'h60000001cffff07ff000004fdffffffedfffa780886140048cb02a3002020202000000000419000000000000000000000000000044260490320000000000000000000000000000000
B1[387] <= 640'h3c000000003cfc07fffff81173fffffffff17d528f0108070822603624220000000040a00000000008000000000000000000000000160000200000000000000000000000000000000
B1[388] <= 640'h7000000000009c037f77fc6d7fffffffe07030b87816027940b1236404240500020c00000010040a0000000000000000001000000000004200000000000000000000000000000000
B1[389] <= 640'h1f0000f0cef000c09fff7f13ffffffff0f80019810240111a11162400004040000001047781818580000000000000000000000000000000000000000000000000000000000000000
B1[390] <= 640'hfc000000f7fe007180cb382fffdff002000000000002cbfd0987c400000000000066040080610000000000000000000004800000000000000000000000000000000000000000000
B1[391] <= 640'h33000000000180000004df23ff8fc030008400000000a1589e248000000000000040000040000000000000000000000002200000400000000000000000000000000000000000000
B1[392] <= 640'hc00000000000111003e67c0ebffc003e80400000000016002000c06000000000080000000000000000000000000000000000000000000000000000000000000000000000000000
B1[393] <= 640'h70000021c0f000ffe03eff2d306001ff8040000000000092e0349c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[394] <= 640'h1f00057fe17fe007fbf00fc41ffb0100000000000000001e21200c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[395] <= 640'h7e00000003ff5f801f000bc000000000000000c000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[396] <= 640'h1fc0000000000fef002fa6f0000007f00c0000c030240000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[397] <= 640'he10000000160067fe0079f803e037fc0c8000c030100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[398] <= 640'h3000000003ff00007f8027706f03fff640000fb000921c0000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000
B1[399] <= 640'h600080060fcfc0001fc88877f03ffff60002030005dbf0000000000000000000000000000000000000000000000000fc3000000000000000000000000000000000000000000
B1[400] <= 640'h1c00000000003fc0009fe7fc002ff2060000010049fff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[401] <= 640'h60000000000007fff006ffe000fc0000000c13039fff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[402] <= 640'h6000000000000007f8000070000f0000000c120080cf8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[403] <= 640'h183000000000000000fc00fc0003c0000000000080040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[404] <= 640'hc001f000effff000003fe7e000180000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[405] <= 640'h100030038000e7ff400003f800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[406] <= 640'he0000000000007fff80001e00000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[407] <= 640'h3c0000000000000001c000fc0000000000000000060000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000
B1[408] <= 640'he80000000000000000100bf0000000000000000040000000000000000000000000000000000000000000000000000000001900000000000000000000000000000000000
B1[409] <= 640'h30800003c387fe00000003fc000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[410] <= 640'hc000003e0000f98e0000007000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[411] <= 640'h600000000000000ecce0001c0000000001c000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000
B1[412] <= 640'h18000000000000000000c0fe3800000000cc00800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[413] <= 640'h70000000000000000000001c8000000002300e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[414] <= 640'h18000000017907000000000600000000004601c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[415] <= 640'hc004f9072000380407f80010000000000310000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[416] <= 640'h1000e001000000000000000e783000000062000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000
B1[417] <= 640'hc0000000000000000000001840000000013c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[418] <= 640'h30000000000000000000000000000000006980600000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000
B1[419] <= 640'hf00000001ff83800000066100000000000920180000000000000000000000000000000000000000000000380000000000000000000000000000000000000000000
B1[420] <= 640'h3003fec3fc0000000000000400000000002e8070000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[421] <= 640'h1800f000000000000000000600000000000b801c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[422] <= 640'hc00000000000000000000008000000000027407000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[423] <= 640'h18000000000000000c000002000000000008180800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[424] <= 640'h7000000001c000000000000800000000003020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[425] <= 640'h1c000000000000000000000700000000000c0c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[426] <= 640'h6000000000000000000000080000000000183000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[427] <= 640'h30000000000000000000000007ffc00000071000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[428] <= 640'hc0000000000000000000000000001e1e000e000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[429] <= 640'h38000070000000000000000000001e010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[430] <= 640'he00003880000000000000000000003c8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[431] <= 640'h30000000000000000800e0000001fc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[432] <= 640'hc000000000000000000000079fc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[433] <= 640'h700000000000000000000005ff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[434] <= 640'hc00000000000000000003f8fc00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000
B1[435] <= 640'h38000fffcc000000001ff800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[436] <= 640'hf800c00000000000ff00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000
B1[437] <= 640'h38000000000001ff8000000000000000000000000000000000000000000000000000000380000000000000000000000000000000000000000000000000
B1[438] <= 640'he00000000007f800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[439] <= 640'h300000000fff8000000000000000000ffc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[440] <= 640'hc000013fc000000000000000000000ff7ee0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[441] <= 640'h3800fff40000000000000000000000ffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[442] <= 640'hf3f800000000000000000000000007fffc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[443] <= 640'h3fe000000000000000000000000007fffc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B1[444] <= 640'h7fe000000000000000000000000000000000000000000000000000006000000000000000000000000000000000
B1[445] <= 640'h12000000000000000000000000000000000000000000000000000000e000000000000000000000000000000000
B1[446] <= 640'h13000000000000000000000000000000000
B1[447] <= 640'h1f00ff800000000000000000000000000000000
B1[448] <= 640'h803860c00000000000000000000000000000000
B1[449] <= 640'h180000000000000000000400000000001808180000000000000000000000000000000000
B1[450] <= 640'h2000000000000000000000000000000000c000000000000000000030000000000067c300000000000000000000000000000000000
B1[451] <= 640'h2000000000000000000000000000000000600000000000000000001800000000601e3e00000000000000000000000000000000000
B1[452] <= 640'h8000080000000000000000000000000000000000000000000000000000000000000
B1[453] <= 640'h3f0000c0000000000000000000000000000000000000000000000000000000000000
B1[454] <= 640'h220000000000000000000000000000000000000000c7c0000000000000fc11000000000000000000000000000000000000000000000000
B1[455] <= 640'h20000000000000000000000000000000000000000013fc1018007f3bc00130000000000000000000000000000000000000000000000000
B1[456] <= 640'h6000000000000000000000000000000000010000000e3ff80ff001809fe2c000000000000000000000000000000000000000000000000
B1[457] <= 640'h7000300000000008000000f80000600003ffee88ff90328000000000000000000000000000000000000000000000000
B1[458] <= 640'hf0107e3fffc04000000000180000e603ffc00bf27f70328800000000000000000000000000000000000000000000000
B1[459] <= 640'h3ff800000000000000000ffffe00000c880c3e38000000000000000000000000000000000000000000000000
B1[460] <= 640'h88020c060006c000010080000000000000000000000000000000000000000000000
B1[461] <= 640'h3700000ff80fe000000780000000000000000000000000000000000000000000000
B1[462] <= 640'he0003f00c07e00000097e000000000000000000000000000000000000000000000
B1[463] <= 640'h33f00000000000000000007000fe33003e00000c104380000000000000000000000000000000000000000000
B1[464] <= 640'h2600900000000000000000000000000001ff83f2e0000f80000c10c220000000000000000000000000000000000000000000
B1[465] <= 640'h400000000000000000000000000000001ff07e0000007f8001851cc18040000000004000001800000000000000000000000
B1[466] <= 640'hd00c000000000000000000000000000000000000000000000000000000000000000000000000000000000007000831c422000000000004000001000000000000000000000000
B1[467] <= 640'h7fff0fe001000000000000000000000000000000000000000013800000000000000000000000000000000000000074bc33fff000000000000000000000000000000000000000000
B1[468] <= 640'h23fffff76d60ff800000000000000000000000000000000000004010e000000000000000000000003f8c000000000000e0410a008e00000000000000000000000000000c00000000000
B1[469] <= 640'h3ffffffe37c38b7000000000000000000000000000000000000080004f8000000000000000000000002000000000000000f47a1c000c0000000000000000000000007c01c00000000000
B1[470] <= 640'hf3fff80015430f8000000000000000000000000000000000000000003b600000000000000000000000ff0000000000000004b07400038000000040000002010000780400000000000000
B1[471] <= 640'h1ffff00000194e00000000000000000000000000000000000000000000788e0000000000000000000003fef0000000080000000fe00180c000000000000287018007c00d30680007e00400
B1[472] <= 640'h7f00000003f840000000197080000000000000000000000000000000000000000000703f0000000000000000000007fff880000044000000000fc00088000038600008169ff390000f0ed40079e80000
B1[473] <= 640'hff800000c600000000001900c00000000000000000000000000000000000000000007018000000000000000000000300f80000004000000000003e006b000018e0000000180f500009fffe007b400000
B1[474] <= 640'h3c107ff440000000000190040000000000000000000000000000000000000000000701c00000000000000000000071fc000000000000000000001fe6300000000000007f00f88000800fe0010000000
B1[475] <= 640'hffffff440000000000110000000000000000000000000000000000000000000000308c0000000000000000000007fe000018000000000000000001e0c000000001e0c0000f080e1805270000000000
B1[476] <= 640'h6ffffc41c000000002f00000000000000000000000000000000000000000000003efc1c0001f000000000000003f800000900000000000000000000000000817e00400001c007fe3b9f0000000000
B1[477] <= 640'hfffffffc640c000000006c00000000000000000000000000000000000000000060001fc036000208000000000000000000000000000000000000000000000001a14000c060016fff1c0fce00f8000000
B1[478] <= 640'h1fffffb0240000000006c0000000000000000000000000000000000000000000600007c004000208000000000000000000000000000000000000000000000000c1400074000b0fc7e0000000f90e000f
B1[479] <= 640'hfffffff004800000000fc18c0000000000000000000000000000000000000000200000000000020c000000000000000000000000000000000000000000000000007fe0f0c7ff8ffc0000000067c10400
end
always @(posedge vga_clk) begin
B2[0] <= 640'hffffffffc7fcfff77ff0000e00000102000001000000000000000000000000000000000000000400000c00000000000000000000000000000000000000000000000000000800000003c0000000000000
B2[1] <= 640'hffffffffc73ffffffffe00ff00000060000001000000000000000000000000000000000000010000008000000000000000000000000000000000000000000000000000000000000001c0000000000000
B2[2] <= 640'hffffffffbf1fffffffce00ff00c000e000000100000000000000000000000000000000000000000000800000000000000000000000000000000000000000000000000000010000000100008000000000
B2[3] <= 640'hffffffff3ff8ffffe78e02bf008000e000800100000000000000000000000000000000000000800000000000000000000000000000000000000000000000000000000008804200000100000000000000
B2[4] <= 640'hffffffff3ff87fffefce033f800003670000010000000000000000000000000000000000008c180000180000000000000000000000000000000000000000000000000018004200000000000001000000
B2[5] <= 640'hffffffffff3ffffffffe027f830007070000000000000000000000000000000000000000000c080000000000000000000000000000000000000000000000000000000000004200c00080000100000000
B2[6] <= 640'hffffffffffffffffffff00ff1fce076700300001008000000000000000000000000000000000000020018000000000000000000000000000000000000000000000000000006600000001000080000000
B2[7] <= 640'hffffffffcffffeffff3f007f87efc0e600300001008000000000000000000000000000000071060060608000000000000000000000000000000000000000000000010100036600008001010001000000
B2[8] <= 640'hfffffffffff9fffffffe18ff83f9c7038f3c831e0000000000000000000000000000000000000066002080000000000000000000000000000000000000000000000000012010c600c000048000000000
B2[9] <= 640'hfffffffffffffffffffe02ff339fff0f0100001e00000000000000000000000000000000000000000001800000000000000000000000000000000000000000000000000000100100c000040000000000
B2[10] <= 640'hffffffffffffffffffff03ff7eff7eff21801c0f00000000000000000000000000000000180000000c03000000000000000000000000000000000000000000000000000880103100c306602000000000
B2[11] <= 640'hffffffffdffffffffdff03ff76ff7eff21000c8700000000000000000000000000000000000100998c00000000000000000000000000000000000000000000000000008c0e601100e707603000000000
B2[12] <= 640'hfffffffffffbfffffdff83fff7ffffff863883030000000000000000000000000000000000010099843800000000000000000000000000000000000000000000000000840ce0c7007c07620000000000
B2[13] <= 640'hffffffffff7fffffffff83fffffff3ff8438c3410000000000000000000000000000000080010099001cc0000000000000000000000000000000000000000000000000c01ce0c7fff807660000000000
B2[14] <= 640'hffffffffffffffffffff83fffffffbffc0fcc7f30000000000000000000000000000000104070066010ec00000000000000000000000000000000000000000000000006060e307fff807c60008000000
B2[15] <= 640'hffffffffffffffffffffcffff9fffbfbf3f33fff008800000000000000000000000000010e073c6673c0c000000000000000000000000000000000000000000400c00070e1e313ffec07848808800000
B2[16] <= 640'hffffffffffffffffffeffffffffffffefc1e030481000c0000000000000000000000000f67d19ecf6600600060010000c000000000800000000000000000000000000807c366f37b6099804800000000
B2[17] <= 640'hffffffffffffffffffffffffffffff66ffff0380003c100000000000000000000000001f6799dfce6700600000000000e0000000000000000000000000000000000080f0c366e300fc99000000000000
B2[18] <= 640'hffffffffffffffffffffffffffffffc7c3ff3ffc3f7c700000000000000000000000003f7fb8ef9e9900600000000000008000000000000000000000000000000000c0008166c7338c00000000000000
B2[19] <= 640'hffffffffffffffffffffffffffffffe7e1ff3ffcffc3e0000000000000000000000000ff7ff9ffc79900600010000000008000060000000000000000000000000000c00f0000ce7f8024004000800000
B2[20] <= 640'hfffffffffffffffffffffffffffffffffc7f7ffcf6c7c0000000000000000000000000fc1bf9ffc39900000030000000dc000002c0000000000000000000000000009cf00000df01fb64c04000000000
B2[21] <= 640'hfffffffffffffffffffffffffffffffffc79fffee73e840000000000000000000000003e99fb7ff39fff900010000000de000000c0000000000000000000000000001cf81899ff7b7160c00000000000
B2[22] <= 640'hffffffffffffffffffffffffffffffdffffbfffffffef00000000000000000000000007fffffff7fffff900000000000c40000000000000000000000000000000000041f3c99ffff0000004000000000
B2[23] <= 640'hfffffffffffffffffffffffffffffffffffbffff67fcf0800000000000000000000001fffffdff7f7fff908011000000c0000000000000000000000000000000000003f83c997133ce03264900000000
B2[24] <= 640'hffffffffffffffffffffffffffffffffdeffff7ffffff1808000000000000000000004ff3f7fffff977e0300ee000166f080000000000000000000000000000000000000c78efffe1806000000010000
B2[25] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffe000000000000000000000006ff7ffffffff67f3000e4000066f3c0000000000000000000000000000000000000f7cff1ff38000000c0000000
B2[26] <= 640'hfffffffffffffffffffffffffffffffffefffffffffffe610000000000000000000006fffffffffff67ffc80f00000467300000000000000000000000000000000002000fcff71f71880000080000000
B2[27] <= 640'hfffffffffffffffffffffffffffffffffefffffffffffe600000000000000000000007ffffffffffffff1e00f0c000077300000000000000000000000000000000003003fef3ffff0080000000600000
B2[28] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffcc0000000000000000000003fffffffffffffffe00f0c0180773000000000000000000000000000000000031077f73fffe8001708100600000
B2[29] <= 640'hffffffffffffffffffffffffffffffffffffffffffffff9c8000000000000000000001fffffffffffffffc017800fc8ff9c000000000000000000000000000000001300f3ff3defec000308100000000
B2[30] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffdc0000000000000000000019fffffffffffffff3017fc0ff9effc000000000000000000000000000000001301feffffefec020310000000000
B2[31] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffff1000000000000000000003bfffffffffffffff3307fffff9efe0000000000000000000000000000000000301fe3ffffff08673100c0990000
B2[32] <= 640'he7bffffffffffffffffffffffffffffffffffffffffffdc08010000000000000000e3fffffffffffffffbfffb88f03fffb0000008000180004000000000000000000033f7de6c7e20cfe9c0010000000
B2[33] <= 640'hffffffffffffffffffffffffffffffffffffffffffffff9e00000000000000001cff7ffffffffffffffffeff07cf73fffd0000008400000000000000000000000000033f7de77fe6833f080096000000
B2[34] <= 640'h3ffffffffffffffffffefffffffffffffffffffffffffffe00000000000000001e3f7fffffffffffffffbfffe3cefffffd40000004c08100000000000000000000001efb7fe77fff83879cc092000000
B2[35] <= 640'hff7ffffffffffffffffc9fffff3ffffffffffffffffffffc0000000000000000c7337ffffffffffffffffffef1fffffffc61000000c08100900000000000000000001eff7ffffffe23f3ff0092000000
B2[36] <= 640'hff7fffffffffffffffff9ffffffbfffffffffffffffffff0c000000000000000c3fffffffffffffffffffefeffffffffff600000000000001100000000000000000003ffcd3cfffc30fc800092000000
B2[37] <= 640'he7ffffffffffffffffe3ff7ffff3fffffffffffffffffff7e000000000000000fcffffffffffffffffffffffffff0fffff4000000003000001000000000000000000439fcd3cf398383f110010000000
B2[38] <= 640'h3ffffffffffffffffe166ffff3fbfffffffffffffffffffe0000000000000007cffffffffffffffffff3fffffffdfffff4000000002000000000000000000000000009fcf9df399083ffb0030000000
B2[39] <= 640'h18ffffffffffffffffe066effefbffffffffffffffffffff0380800000000000fffffffffffffffffffefbffcffffffffec48000e31800000400000000000001000000ffcf9b7f9980ff010032e0c180
B2[40] <= 640'h3bfffbffffffffffff8019bb3f99efffffffffffffffffff7f180000000000007fffffffffffffffffffffffffffbbfffe8020c03c67811800001080000000000000010f3fc7f967000e80c1e30f9c00
B2[41] <= 640'h3bffffffffffffff7f8098bb07098fffffffffffffffffffff180000000000007fffffffffffffffffffffffffffffffffc070c0c16700100000000000000000000001be3f0ff067000e0000e1048800
B2[42] <= 640'h3bfffffffffffe9f7f00009c03067ffffffffffffffffffef818000000000000ffffffffffffffffffffffffffffffffffe0f1e1e06700000000010000000000000000ff3f0f706600871000e0c08000
B2[43] <= 640'h3bfffffffffffefff800009c3066fbfffffffffffffffffff000000000000000ffffffffffffffffffffffffffffffffffe0f0637c663c0007000000000000000000003f3f0ff86600cf1810e0c00000
B2[44] <= 640'h3bffffffff3ffffffc00000cc06627ffffffffffffffffffc300000000000001fffffffffffffffffffffffffffffffffff080373c663c0000000000420000000000003f00c1fc60008f0000fc800000
B2[45] <= 640'h3bffffffbfffffe61c000000830003ffffffffffffffffffc700000000000001ffffffffffffffffffffffffffffffffffe0803fc76600000000000000000000000000ff00e0fe60000e0000fe000000
B2[46] <= 640'h3bffffff88feff660c0000200300807ffffffffffffffffffe00000000000001ffffffffffffffffffffffffffffffffffe0cc31e366000000000000000000000800003800e39e60001c0000fe1c0000
B2[47] <= 640'hfffffffffc3ffe66c00000203c800e3ffffffffffffffffffe00000000000000fffffffffffffffffffffffffffffffffbe08e207826008000000000000000000300000700078c60001c00010c3c0000
B2[48] <= 640'hffffffffffc4fe8cf8800000008400ff7fffffffffffffffff00880000002001ffffffffffffffffffffffffffff7ffffffe8c2002a83000000000000000081000810007183c77c00081030008030000
B2[49] <= 640'hff7fffffffc03f873e100000000000ff6fffffffffffffffff00800000000018ffffffffffffffffffffffffffffffffc3ff80000001200000000000000080000018000381f077000001010000000000
B2[50] <= 640'h7f7efffffff0ff071f1000000000013fffffffffffffffffffc0800000000018ffffffffff7fffffffffffffffffffffffff808000010000000000000000810100000003818104080001e00000000000
B2[51] <= 640'h3e67fffffff1f938f08000004000009effffffffffffffffff808000000000c3fffffffffffffffffffffffffffffffffffe8000803800000000000000000000008100033881040c0020e00000000000
B2[52] <= 640'h3ee7ffffff31f931f08000000000008ebdffffffffffffffff000000000000c3fffffffffffffffffffffffffffffffefffe800080380000000000000000180000030003380004000022100000000000
B2[53] <= 640'h3fe7ffffff1339c1e0000000000000033ffffffffffffffffc0000000000000effffffffffdfffffffffffffffffffffffff603000c30000000000000000000080060003631c04000022180000000000
B2[54] <= 640'hff7fffffffcf9981c3000000000000312ffffffffffffffffc0000000000012efffffffffffffffffffffffffffffffffffe701000800000000000000000000000000003630020800022000000000000
B2[55] <= 640'hef7effffffcf981ce08000000080013147ff67ffffffffffff80000000003167ffffffffffffffffffffffffffff7ffffffc780c000c0000000000000000000004400007340160000022003000000000
B2[56] <= 640'hc378dfffff3f6e0060000000c00000869ffffefffffffffffcc0000000000c0effffffff3fdfffffffffffffffffffffffe3000f600080000000000000000000000020023880e3000001000000000000
B2[57] <= 640'h3ce3ffffffff6e00200000000000000389ffffffffffffffc00000000000048fffffffff7ffffffffffffffffffffffffff000002000000000000000000000000100013e000162000001000000000000
B2[58] <= 640'h3ce7ffffffff9801000000030000002081ff7ffffffffffec0000000000001cfffffffe7ffffffffffffffffffff3efffff8c0000001000000000000000000000000033f000000000000000000000000
B2[59] <= 640'h3ccf7fffffff9801800000000000000001e7f7ffffffffff3c000000000001fffffffffefeffffffffffffffffffff7ffff8c0000001000000000000000000000000073f830000000000000000000000
B2[60] <= 640'h1f7fffffff980098000000010000070067e7ffffffffff3c000000000001fffffffffedfffffffffffffffffffff7ffff818030000000c00000000000000000000823e810000000000000000000000
B2[61] <= 640'h813c7ffffffffd001800000000000000001fe7ffefffffffc00000000000017fffffffe7dfffffffffffffffffffe7ffffc03cc30000820c00000000000000000000e03e000000000000000000000000
B2[62] <= 640'h3cffffffffee01100000000000000002997377ffffffff800000000000077fffffffffffffffffffffffffffffefffffe078800000a8a800000000000000000000213f000000000000000000000000
B2[63] <= 640'h1cffffffffffe7c10000000000000000009831737effffff00000000000087f3fffffffffeffffffffffffffffff6ffffff0c000080018c00000000000000000080023ffc01e06000002008000000000
B2[64] <= 640'hdffeffffffff7fc00000000018000000000001eeeffffffef800000000003f3fffffffff4fffffffffffffffffff3ffffffc010000108003000000000000000100816f78308130800000000000000000
B2[65] <= 640'hffffffffffffffc0f00000000000000000000006fffffffecc00000000003ff9fffffffffdfffffffffffffffffebbffffff000fc0000000000000000000000f8088f678710000000000000000000000
B2[66] <= 640'hffffffffffffffe4000000000000000000000000ffffffff0000000000007ff1fffffffffffffffffffffffffffedbbfffff000fc0000000000000000000001f80987ff1711c00000000000000000000
B2[67] <= 640'hfffffffffffffee6000000000000000000000006fffffffd8000000000007fc7ffffffffffffffffffffffffffff9fbffffe000f00000000000000000000001fc09c0fe3a00b04000000000000000000
B2[68] <= 640'hffffffffffffff768000000000000000000000273ffffffdc000000000007fffffffffffffffffffffffffffffff8ffffffe000307300000000000000000001ff09ce8a0000300000000000000000000
B2[69] <= 640'hfeffffffffffc7760000000000000000000000223fffffffc000000000007fffffffffffffffffffffffffffffff8dffffff000203100000000000000000003fff9f9960000100000000000000000000
B2[70] <= 640'hffffffffffffcf76000000000000000000000022ffffffffc00000000001ffffffffffffffffffffffffffffffff91bfffff0000001000000000000000000003ff9f1b70800000000000000000000000
B2[71] <= 640'hfffeffffffff3e72000000000000000000000076ffffffff840000000001fffffffffffffffffffffffffefffffff0beeefe0000000000060000000000040003ff9fd878ce0001010000000000000000
B2[72] <= 640'hfdff7fffffffff0c00000000000000000100060ef3ffffff800000000101ffffffffffffffffffffffffffffffff8e63fffe0080c00000000000000000000023cfff84038c000c000400000000000000
B2[73] <= 640'hfffffffffffffcc0c000000000000000200000037fffffff800000000001fffffffffffffffffffffffffeffffff899ffeff0000800018200000000000000023cfff8fb72a8000000000000000000000
B2[74] <= 640'hffffffffffff7cc00000000000000000000000137fffffff800000000007fffffffffffffffffffffffffe7ffffc119e1c7b800004000c600000ff0000000001fcffffff73ef00002000000000000000
B2[75] <= 640'hfffffffffffff81c000000000000000000000103ffffffff00000000000fffffffffffffffffffffffffe37ffffc11be3e7380000000032000003f0000000000f9fffffffbff70000000000000000000
B2[76] <= 640'hffffffffffffc0180000000000000000c0000107ffffffff000000000007fffffffffffffffffffffffff37fffff80f3fff7c0002000030300007ffc000000007fffffffffff80000400000000000000
B2[77] <= 640'hffff7fffffffc1c000000000000000000000000fffffffff800000000003ffffffffffffffffffffffff783fffff887323efc00030003c170081fffc00000000ffffffffffff80008400000000000000
B2[78] <= 640'hffffffffffffe0c000000000000000000000000fffffffff800000000003fffffffffffcfffffffffffff80f7fff013f3ffee00000003c700081fffe00000004ffffffffffff00008000000000000000
B2[79] <= 640'hfffffffffffff800000000000000000080000037f3ffffff800000000003ffffffffffffffffffffffffc00ff3fc011f3ffee0040000c1f0101efffe000f0000ffffffffffff00000300000000000000
B2[80] <= 640'hffff7ffffff73c80000000008000000000000046c7ff7fff800000000003ffffffffffffe3fffffffff9e63bffe60063837f78400000393e01f3ffffc06680037fffffffffff08001c09000000000000
B2[81] <= 640'hfffffffffffff00800000000000000000000000406fffffec0000000000fffffffff7fffe1ffffffffffee39ffc0183889fff0000000383e017fffffc8e60001ffffffffffff00000089000000000000
B2[82] <= 640'hffffffffffffc01800000000000000000000000000ffffffe0000000000ffffffffffffe1c1ffffffffffd3dffc0183e19ffe300200038e0187fffff8cdf8000ffffffffffff00000098000000000000
B2[83] <= 640'hffffffffffffc00000000000200000008000000100fffffff0000000000fffffffffffe61ccfffffffffd93dffc007e31bfff780000000c0187ffffffc99ff28fffffffffffe80800199000000000000
B2[84] <= 640'hfffffffffff7fc8000000000200000000000000001ffffffe0000000000ffffffff79fe68cfffffffffff93fff1803e323ffff808c0000c0017ffffffc99ffeffffffffffffec1801f1f000000000000
B2[85] <= 640'hfffffffffff73c00000000004000000000000000000fbfffe0000000000ffffffff7fffece7fffffffeff19fff1cc37ee77ffe008c8000c001fffffffeffffffffffffffffffe1801a1f000000000000
B2[86] <= 640'hffffffffffff3c00c0000000000000000000000000061fffe00000000007fffffff7ffffff7ffffffffee3cfff9df7fffffffe007080043801fffffffffffffffffffffffffffb840ffd000000000000
B2[87] <= 640'hfffffffffbfe0080000000009c0000000000000000001f7fe00000000003ffffff377fff7ffffffffffee3cfffdffcfffeffff62711c043c007ffffffffffffffffffffffffff9f007f8000000000000
B2[88] <= 640'hff7fffffffccbf8100000000f000000000000000008efeffc0000000000ffffffefbffffcffffffffefff97efffffffffffffff00900000003bffffffffffffffffffff3fffffe99e7ff000000000000
B2[89] <= 640'hffffffffffdcb38000000000100000000000000000047fffe000000000dffffffffbffffffffffffffffffffffffffffffffff3fd902008c03fffffffffffffffffffffffffffff8ffff000000000000
B2[90] <= 640'hfffffffffffe92000000000038000000000000000000fffff0000000001ffffff7f9ffffffffffff7ffffffffffffffffffffff8fdff03fe0ffffffffffffffffffffffffffffffeffff000000000000
B2[91] <= 640'hfffffffffefe820000000070f8000000000000000001fffffc000000003ffffffffffffffffffff39ffff6fffffffffffffffff03ffff3de0efffffffffffffffffffffefffffffffffe000000000000
B2[92] <= 640'hfffffffffee0be7800000071fc0000000000000000637ffffc00000000fffffffeff1fffffffff71ffff7fff7fffffffffffff077efef3debeffffffffffffffffffffffffffffffffff800000000000
B2[93] <= 640'hfffffffff7e0bef000000070fe0000000000000004f7fffee500000000e7ffffc1ff0fffffffff79ffffffffffffffffffffff87fefef1f89fffffffffffffffffffffffffffffffffff800000000000
B2[94] <= 640'hffffffffffe1b7c000000179ff000000008e000006fffffff00000000017ffffffffcfffffffffe03ffffffffffffffffffffff8effff171cfffffffffffffffffffffffffffffffffff800000000000
B2[95] <= 640'hbffffffffef3b7e08000007bfe46000000fe8000047fff7f30000000023bffffffe7ffffffffffe07f7fffffffffffffffffff1f47ff71718fffffffffffff7ffffffffbefffffffffff800000000000
B2[96] <= 640'hfe7fffffe6cffefc000000fbfee00000833fe000003ffff9300000000007fffffffeffefffffffdb1fffffffffffffffffffffe1dfdeff7086ffffffffef73fffffffff731fff7ffffffa00000000000
B2[97] <= 640'hfffffffff7efffff000000f9ffc000003cff600000bffffd700000000006f8fffeffffffffffffe01f7ffffffffffffffffffbf1ffcfff6006fffffffffefffffffffff008ffffffffff800000000000
B2[98] <= 640'hffffffffffffcff3800001ffffcf00003fff000011fffffce00000000008fffffefffffffffffec11f3ffffffffff1fffffff99cffcfffc00efffffffffccffffffffff08c7fffffffff810000000000
B2[99] <= 640'hffffffff99ffeff3000007fffffe00800ffc00001ffffffc00000000001cffffe7ffffffffffffdf1f07efffffff0070fffff18ce3df3fc00efffffffffee7fffffffef0803ffdffffff610000000000
B2[100] <= 640'hffffffff9ff9fffb00001ffffff8003b87fe00010ffffffc000000000007fffffffffffffffffff807c3effffffc003003fff380c03c3f800efffffffffff37ffffffff0003df97ffffff00000000000
B2[101] <= 640'hffffffffbff9ff7e00001ffffff8003fffff0000cffffefe000000000007ffffffffffffffffff980710efe7fff8000007ffff80f838f8180ffffffffffff37fffffffc00038717ffffff80000000000
B2[102] <= 640'hffffffffeff9fe7a000003fffff8003fffff0000fffffee4000000000007ffffffffffffffffff190600edc3ffc000000fffff007c00f8981ffffffffffffffffffffd000000607fffffcc0000000000
B2[103] <= 640'hffffffffc6fb8ef3000003fffff8001eff7c0004fffffee000000000003fffffffffffffffffdff96603e00099c0000004ffff3818033f881fbfffffffffdffffffff0000000647fffff8e0000000000
B2[104] <= 640'hffffffffffff9970800003fffffe018eefd80019fffffe0000000000097ffffffffef1ffffffe7c1630001806c80000000fffe00c0000d804dffffffffffffffffff00800000f0cfffffb00000000000
B2[105] <= 640'hfffffffc7fff8920800007fffff0000eefd80019ffffff7800000001007fffffffff07ffffffe7ff0700010041000000007fff0000000fc0edfffffffffffffffffc00000000f1ffffff100000000000
B2[106] <= 640'hffffffff7fffe620000007ffffe00013ffc0001fffff7be00000000000efffff7fdfc4ffffff7fdc0600000041000000003fffc000800d00fffffffffffffffffe00000001015fffffff900000000000
B2[107] <= 640'hffffffffc7ffe600000003ffffe00003ffc4000fffffff000000000040efffff7ec0c07fffff7fcc0000000040000000003ffff0088c48134ffffffffffffffffc00000000c3cfffffff960000000000
B2[108] <= 640'hfffffefee7ff6e00000003ffffe00000ffe40007fffffef80000000067fffffde080001f7ff331c00000000040000000001ffff8000c40f94fffffffffffffff7000000000ffcfffffff960000000000
B2[109] <= 640'hfffffece7fff0c00000007fffffc080cfffc0007fffffefc840000006ffffffcc000000f7df100800000000000000000000ffff8800009fffdfffffffffffffb6000000000c7ffffffff820000000000
B2[110] <= 640'hffffffff1eff8080000003ffffec000efff80007fffffffcce000000edffffff0000000e410101000000000000000000000fffff00000d0f7cfffffffffffffe0000000400ffffffffffb00000000000
B2[111] <= 640'hfffffffc03ff80000000018f7600810fdf800027fefffffcff000000c9ffffcd000000000104010000010000400000800007ffff000108c07cff7ff7fffffdbe8000000401fffffffffef20000000000
B2[112] <= 640'hffffff7099ffc000100000121000000ebf980003f9fffffe9d000422e17fff7c000000000000000000048001200000003003ffff61018c79df7f3ffbfffefffe80000001001fffffffff000000000000
B2[113] <= 640'hfffffffc11ffc0000800000000000004df9800017dfffffffc000000c3ffff60000000000000000002400000000000001007ffff01000b09dfffffffff36fefc8000000103ffffffffffc40000000000
B2[114] <= 640'hffffffce33ff00000400000000000000f33c00017cfffffffe00018087ffff60000000000000000003400000000079001007ffffe000015dffffffbfff337c380000001ff3ffffffffffc40000000000
B2[115] <= 640'hffffffcc63ff000006000000000034003f7e00007cfffffff600038003ffffe80000000000100000034000000000fd003007ffffe0c0e0fcffffffffe01303700000001ffbffffffffff000000000000
B2[116] <= 640'h1ffffff887ff80000400000000003c00237600006f3ffffff680cf9131fffffc00000000001c000000c000000000e880f003ffff86800efcfffffffff08003f00000003ffffffffffff7000000000000
B2[117] <= 640'h7effff300eff8000000000000000e30003fe00006f3fffff7700dfb1303fff4c0000000004fd000000cc000000017f80f001ffff8c000eddfffffffec00018600100003fffffffffffffe00000000000
B2[118] <= 640'hfcffff0006ff8000000000000011fb80003e00000cbfffffff00ff98000fff78000000000ffc00181ffd00000003ff818001fffff800e47dffffffefc00010000000012fffffffffffff700000000000
B2[119] <= 640'hcf9fd80007ff0000000000000061fef90038000009bbfffffb07338c808fff71000000003fff0f181fff800000047f80800038ffff004779effefffffc1001000000000fffffffffffff708000000000
B2[120] <= 640'hfcfefc00027f80000000000000707ee00000000000c0ffffffe38b80181fff88000000007f7f9c1e9bff20000007ffc0000272ffddcc67fffeffffffffc680000000003ffff9fff9ffb9f00000000000
B2[121] <= 640'h1cff3e0000ff8000000000000020e3f30000170020007fffeb389980810ffff8000000007ffffc1fffff000000077fc0000002fffdcc6ffffffffffffffe00800000033fffffff99ff19fc0000000000
B2[122] <= 640'h1e0f3c0000ff90100c010000000003f00000bfdf80007fffe33c8b800103fff8000000007fffffcfffff8000000fff80000003ffffcd7ffffffffffffffe03c0000003ffffffffbfff18fc0000000000
B2[123] <= 640'hc600c00001ffd0000c200000000000000001fbfffcfffeffc08b0b800003ff3800000000ffffffffffffc0000007ff000000037fff6dfefffffffff0fffff300000003fffffefeffdffdfc0000000000
B2[124] <= 640'h8000030001ffc980771c0000001c000f0020bffffffffce0000000000001ff0000000003ffffffffffffc00210062f000000167ffffdfffffffffff0fffffb18000003fffffefffccf70100000000000
B2[125] <= 640'hffff8073c008000000800000107ffffffee3c0000000000001ffc000000007ffffffffffffc004003e3c00000010fcfffc3fffffffffe17efffff0000003fffffeffc6ff60300000000000
B2[126] <= 640'hfffc307fc31c0000000100b001767ffffff3000000000000017ff900000006ffe79fffffffc004001ffc40000000e037fdffffffffffc0227ffffc00008fffffffff06f960300000000000
B2[127] <= 640'h10001fffe7f3ef30001068ff8fe3881773fffc77e880000000000007ffbe000004ffee01fffffffc006001c81600000008023ffffffffffffc063fffffc00023ffffffffc467866700000000000
B2[128] <= 640'h11ffd5effdfff60037ff7fbdce0f9ffff99cc800000000000003ffff000003ffc003fffffffe080026f230000000000007ffefffffffff000fffffe800f3ffffffffef81ffb790000000000
B2[129] <= 640'h3ffdffffff7e0003fff7fffd61f1fffff9cf000000000000003ffff000021ff8000fffffffc0040226001000000000007ffffffffffffc07fffffe800ffffffffffff0fef3fc0000000000
B2[130] <= 640'h167fdfbfff83f8021fffe9f79f1fe7fffffef0000000000000007ff6000001ff8000fffffffc000020e003000000000003bbfffffffff1c8fffffff80ffffffffffffc7fcffde0000000000
B2[131] <= 640'h16ffff9fff8338470fffc103339ffff7ffffe8000000000000007f7600000fffc0007ffffffc400022f80b200000000001b0fffffffff9ebf7fffff00ffffffffffffffff7efe0000000000
B2[132] <= 640'h1000000007fff9cefce03c07fff980000097efffffffe000000000000001ff3e08016fffc0007f3ffffc400022f01f7000000000000007fffffffcf7effffffc77fffffffffffffff7efb0000000000
B2[133] <= 640'h71c00000007fff9cc0cf00e0dfff90000081fec7fffb1c040000000000063ff30080b7fffe001ff3ffff7c000000117e000001000000003fffffffff7ffffffffffffffffffffffeffeff30000000000
B2[134] <= 640'h7b000000009ffd6400cf9e20fefff0000000f9007fff00ec000000000004ff30001db7f3ff003fe0fd01000000003ffe00001d000080000037fffffffffffffffffffffffffffeffffdffd0000000000
B2[135] <= 640'h37fc000008fff66007fcf00fffff000000081001c7dffc6000000000080ff10079f3f7fff00ffe0380e0000000067f20001fe000389600003ffffffffffffffffffffffffffffff7ebfce0000000000
B2[136] <= 640'h878680000026fc20111983387ffff80000008000003ffee8000000000073fc001f73c3e37fffffc04400000000083ef90001fe0009afe00001ffffffffffffffffffffffffffffffe7fff08000000000
B2[137] <= 640'h9ef8f00c0007ffc0011807c17fff180000000000003ffffdc00000201c7fffc012f207387ffffec0040000000000fef00007fe0001fffee0007ffffffffffffffffffffffffffffffffffd0000000000
B2[138] <= 640'h1eff704d8006c18080000c83d9fffc00000000000007ffffcc0000fc0ffffe0003e00c183f9fff80000000000001fee0000fff6003fffff00000f3ffffffffffffffffffffffffffffffff0000000000
B2[139] <= 640'h6bf74c1000000000000800099ffec00000000000017ffffce80e6e7c7fffe0003c000003f9fff00000000000001ff00000fffe002fffff0000033fffffffffffffffffffffffffffffff80000000000
B2[140] <= 640'h83fde461000280000000800099ff0600000000000016e7ffff00eeefcffff60003e000003ffffe00000000000000ff000003ff8000fff900000007fffffffffffffffffffffffffffffff80000000000
B2[141] <= 640'h33ffce3f00000000000000001bffec00000000000003ffffffcfff7ffefff30012e000001ffff00000000000000318000013ff8011fff800000003fffffffffffffffffffffffffffffffc8000000000
B2[142] <= 640'hb37fff7f0000000000000100037ff8000000000000069ffffffffffffffff300330000001fff900000000000000700000017ff8001fff000000001ffffffffffffffffffffffffffffffff0000000000
B2[143] <= 640'h8277fbeb0001000000000000003f19000018000000069fbfffffbff7fffffe801310000003f9f000000000000000f100000ffee019ffe000000018fffffdffffffffffffffffffffffffff0000000000
B2[144] <= 640'h19efffff8800080000000000000020000003080010426837fffffffffffff008300000001fc000000000002400074000025384002ff8000000000ffffffffffffffffffffffffffffffffc000000000
B2[145] <= 640'h11feffffc00000000000000000000800000f000008000007fffffffffffffc0100000000000000100000000000000000000804003fc000020000ffffffffffffffffffffffffffffffffff000000000
B2[146] <= 640'h7eff766000000000000000001008000218080000000002fffffffffffffc0000000000000000000000000180000000000800003fc000000000ffffffffffffffffffffffffffffffffffc00000000
B2[147] <= 640'hefff26000000000000000001000000e386600000000067ffffffffffff8000008000000000c0013c9180b80000000000000001cf000040017ffffffffefffffffffffffffffffffffffe00000000
B2[148] <= 640'hccf820000000000000000000080003f3b22200000001f7fffffffffffd0000009f000000000ffe11f982110000000000000000c40000cc83e0fffffffffffffffffffffffffffffffffe00000000
B2[149] <= 640'hf3c00000000000000000000000003ff322000000001ffffffffffffed000000dfc30000000ffffff9b70100000000000800007c0003ffe3f0fffffffffffffffffffffffffffffffff200000000
B2[150] <= 640'hd0891000000000000000000010003ff33e0000000013ffffffeffffcd000105e4c00000005ffffffffff08c810020000d88003e0001fffff9ffffffffffffffffffffffffff190ffffe00000000
B2[151] <= 640'h8099000000000000000000010007fff38300008011e3ffffff7fffc981000864180000004ffffffffefe8f1bf0c6000999000000003fffffffffffffffffffffffffffffcc39017ffec0000000
B2[152] <= 640'hc000080010010000000000000007ffbee48c080084deffffffffffc10000836d800000010fffffffffe707e3ff00c83b8fc00000007fffffffffffffffffffffffffffff0001017fff80000000
B2[153] <= 640'h10000000000000000007fffff8bec0000ffefffffffffff80600007c800000007fffffffffe70ffedf0f40fdf03ec000003fffffffffffffffffffffffffffff000101ffff80000000
B2[154] <= 640'h100000000000010001800000000000007ffffff3f400007fcfffffffffffc0700007c000000007ffffffffffffffeffff69fe73668001c0019ffffffffffffffffffffffffffe000000fffe00000000
B2[155] <= 640'h88000000000000200000000000000000fffffff7f000003fffffffffffffc06010168000000007fffffffff7edefffffffdff73e23c00fc000ffffffffffffffffffffffffffe400000dffec0000000
B2[156] <= 640'h18c000000000000203000000000200000ffffffeff0000017bfffffffffffffec00040000000027fffffffff78840fffffff7ff1e7fc001e01005fffffffffffffffffffffffff400081ffffe0000000
B2[157] <= 640'h98100000000000383c00001000600000ffffffffe8000007bffffffffffff7fe00c40008000037ffffffffe810001ffffffffff7fe40003c1601fffffffffffffffffffffffff000081ffff80000000
B2[158] <= 640'h9b27000000000003fffc0001000000000ffffffffe800006737fffffffffff7fff3c4000c100037ffffffffe8000007ffffffffffdf3010700603ffffffffffffffffffffffffe8000017ffe20000000
B2[159] <= 640'h18f0800000000003fffc00188100000007ffffffff000002e17ffffeffffff7ffef34c187374077fffffffe400000007ffffffffdfff813e3d761ffffffffffffffffffffffffc8000017ffff3800000
B2[160] <= 640'hcf8402000000003fffe0000008100003fffffffffe000008ffdffffffffffffffe0f8b83fff1fffffffffc80000003fcffffffeefffc0ffcfc318fefffffffffffeefffffffd8000000fffff8800000
B2[161] <= 640'h87f8400001000003ffff80000000000037fffffffff00000007fffffff7ffffffffde739ffff1ffffffffff80000003f3ffffffffeffc0dffefc0197fffffffffffffefffffff80000003fffff800000
B2[162] <= 640'hc7b84c0001000003ffffc000000000001ffffffffff8000001fffffffffffffffffffff9ffff7ffffffffff00000003f7fffffff7fffc1fff8f80107fffffffffffffef7fffff80000009fff7fc00000
B2[163] <= 640'h6e1b6c0010000001ffffe100600000009ffffffffff8000003fdfffffffffffffffffffffffffffffffffff0000001fff3fffff97fff013ef3e000037bfffffffffffffffffffc8000008fffffc00000
B2[164] <= 640'h7e83fd0000000000ffffe000600000009ffffffffff80000006d7ffffeffffffffffffdffffffffffffffffc000001effffffffbfffe487fefc00803f9ffffffffffff3efffffc0000008ffffcc00000
B2[165] <= 640'h6781cd80810000007fff9800000000001ffffffffff800000049ffff3f7fffffffffffdffffffffffffffffe4c30010fffffffffffe00c831e000011ffffffffffff3dfffffff40000001ffffcc00000
B2[166] <= 640'he391fd80010000277fff8e00800000003effffcffff000800000ffff7f7dffffffffffffffffffffffffffff6ff801bfffffffff7d00000338000010ffffffffffff3fcffff9e41000003bffffc00000
B2[167] <= 640'h62bffd1c18800007ffff84009800000036ffffdecf1800800001ffffe6f9fffffffffffbffffffffff7fffffeffe19ffffffffffe100000021c000101dffffffffffffffffff06000000c3ffffc00000
B2[168] <= 640'h9c6fffc000643007ffffff60c00000001fffffce008000000001ffffccffffffffffefffffffffffffffffffffffffffffffffee60000000208000019ffffffffffffffbfffff600000001ffffc00000
B2[169] <= 640'h83fdffc000fe080efffffc23060000001cffffe40000000000007fffffc0ffffff7ffdffff7fffffffffffffffffffffffffffee00000000000000001ffffffffffffffffffff600000007fffffc6000
B2[170] <= 640'ha3cdffcc1ef88edefffffc22020000000cfcfe00801000000006ffffefe07ffffffffdfffffffffffffffffffffffffffffffffc00000000000000000b7fffffffffffffffffff00000007fffffc7000
B2[171] <= 640'h770fffee1ef98efffffffff0e00000040e807e00800000000007ffffeffcfffffffffdfffffffffffcffffffffffffffffffffc00000000000000000005fffffffffffffffffff00000000fffff3f800
B2[172] <= 640'h764ffff203fffffffffffffe34000000078126c0800000000003fffffdfcffffffffd9fffeffffffefffffffffffffffffffffc00000000000000000005effffffffffffffffff00000000fffffffc00
B2[173] <= 640'hf2fdff6303ffff7ffffffffe3c00000003182600800000000007fffffdfc3ffffffff93fffffffffffffffffffffffffffffff800000000000000000000cfffffffffffffffffd800000007ffffcfc00
B2[174] <= 640'h8279ff7003ffff7ffffffffe700000000198600000000000001fffff7dec1ffffffffc1fbffffffffdfffffffffffef7ffffff8000000000000040000004ffffffffffffffffffc00000037ffffefc00
B2[175] <= 640'h9a61ff7e33fffffffffffffc638004000188600000000800001fffff7feffffef9efe77fffffffff7ffffffffffffe7f7ffff99000000000001000000004fffffffffffffffffff0002007ffffffc000
B2[176] <= 640'hf973ff7f36ffffffffffffff731c000004679c0000000008001fffff7fff7ffffffff9ffffffffff7fffffffffffff3effffffc000000000000000000001ffffffffffffffff87ff000007fffffffc80
B2[177] <= 640'hbf79fc7f67ffffffffffffff73cc000000f08f3000000000000fffffffedffffffffff1ffffffffffeffffffffffffffffffff0000000000000000000001fffffffffffffffffffe0012cfffffff7c00
B2[178] <= 640'h1d383ceee7ffffffffffffffe7c400000039df3000000000000fffffffebffffffefffffffffffffe7ffffffffffffffffffffe000000000000000000000fffffffffffffffffffc0002cfffffff7800
B2[179] <= 640'h988001ce27ffffffffffffffffc7900000197ff600000000003fffffffedfffffffeffffffffffffc7fffffffffffffffffffff800000000000000000000fffffffffffffffffffc0012ffffffffe340
B2[180] <= 640'h8180808f67fffffffffffffffefef1e000907ffe06000001003fffffffecfffffffeffffffffffff0ffffffffffffffffffffffcc00000000000000000003ffffffffffffffffff800bffffffffffc00
B2[181] <= 640'h8100789fe3fffffffffffffffefe1bf00001fffe06800000007ffffffffcfffefbdffffffffffffe9cfffffffffffffffffffffde04000000000000000003f3ffffffffbffffffc00016fffffffffc00
B2[182] <= 640'hc1001099e7fffffffffffffffffe9b700007fffe00900000003ffffffffdfffeffdffefffffffede9cffffffffffffffffffffff6c4000000000000000003ffff9fe7600ffffffe00102fffffffffe00
B2[183] <= 640'hf83003b93cfffffffffffffffffefbf00124bffe01160000003fffffff7bffffdffffefffff8fede9fffffffffffefffffffffff7d6000000080000000003fff81016000cf9ffffc01bfffffffffff10
B2[184] <= 640'he0010086c6fffffffff7fffffff9f7fc0000bff804f8000002f9ffffffcf7f3fef7fffffffcf79f063bf9ffffffffffffffffffffe1c00800000000001003f8300000001303cffc09876ffffffffff00
B2[185] <= 640'h1c06ffffffffffffffffffeff80000fffc05f8e398007b7ffffdc07ff8feffffffffffefc360bfffffffffffffffffffffff1f01180030000000037f92000000000111ffc099e7ffffffffe700
B2[186] <= 640'h1c00ffffffffffffffffffffec0000bffc0fffe380004ffffff9e0fffefecfffbfffffcf0760bf7fffffffffffffffffffff87811e7c7000000003ffb00000000000003ffc1fdfffffffffe780
B2[187] <= 640'h8100ffffffffffffffffffffce00003ff80ffffff9006ffffff9014fffffdffe9fffffed0362be7ffffffffffffffffffffffeffe6fe00000000ffff9000000000000007f89bfdfffffffff6c0
B2[188] <= 640'h8100fffffffffffffffffffffe00003f784fffffff906ffffff800cf7cfffefeffffffe000c7b7f7ffffffffffffffffffffff3fe6ffff000001ffff80000000000000033bfbfdfffffffffcc0
B2[189] <= 640'h3ffffffffffffffffffffe0000b2f84ffffff8907fffffe000e779fffffffbeffee000c7bfffffffffffffffffffffffff7ffff8ff0000033fff800000000000000003b9dffffffffffcc0
B2[190] <= 640'h3ffffffff3feffffffffff00003080df7fffff907fffffe0c0e607ffffffffe7fec1000ebfbfffffffffffffffffffffffffff3cff060001ffff80000000000000003339e7fffffffffe00
B2[191] <= 640'h3ffffffff37fffffffffff60001000fffffff3915dfffb200002c0fef7ffce7fffcd001ebfffffffffffffffffffffffffffd93eff060718ffffb00000000020000071397effffffffff00
B2[192] <= 640'h7fffffffedfffffffffff81000001ffffffff7c3f7ffca0801cc107fc38200fffb320ff77ffffffffffff7ffff7ffff9ffffff97fe3fed3ffffc800000000000000882e0fcfffffff7e00
B2[193] <= 640'hffffffffffffeffffffff81c00001ffffffffe7fffff9830031f06ffff83887ffe3e0fff7fffffffffffffffffffff3ffffffffffffffffffffc80000000000000000c01ffeffffffcc00
B2[194] <= 640'h3ffffffffff7fdfffffff63c00003ffff7fffe7ffff71377173fceffffe1c83fff2c6bdf7ffffffffffffffffffffe1fefffffffffffffffffffdcc00000000000000001fffffffffc480
B2[195] <= 640'h1ff7fffffff3f3fffffff76007003fffffffffffffff83e7973fecefee60007fffecf9fffffffffffffffffffdffef067fffffffffffffffffffffc00000000000000009f7ffffffe7c80
B2[196] <= 640'h1fffc3fffffff7effffff7680c3e3fffffefffffffffc329f7ffffffee6801ffffe7f9fffffffffffffffffffdfffe0277fffffffffffffffffffff008000000000200007fffffffe3b00
B2[197] <= 640'h27ec1ffffffffffffffffec1c77fffffffffffffff9fb38ffffffffee6c003fff7f9fffffffffdbffffffffffffffe3e3fffffffffffffffffffffc1f200000000000007ffffffff0300
B2[198] <= 640'h1780000400fffff9ffffffffffcffff7fffffffffffffffffb7f7fffffffef90003fff3f9fffffffffffffffffffffffffc98037ffffffffffffffffffffff600000000000007ffffffff8000
B2[199] <= 640'h2016000fc0020000ffff3feffffffffdf1ffffffffffffffffffeff3ef3ff7fffef9100137fffdffffffffffffffffffffffffffc81c403ffffffffffffffffffffffc000000000001ffffffffe8c00
B2[200] <= 640'h183fc1fde00000007fffffffffffffff67f7ffffffffffffffffffcfb7cffffffff7e0c23dfffffffffff7bfffffffffffffffff0006081ffffffffffffffffffffffde20000000001ffffffbf90000
B2[201] <= 640'hfffe9fff80000003fffffffffffffffefffffffffffffffffffffeffffffffffffe30477fffffffffffffbfffffffffffffffff8004000fffcffff7fffffffffffffff00004000000fffffffff0003
B2[202] <= 640'h3effffffffc0000003fffffffffffffffc7ffffffffffffffffffffffffffffffffee300ffffffffffffdbf37ffffffffffffffffc0000000fdfffff7ffffffffffffffff8004800003fffffffff0000
B2[203] <= 640'hffffffffffe0000001fffffffffffffff33ffffffffffffffffffffffffffffffffe6080fffffffffffe81017fffffffffffffffff8001183b1f9fbffffffffffffffffffe0f7d00007efffffeff0030
B2[204] <= 640'hfffffffffff032f800fffffffffffffff13fffffffffffffffffffffff7fffffffff7680fefbfffffffed8007dffffffffffffffffe0001f38fff1bffffffe7ffffffffffff8fdf0007fffff3ff30000
B2[205] <= 640'hfffffffffffc3ffc00bffffffffffffffc3ffffffffffffffffffffffffffffffeffe300fce1fffffffc98187c3ffffffffffffffff9480bfc3b7fffffffff7fffffffffffffff9330efffff3ff20080
B2[206] <= 640'hfffffffffffffffe00fffffffffffffffc3ffffffffffff77fffffffffffffffff9c0000fcc07fffff798080003ffffffffffffffff9c481fe1f3fffffe7ff7bfffffffffefffffb7bffffff9ff60080
B2[207] <= 640'hfffcfffffffffffe007ffffffffffffffc3fffffffffffff7ff7ffffffffffffff1c00001c0466fefee181000077fffffffffffffcb9e6c9dffbfbfffefffff9fffffffffffffff9ffffffff9ce60000
B2[208] <= 640'hfff97ffffffffffe00ffffffffffffffff7fefd8ffffff7ffff8db7ffffffffffc00000042903df0ff000400007fffffffffffffff7800667cfc39ff7eff0f3f7ffffffffffffbeffcffffff163f8000
B2[209] <= 640'hfff9ffffffffffff000ffffffffffffff83f7fff7fffffffffdffdfffffffffcff800000400013f97c000000001fffffffffffffff000072741ff8ffff7f3eefffffffffffffffcfffffffff84031000
B2[210] <= 640'hfffffffffe3fffff801fffffffffe33ffe7ffd9ffffffffffffffdfffff3fffeff810000380003387800000000037ffffbffffffff8f0039c2f9f8e7ff7ffcff3fffffffffffffffffffffff80033800
B2[211] <= 640'hfffff3ffdc7fffffc003ffffffff00001cfff9ffffffffcffffffffffff7ff7ffc000001980000383800000000003fff810007fffeffa019c6ffffffffffff7e3ffffffffffffffffffffff910038000
B2[212] <= 640'hfffff3fc01ffffffc001ffffffff000038fffffffffffff0ffffffffffffffe67c0000079800203800000000000010fe000001fffffef08f8c1ffffffffffffff8fffffffffffffffffffff9510e8000
B2[213] <= 640'hfffeffcc0107dbffc0017ffffffe000038fffffffffffe307fffffffffb7ffe40700000398000030800000000000033c0000003ffffef086be3fffffffffffffffffffffffffffffff7ffffc700e0000
B2[214] <= 640'hfffffe8000049ffff0000b7fe018000000fffffffffffc0307fffffffff7fe0f030000017e000100800000000c00000800000001fffff386bbfffffffffffffffffffffffffffffffffffffcb88c1000
B2[215] <= 640'hffffde80001000fff800003cc0000000001feffffffff80007fffffffffffe98000000017e000800000000003b000000000000003ffffffffbffffffffffffffffffffffffffffffffffffecf884e000
B2[216] <= 640'hffffff000000009ffc00000460000000007fffffffffec8000ffffffffffff86000000000f000000000000077c600000000000000fffffffffffffffffffffffffffffffffffffffffffffb3ab0700a0
B2[217] <= 640'hfffffe000000000fff80000000000000003fffffffff400000fffffffffffe07000000000f0000000000003ffffc0000001f000007ffffffffffffffffffffffffffffffffffffffffffffd36e148000
B2[218] <= 640'hfbfffc000000001fffc0000000000100003fffffffff0000007fffffffff7e0000000000070000000000007fffff000000fffc0000efffffffffffffffffffffffffffffffffffffffffff77df168450
B2[219] <= 640'hf7ffc0000000001fffe400000000300000fffffffffc8000003fffffffffff800000000003c00000000000ffffffe00001ffffe0004fffffffffffffffffffffffffffffffffffffffffffa0d8178448
B2[220] <= 640'hfffffc0000000003fffe800000003000007ffffffffc8000011e0ffffffeff8000000000c3e00000000001fffffff001fffffffc000dffffffffffffffffffffffffffffffffffffffffffa01c10c010
B2[221] <= 640'h7e7c3c0000000020ffff90000000ff00001fffefffb80000008c03b9dffffc0000000000e1c00000000003ffffffffffffffffff00017ffffffffffffffffffffffffffffffffffbffffffe08394f814
B2[222] <= 640'h4e1800000000002003fff8000006ffc0003fffefff800000000100110eff38000000000020000000001800ffffffffffffffffff00017ffffffffffffffffffffffffffffffffffbffffff71a7d73084
B2[223] <= 640'hc68000000000000001ffff800000cfc000ffff7cff80000000010000dc7e80000000000020180000003c003fffffffffffffffffc001ffffffffffffffffffffffffffffffffffffffffffff9282105e
B2[224] <= 640'h8900000000000000007fffff80000e0001fffff018000000000000005c6f98000001000000c00000003e003fffffffffffffffffc0007fffffffffffffffffffffffffffffffffb93dffffd0d828bb85
B2[225] <= 640'h9800000000000000007fffffff000e0000ffffc00000000000000000083e98000000000007300000007f803fffffffffffffffffc0003fffffffffffffffffffffffffffffffffa978ffffd8e2769382
B2[226] <= 640'h7ffffff168e0000ffff000000000000000000003c6000000000006018008001ff803fffffffffffffffffe0000ffffffffffffffffffffffffffffffffec325fffeca454710a3
B2[227] <= 640'h6000000000000000000ffffff3fde0001fffc0000000000000000000000600000000000e00001f003ffc03ffffffffffffffffff00007fffffffffffffffffffffffffffffffed5e71fffdcb0a3ee86
B2[228] <= 640'h2000000000000000000ffffffb8ff0001fff000000018000000000000000000000000000000017801ffcc7ffffffffffffffffff00007fffffffffffffffffffffffffffffffe98e45fff50901eac97
B2[229] <= 640'h7fffffe3eb0001ffe000000000000000000000000000000000000000003800fffe7ffffffffffffffffff00007ffffffffffffffffffffffbffffffffe03884ffe41e1385aa7
B2[230] <= 640'h1fffffe3e200007f00000001c2000000000000000000000000000000000000fffe3fffffffffffffffffe00007fffffffffffffffffffffffffffffffe416a4ffa6c710de267
B2[231] <= 640'h1fffffe7c000007e0000000038000000000000000000000000000000008303ffffffffffffffffffffffe00007ffffffffffffffffffffffc7ffffffff7cc78ffa668b01a6e3
B2[232] <= 640'h1fffffffcc00007c00000004e00000000000000000000000000000000000003fff001fffffffffffffffc00003ffffffffffffffffffffffffffffdffe713afdf4523062672c
B2[233] <= 640'hffffffffe00003800000003e0000000000000000000000000000000001f033ffe0019ffffffffffffffc00003ffffffffffffffffffffffffffff7fefd496e7e460e81b9371
B2[234] <= 640'h5ffffffefe0000000000003c000000000000000000000000000000000870307fe00017fffffffffffffe00003fffffffffffffffffffffffd7fff7ecf32a21da044200b7c47
B2[235] <= 640'h1fffffffff0000000000001e000000000000000000000000000000000000307fff0017fffffffffffffe00003ffffffffffffffffffffff3c7fffffc89590cfe6311b7af492
B2[236] <= 640'h7ffffffffe08000000000000000000000000000000000000000000000000000ffe0003effffffffffffc00003ffffffffffffffffffffff38fff5ff8c38d67f779808274df3
B2[237] <= 640'h1007fffffffff080000000000000000000000000000000000000000000001e0000fff00406ffffffffffffc0000ffffffffffffffffffffffeefffff7edca2a4ddb7a23cc03abc
B2[238] <= 640'h2007fffffffffc00000000000000000000000000000000000000000000000c00003ce00006ffffffffffffc0000fffffffffffffffffffffffeffffffe78965f269797d20170b3
B2[239] <= 640'h1effffffffffc0000000000000000001000000000000000000000000000000081000002027ffffffffffe80000ffffffffffffffffffffffffffffffc7804609bc3a134443383
B2[240] <= 640'h7fffffffffffe00000000000000000000088000000000000000000000000000008fc000000ffffffffffe00000fffffffffffffffffffdfffa7ac2ee565d806df81d3040eeae1
B2[241] <= 640'heffffffffffffe0000000000000000000078d800000000000000000000000000018400000003fffffffffe00000fffffffffffffffffffffffffafbb849aab067fa31cb03c7edb
B2[242] <= 640'h3fffffffffffffff00000000000000000000f0f800000080000000000000000000010000000003fffffffffe000003fffffffffffffffffffbffffbfbbef0fc0d283f761f8072d7e
B2[243] <= 640'hc13fffffffffffffff80000000000000000000e7fc003e71fc000000000000000000000000000000fffffffffe000003fff7fffffffffffffff9ffddbebff4c90dac68f02768381095
B2[244] <= 640'hc01fffffffffffffff8000000000000000000087fe01fffbff800000000000000000000000030000fffffffffe000000ffeffffffffffffffffdffdd9fee67fb76287ef5c3886ad8d4
B2[245] <= 640'h3c07ffffffffffffffc000000000000000003c0fff07ffffffc000000e00000000000000e007e0003fffffffdc00000000effffffffffffffffdbbfcdfee7784d26c897d0058ef7d4f
B2[246] <= 640'h3edfffffffffffffffe000000000000000863c87ff0ffff7ffe00000bfb8000000000001710fe00003fffffc0000000000fffffffffffffffffbbbfd5ffe761c20246a5e9284eb2f48
B2[247] <= 640'h7fffffffffffffffb000000000000013fff7effff1ffffffff80001fff80000000000017bbee00003fffffc0000000000fcfffffffffffffffbb3f74f7e45b6648174e4c1e046981a
B2[248] <= 640'he0033001003c07ffffffffffffffff00000000000007fffffe7ffffffffffff0000ffff80000000000001ff8000000fffffc800000000ffffffffffffffffff3fb1c4f3f75418416a2cdc384017626
B2[249] <= 640'hce3007800000fc0fffffffffffffffe00000000000000ffffffefffffffffffff8001ffff80000000000003fa8000000ffffff040000000ffffffffffffffffffad960cebf252f1401eb5c41f832c05d
B2[250] <= 640'hff3f7fe100007cffffffffffffffffe0000000000004ffffffffffffffffffffff003ffffc0000000000001fe8000000ffffff0800000003fffffff00407d59f9e62de331f7c66a0bb840d4b8c20480e
B2[251] <= 640'hfffffff0000000ffffffffffffffff8000000000001fffffffffffffffffffffffe0ffffff1800000000001fe8000000fffffff800000000fffff0000000000765b08aa19fda50938007cee01c1630c1
B2[252] <= 640'hffffffff8000037fffffffffffffff800000000000ffffffffffffffffffffffffffffffff7f0000000000ffc0000000fffffffc00000000ffffc00000000003dc8e1cb2bf1e890c1082dee96b218849
B2[253] <= 640'hffffff7fec00003fffffffffffffff800000000023fffffffffffffffffffffffffffffffffff800000000ff00000001ffffffff0000000000ff000000000001168e209b7ea9269485aeeb0e403d1928
B2[254] <= 640'hfffffffffff000ffffffffffffffff800000000077ffffffffffffffffffffffffffffffffffc0000000007f00000003ffffffff8000000000fe0000000000016771306dfb8df03914d0e2a248daedc3
B2[255] <= 640'hffffffffffffffffffffffffffffff800000000021ffffffffffffffffffffffffffffffffffc0000020000000000007ffffffffe0000000000000000000000d1e760c1c7f8cf49e39047bb121882085
B2[256] <= 640'hffffffffffffffffffffffffffffffa00000000000fffffffffffffffffffffffffffffffffffc00000000000000000fffffffffe380000000000000000000166aba24397d1290990242edfc871b104a
B2[257] <= 640'hfffffffffffffffffffffffffffffff000000000001ffffffffffffffffffffffffffffffffffffc000000008000400ffffffff8e000000000000000000000452af534b869120514008cd4eea602c893
B2[258] <= 640'hffffffffffffffffffffffffffffffffc000007f000fffffffffffffffffffffffffffffffffffffffa80000c000e00fffffffe000000400000000000000608b7010e28b59cc718213bcdab9a16ba9f8
B2[259] <= 640'hfffffffffffffffffffffffffffffffffc001cff8007ffffffffffffffffffffffffffffffffffffffff0000fe03f81fffffffc000000ef000000000000000023f2d830518e62c265c82c179e44ee068
B2[260] <= 640'hfffffffffffffffff03fffffffffffffffc0fffffc03fffffffffffffffffffff3ffffffffffffffffff0c0ffffffeffffffff8000013fff0000000000000008130c0eb3fe31100e4064027ce338a7c0
B2[261] <= 640'hfffffffffffefffff81cffffffffffffffffffffff23ffffffffffffffffffffe7ffffffffffffffffffc7ffffffffffffffff8000007fff0000000000000024d90cabdf064b80e14d0364f3a3421209
B2[262] <= 640'hffffffffdffc031fffffffffffffffffffffffffffe3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000010c000000000000009a5a288927a08aa719fca06d54631ac725
B2[263] <= 640'hffffffff9ff00000ffffffffffff011fffffffffffe03fffffffffffffffffffff7fffffffe7fffffffffffffffffffffffffffc0000000000000000000001c56a99da30e44502e49398ef97324e02a1
B2[264] <= 640'hfffffffffffe00007ffffffffff800017fffffffffff8ffffffffffffffffffffffffffffffcfffffd7fffffffffffffffffffffffc0000000007fc000000c0f482f1b902d9e07a668ab0cdf8904af2a
B2[265] <= 640'hffffffffffffc0007ffffffffff800001fffffffffffdffffffffffffffffffffffffffffff00700e00ffffffffffffffeffffffffffffff0000ffff800045a8032cc020fa1ed27349a201a410050de7
B2[266] <= 640'hffffffffffffff37ffffffffe0000000001fffffffffffff7fffffffffffffe3ffffffffff0000000001ffffffffffffbfffffffffffffffffffffffc00009b3dc304c08462749666080ec2f25b2004b
B2[267] <= 640'hffffffff80ffffffffffffffc00000000007fffffffffffe3fffffffffffffc07fffffffff0000000001ffffffffffff0fffffffffffffffffffffff3e839a9c6889d3086569ecd3060400aee4862672
B2[268] <= 640'h7ffffff001fffffffffffff8000000000007effffffffee3fffffffffffff801fffffffff007f800000fffffffffffe8ffeffffffffffffffffffffffff415613ef0b0ec9765d252ea632d51d108a18
B2[269] <= 640'h7fffff000ff1fffffffff800000000000000ffffffffc43fffffffffffff000ffffffffe00ff800000fffffffffffe3ffc1fffffffffffffffffffffff01969edb55138223922dfa4ad85ac8a1c581
B2[270] <= 640'h1fffff030e003fffffff300000000000000000ffffff003fffffffffffff0003fffffffc00ffe000008003ffffffff7fe0001fffffffffffffffffffff9413dbb117c138d922cacb4141abb0a44ec0
B2[271] <= 640'h7ffffff8e007bffffff0000000000000000007ffef9003ffffffffffffd0003fffffffc00f8f000000000ffffffffff800003fffffffffffffffffffff85ef671a4f16e0f331cf14f9345388ed100
B2[272] <= 640'hffffffff8000cfffc00000000000000000000fffff0001fffffffffffffc01ffffffffff8f8000000000003fc3ffdf0000000ffffffffffffffffffff90315cdb86d5d779e9c40048a901a49a2510
B2[273] <= 640'hfffffff3800003c00000000000000000000007ffff0003fffffffffffffe03ffffffffff8f8000000000001ff9ff00000000000ffffffffffffffffff85e363f74ed3043997a420828e7970012e72
B2[274] <= 640'h7fffffe0000001800000000000000000000001ffff806ffffffffffffffe078fffffffff8ff8000000000000f83f00000000000ffffffffffffffffff58811d8333086be1b38d25a85c037f89a148
B2[275] <= 640'h7fffff83800000000000000000000000000000fff3f07fffffffffffcfffff8fffffffff8fc0000000000000011f00000000000ffffffffffffffffff7c9b2d537613028e04df478b2471569918d2
B2[276] <= 640'h38fffffffff8000000000000000000000000000003ff1ffffffffffffffefffffffffffffffef80000000000000039e000000000000ffffffffffffffffff4680d9c31956f43ba1b845f4671a55391e4
B2[277] <= 640'hfffffffffff0000000000000000000000000000001fb1ffffffffffffffffffffffffffffffef00000000000000003c0000000000001ffffffffffffffff3c8a4c5be10204c2b412c411f216c8573c5c
B2[278] <= 640'hffffffcc0700000000000000000000000000000000713fffffffffffffffffffffffffffff7effe00000000000000100780000000000ffffffffffffffff006d8c3f62530187b08e4240499a68202438
B2[279] <= 640'hfffffe000000000000000000000000000000000000201fffffffffffffffffffffffffffff3fffe00000000000000000fc0000000000ffffffffffffffffdf2191750082127a03aaa47e8fa6a446601c
B2[280] <= 640'hfffffe000000000000000000000000000000000001c00fffffffffffffffffffffffffffffffffe0e000000000000001ff80000000e0ffffffffffffffff4a42f185a4ba745559a86100b98d17ad031b
B2[281] <= 640'hf007fc0000000000000000000000000000000000010007ffffffffffffffffffffffffffffffffe0c000000000005807ff8000000000ffffffffffffffff3504b2c478a81174f165e275f2e07a03008b
B2[282] <= 640'hfc0000000000000000000000000000000000000007ffffffffffffffffffffffffffffffffffffe00000e001f81fffc000000000fffffffffffffffdf26236c3b849da23b0037041ba2c1e83391d
B2[283] <= 640'h3c8000000000000000000000000000000000000000fffffffffffffffffffffffffffffffffffce1c000f01ffefffff800000000ffffffffffffffdc148ec4e6fd84aedd651870e0e379cb6b5582
B2[284] <= 640'h8000000000000000000000000000000000000000fffffffffffffffffffffffffffffffffff8e1ffe0f89ffffffffc7f00ffffffffffffffffffd96c42e8f338ffff5e839267af6402c3c6d739
B2[285] <= 640'hfffffffffffffffffffffffffffffffffff0e1fff1f99ffffffffcfffffffffffffffffffffffb327374a1e658d3a7633091ae044a0b209c04
B2[286] <= 640'hffffffffffffffffffffffffffffffffffffe0e1fff9fffffffffffffffffffdffffffffffffffedb1ad0f23a2848c692e92c5c4e0991c022805
B2[287] <= 640'hfffffffffffffffffffffffffffffffffffff5f5fffdfffffffffffffffffffffffffffffffffff88091e080c8818c31f8fa30ada3280b31a1ef
B2[288] <= 640'h737ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffad331f339c60024523963325e443865c49985
B2[289] <= 640'h717fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7d6502c87e43c80941072d052c5526f6110c35
B2[290] <= 640'h30007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbf9c691a348b4b984533f524d2b47d4f61828b
B2[291] <= 640'h78017bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8c9e6415194a49595746af023842f278780666
B2[292] <= 640'h7cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb82e946ec2387086268902c55fd8eca51192b4
B2[293] <= 640'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdccfae227846d29110274fb7017e2b6c0578c6da
B2[294] <= 640'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80ffff80080782f83d540311a08d6c1d9229a0a0f1070d628
B2[295] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8f1fffffe00000000000002ddf0e3809450acbc5f17b47b7925f81709293
B2[296] <= 640'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcc001ffff800200000000000215be951d2748a7b1a2f862f229bd42b09970
B2[297] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffee80000000000000000000000c0184fec8c5299de0ac9f2a3a2a03e20043b10
B2[298] <= 640'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffffeea0000000000000000000000001e3d275bc13822a2b1c6190d974fe9088f590
B2[299] <= 640'h13fffffffffffffffffffffffffffffffffffffffffffffffffffffff880000000000001c00000000001284d30968929216eafe678259c9bc8d28e277
B2[300] <= 640'h17fffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000041ec04000c010505e07a4a600cd277c1740c6527a6b38a9db22
B2[301] <= 640'h7ffffffffffffffffffffe7fff3fffffffffffffffffffffffe30faa0000000000001fdcc0085ff4551ecd98c67480048899fe8a11900b394e04a200
B2[302] <= 640'hffffffffffffffffffffff3ffbffffffffffffffffffffffff080000000000000000ffd0e40cffffffc7fbc2035872807e0c645e1101072b88852706
B2[303] <= 640'hfffffffffffffffffffff01f82cffffffffffffffffffffe7d3c0000000000000000ff46ee9eff7fffe035d2118a77291a5dfec2e3508c2ce788f57c
B2[304] <= 640'h500000000000000000000000000000007fffffffffffffffffff382fc7f9fffffffffffffffffff91e19e0000000000000077f37b76a827fff41945c5cdb0823fccd204162c441898b541d15
B2[305] <= 640'h780000000000000000000000000000007ffffffffffffffffffca02f43ddfffffffffffffffffc00fe11fc0100000000201cffef2fb80007fec4ec90ec8c620b77220fe0923f5acd39ec114b
B2[306] <= 640'h788000000000000000000000000000001fffffffffffffffffe509cfc3c1fffffffffffffffffff9fffff80000020000001c4f216be7003e01a590100c89134acafb07a462c0148f9ef46c40
B2[307] <= 640'hf8e000000000000000000000000000001fffffffffffffffffd40360feddffffffffffffffffffffff01f800030fc8b000001efdd078000eff8a71476a04aa4f6306e8760067ca0546c048b0
B2[308] <= 640'h7e0000ffffcc000000000000000000000000000fffffffffffffffe395e453bfe07fffffffffffffffff1ffffffc007ffff80ffeffe0261ebafffffc233060a500800652ac49d7b131f64264309021
B2[309] <= 640'h7e0001fffecc000000000000000000000000001fffffffffffffff986266fffff007fbfffffffffffffeffffffff1e80009efffe3f0970d0ce7ffff806ecb04f19483787418e39019c683f100c1c09
B2[310] <= 640'hfffff8fffff0cc0000000000000000007f000000ffffffffffffffff9cdfc5fbfefb079dfffffffffffffffc00000fe0ff00fac0600000e5b032fffe7d0bcb191d04e081f3e2059549d82534e0bc0480
B2[311] <= 640'hfffff8ffffc0cc000000000000000000ff000001ffffffffffffffff8040fefefff8186efffffffff8007cf0000000003ffffaa79c000074399b13303d232a8109e0a465341a08041035396c1355a881
B2[312] <= 640'hffffffffffe7fffffcffff0000000000ffffe003fffffffffffffffc0081ff9ffffdfe72ffe000f902fc763fffffffc000fe1dc900020132539f100045d685e2278030e20c92dac76199dca37598c830
B2[313] <= 640'hffffffffffffff1f000000ffff040303000000ffc0ffffffffffc3ff000cfc180001600c00830007ffff84bffff9fe000066f3df00804025e66370000751f92c308209e313dc76f14130139386cce250
B2[314] <= 640'hffffffffff7effffffffff00d0f0fe00feffffc0ff00003ffffff800fffe03800001e079066cfffffffff0f87a30f8000013c7b6000042011aba2800336bbc00d041910044349c43417af9f537c89003
B2[315] <= 640'hfffffffffffffefff00f00ffffff0000000000000cfff0000000003ffffe1f7fe7e0fff07859ff7f6083f8087c6cfb0000107dc0000b01ed2593100e92db821560c945700235259023588149698c8a0e
B2[316] <= 640'hffffffffffc180000000000000030ffff800000000000000000000080000007fffff1c9f7c7f3ef9607ffc0000c401e0001f8000000300f5b6f3800ee7ce6cb208fc24a04c6631eb4163904338426164
B2[317] <= 640'h3fffffffffffffffffff00000000003fffffe00000ffff0000000407ffcfff0fffffffc48f407ce600800001e0000800000001013541585003a6c83ebf08a16c454dda0891cb5427a75c8c08e1
B2[318] <= 640'h7f30000000000000fffffffffffffe000000000fffffffffff0c0000000f8ffefffeff37ee330c08e6c083080000300006103a00008f77609971e011d6b7c56e44196e8496538216022dfad2a404859
B2[319] <= 640'h7fffffcc0000000ffffffff7ffffffffffffffffffffffa0000000000dffffff6e07f4e0f886f9003df80000000006000000009e100a53094001a994e5712181058c360b1b0e222345197289d0c
B2[320] <= 640'h3fffffffffffffffffffffffffffffffffffffffffffffffff8c000180000cffffffee03cff20201dc0fff1670000000000002af06a0d62eee540001fe900fa9328ce085eb00db941c61b15062e460a
B2[321] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffff080001f1f03ffffffff078fff737f80e0fd003a00000000000011c84f3956887444006eeb813adceb6003997e21c6e0c05cd0126460ac
B2[322] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff000007ff07ffffffffff879c000080ffe040006000000000006576bc5a13dab43400601222222611c8612065331761396364c8204648
B2[323] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff000001f803ffffffffff8c080000183f00000009018f8000004e30d2e63a0f4976dbaa49000c43187c480e60721c4841a429e22852d4
B2[324] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffff31c00000e003ffffffffff308000fcf87f0000000600f10000003a0c46431d24a1da20816681821116342833d6117b40c3d2e1e77884a3
B2[325] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffe0080000000007fffffffff20800000007fff000e00fff80000000ddeb07a148a264221c828c988981f5e64425775268107d5af830a4081
B2[326] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffe0000000000003ffffffffff1e07900011dfffffe808077ffe0194df7ac8ce20557ac90595304662202824442385c50118ccc95e1123066
B2[327] <= 640'hf1ffffffffffffffffffffffffffffffffffffffffffffff0000000000001ffffffffffffffffe38000000f0ffffbffeff9fcca9d97c6c01fe7a65b852ec8242a9e750044008ff093e9d3c528620e0
B2[328] <= 640'h1800013fff0fffffffffffffffffffffffffffffffffffffffffffffff00003effffff3ffe000002f1800000fffc003fc7ff9d259db82e381acd0254b1b6684cc1d031144656607ac825420c191a5480
B2[329] <= 640'hc00000ff000000001f1f0007ef000000000000000000008000fffffffffff08000ffffffffffff800000007f5f7f8071ff8000964bac24060576e84c50ea5f1d72728c08043122b380081aa1e1384cc0
B2[330] <= 640'he3ff8007000000fffffd0000c1800000000000f4e03f000000000000000000fff8709fffff800000000fff7f000000fc3f800222a31c6e8904f87802dee80acfd33b2c10086f3a214012ae1a24da4289
B2[331] <= 640'h8fc000000080000000001ef80fffffffffffffffffffffe00000000f3ffffeffffffffffc378ffffffff0000000fe00087fe1871627e03003a995b510c4c38674e4a330c2001640400444f12a0c43c31
B2[332] <= 640'h1ffe600000000fff8008000fe000000000001ffffff7f3ffffc001fff0000000000000000fffcfffff800007033ffff03ff51579f7beb6260e7832d9a4a01e2a1d068101070261ec028378d3028066e
B2[333] <= 640'h87fffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000f807ffff7ffff0c0003c21ffffffffde2b510fc3ed5a3c408932421ffe041c031a1c71439b400016190a70321f
B2[334] <= 640'h3fffffff1f80ffffc0fff0c3ffffffffff003fffff3fffe0fc0000000000000003e007fffffffff8fe003f00f87effff41c1e485ae432a9681ccc37a1d796d46ef0c6c44d62001906a13da4a6c2f
B2[335] <= 640'h8003ffffffffffc0ff7880003c3effff8800f1f0ffff3ffbff800000000000000000000003f7e07fffc0ff7ffffcffffbfffae0a2e0b26052083dd39080a240b182e98040020a27d482de0b5b3a4163a
B2[336] <= 640'hec007cfc00ff0000600000000000ffffffffffffffffffffffc3000000000000000000000130e1ffff00000fffffffffffb733416019c5fa833f50845cccfbc821e6bc4e43027581404ce8333894182e
B2[337] <= 640'hec00000e000000000000000000001fffffffffffffffffffffc3000000000000000000000000007fff803fff1ffffffffc7e3d25289261669c520135766d21005012c20c2044484188338a18fe761b90
B2[338] <= 640'hfcf001e00000000000000000000001fffffffffffffffffcff800000000000000000000000000c3fffffffffffffff9ffffe812e31a984369458708927483022200241c336608db00475b7278544081a
B2[339] <= 640'hfe3e00300008000000000000000000fffffffffffffffff80000000000000000200000000000000f3dffffffffffffffffef65dac007a7f61825912740702c0075a3076239088d5b5818304391881004
B2[340] <= 640'h730001000002000000000000000000039fff801f1fffff800000000000000000ffff0f0000006000100fffffcffffffffff86010d02e0b271827904f923b9eb614919522080c348b18314c8317823028
B2[341] <= 640'h6fff03f800000000000000000000000003fe00030fffffe000000000000000007fff9f800000f000011800ff3bffffff1ffdd3a6de278c1b1548821107701f4244a00082b90e32ac0610886d86c66877
B2[342] <= 640'h49ff818c00000000000000000000000000000000020028000000000000000000fc3f00000000b000039fff3f93efffff60febdb4c33900af1834de58f31237224070360228601dc88208239240116c46
B2[343] <= 640'h32ff983000000000000000000000000000000000000000000000000000000000400600000000d000039fffe3ffe024f3f3c0241087d5245150a14d28e8816736100b9c8098120157002239901b10384f
B2[344] <= 640'h3f00180000000000000000000000000000000000000000000000000000000040a0050008401800231ffc001840c0a06e64dc4063c0053048ab0611a3771d80493b831808802024c207252810f31331
B2[345] <= 640'h700000000000000000000000000000000000000000000000000000000000060c200080080000103c5fd000007f8cb8003b67e81e904a0908c7fa8c82861e4c45b21c109800004943b2006f2880c20
B2[346] <= 640'h40f000000000000000000000000000000000000000000000000000000196c0000acfa0040194006600ffd8cfc01e3ffffc240d7c7c18066d50c6d944ca346401e0790c000e01040062208901b880052
B2[347] <= 640'h3f810000002000000000000000000000000000000000000000000000986f300dce0dee48f259c03c32b8800083fffffff83c110a7a33aa3cab30350a01b845d400a230c61028b01319082210263804
B2[348] <= 640'h7fe000000000000000000000000000000000000000000000000000ef779efff2c0b71680825c303aac001e01f13ffbfff8a69a33734576051b01047442921a00d28000844c38331100140621323d42
B2[349] <= 640'hffe000000000000000000000000000000000000000000000000003fb0ce1f10b9a5c7868ed00001b62000003fc31fdbff20726a2c05644006750615831883cbc4bac608c5c0d110818126040700049
B2[350] <= 640'hcfff0000000000000000000000000000000000000000000000000060e07f807d1806a8e830c9600a362003ff1ffc7e7fffb289a038a0063488048b9ea79cc11dd141a10415c48006404000071a40344
B2[351] <= 640'hdfff802000000000000000000000000000000000000000000000007ffe09c3040480c0006110be0136003ffffffe4000ffe830a90183110a210e00d70708dd629403ae48302012436021066ab060101
B2[352] <= 640'h7ffff83000000000000000000000000180000000000000000000003ff30191ac92c2aab7e452b83a269fdffffbff27f9cfc4b429104201250a1800c44486081c8609620469207207083004c8d740daf
B2[353] <= 640'hfffffe000000000000000000000000003000000000001c002801007ffff8080e511e8624f39ac5d2ac06bfffffff3fe9f850200533d78cb9a225838b19d9ee441a608980401188026418226052e1910
B2[354] <= 640'hbfffff8000000030080000000000fff80000300000003f000007fffffffc0c6418f7acdb19ae4443af7163f7f7fffc781841141415b622240819098c0081604e0624c544d06c5444482422245080018
B2[355] <= 640'hbfffffce8000003fc40001f8000f0c0f8000000ec3f03fff00f7fffffffc005a038b554bacdeeac7f183007fffeff0783dd0ebd711989c1419b8931053369b843254070230011800242890602302122
B2[356] <= 640'hffffffffff6000004000ff8000087ffe78000000fff07fe7fffffffffff6032a58dc82f4732d6d2341293ffff4900020344e838c6aa1d46b08090c709185ba2010e09980081100c4b40318083302924
B2[357] <= 640'h1bffffffffff702ff93804000001f0003c003f7e73ff0ffffffffffffffffeb3c65031dc8d8b081031176fffffc8c000036c2340d0436e2de074d84aca288438191831a102000450630120865900010c
B2[358] <= 640'h1bffffffffffff20ff0001900003000007003fe7bfff1fff3e3ffffffffeffb21c1925401c804240412837ff3fe8e0000360a30c60250883129240cf210126188301480700004400217020002e4a69a1
B2[359] <= 640'h1bffffffffffff79000006606080000000ff00ff0ff81fffffffffffff7ffff9711911506930e2a861d366fc00726000016394708b410069a3ba3f0972f35927201218c3000110188800270180042500
B2[360] <= 640'hffa1fbffffefff880000000000000a0001f0001c0011fffffffffffffff006ca62920c664b41a98318a87f8014691e0012236bc44474491a7e5738cc86b0ca71007800c00c2f01008f0130000004000
B2[361] <= 640'h13c5812f9effffe0f8000000001e000f80000000007ffdffffb9fffffe0700618d1763008080a71ee19f070003d0f4e8fc80ae6064999361a282a1333039601482140000000000100430006049042809
B2[362] <= 640'h159c2fbffb73ffe0ff80f000007e0000200000007fc31ffffff0fffffe038825f75e45b598161cdcf11692004372f47f7eec4a628d1a7430a69d11830468402ad308010041400c89cc10024a18062700
B2[363] <= 640'h162a8f873ffffffdfffffe0001ff00b026800001fffffefffff1ffdbbf19f00995103e2896de6eac82307e00c3e6f00f1f90c5304320e2545a13db0d4930c722108910800131c208023000c019c71100
B2[364] <= 640'h110423c3fffffffffffff80080ee00306c00008300001e3ffffebffb8380f862e74c21e000252d41c74c8806c335ef8607064be0236183a90cb4c19308098f216040004c009046404204004418420108
B2[365] <= 640'h160003e6fffffffffffff000800000002b00003c00003fffffff3bbe01807f388a1e1941841e905a0e2c8d0efbad47860340e0a5753a07292479203001a246426990000580100300420000c080000300
B2[366] <= 640'h1a00001e03ffffffffffc0010000002050000004803cffffffffbf240fc27f570419259a01029308d8ea260feb6623f6614b72ed2050609914cde0d8c162408c2d8000348801a8019201004081820022
B2[367] <= 640'h3fc22fffffffffc0030000003068000000019fbffffe7f9f689effe7a0c50ad842e34dd90c002a8b01c0364391e152c80329804331411ba009210c824a89801a0810d080814820000043001860
B2[368] <= 640'hc01a597ffffe5ff8c0000f6207100000001061ffffff3ee33a2235a6805381586249c7500405a8c808934033fa4d0990a35209800c1a3e905081a025620000c8040805c0282000000002618a8
B2[369] <= 640'h5c01cc63ff98df9f8000070e05800000000068cfffffe3d8fa08345a116e30d9a2e980083a4c00c800e01f56e28f5096453005981a3e0621658aa238a1000002850445e01808400000020208c
B2[370] <= 640'h18401dc3d1cff3c00000078a031005c001e20077fffff1fc1eed8459d4ad38b4011084c89e432d700103c53593fd42ec211046182b1a40ac4a0e5614d940238e0580002100d800000111000a0
B2[371] <= 640'h950000c00dffe6000000001c0fe007f3c0004f7ffffdffa4d51bd1c0004af01538480cda258f0c0011cac19b2a241b08421c282101ec406e11200042490a02ed280000101c020300002000e8
B2[372] <= 640'hf5c20007802ff9fffcfe072fecfff880ff0fffffffc7f84426dee2101a416c0c50514c084439a781485a741c8901060a02c794a40004a68d01c0c80003480028000000007300000080100008
B2[373] <= 640'h5678280663afffffffe10430783ff1f0080ffffff0fe491208e8480746506a538514c67ad188001c30f0004902002b284006119816578819160000c60008080000000002a1c000000620002
B2[374] <= 640'h607d0800aca9ffffa61400418003ff3f80ffff7fdf9029ba8ec89d01b38693c01a11940500d8003a01f0b18091000a042120099b8246824a010203700862010c401218001a06000020000c
B2[375] <= 640'h580e60000347790000380200800000f3063ffcffe0b001051700481aa10865c880c9142623b3ff230c48ff90121a5a4427a4600386366050471a1180c0212ba0001008201a0000000b0000
B2[376] <= 640'h3030f1e0000864200848000080000000f1f78f000615250c1b00980a008649a3428e98021041dc1d4621a089420248402200e8490c06402380d5800008f92920000008001808000000000d
B2[377] <= 640'ha01fff8c0000274003c000100008003fc007fb8607da5cd8ca6b4183b3d1780010525a120039ef0924de20400424440066e10018404b22b20020992088444c0030044000c180000000008
B2[378] <= 640'h3f0073808670409c000100010000f0ffffffdf6945ad4c96d410c1029490620cb6a19449ff70662bd851600422110822c148362683b014430110840090080100440084180000000000
B2[379] <= 640'ha0000961e3fe997e400002c0313e0007ffffffe1c121583e030028a45e8e0c67871001956bffe0b161989830280000001605280832c0016aa81d41868e0c580000000080000000000000
B2[380] <= 640'h4c0101fee0f1e089fc0003c0ffffd80fffffff649150d850fc052163428900c48a5d2002623fe0b965760090b04000000344b96060049a5612046642240c000000000000000000000000
B2[381] <= 640'hf04001fff01b622a8000389fff1001ffffdcf887a11042069dcbc4693c0a647303d8924943fb81020b2009c0034002018048032a4a488040d0484427818000000000000000000000000
B2[382] <= 640'h380ff80beffe058000001003ffffffffce0effdb7399a3a209e60802bca24e251088820b447a48e049c44100004100c5000b10092f60841118484206200200000000000000000000000
B2[383] <= 640'h1a43ff9003f0bfb00000387dffffffbff061fffe78681ec1b0a2882d493833002580990003eed20040060e08000000034323020986420421880c0200000000000000000000000000000
B2[384] <= 640'h68003fe0805fff80e00168b7fffe07ffc103f68e7c31c819d2dc76e83166410430099802079b00040d700000000000000000207c498000800ce0000000000000000000000000000000
B2[385] <= 640'h340003fffc000ff0f6003805fbf807ff5ffece3e59081c0a211d07d3cc0c01ae52405814030be618000000000000000000007ad05a7324118100000000000000000000000000000000
B2[386] <= 640'h1a0000001cffff07feff0083fdffffffedff6e5648d8c0c6147381035a09c098104058131b9a608001000000000000000000000253276fe484c0000000000000000000000000000000
B2[387] <= 640'hcc000000003cfc07fcfc073d73fffffffff50de80191a0009b00643043174308160420d03000004020000000000000000000022200280c5c3e0000000000000000000000000000000
B2[388] <= 640'h3b000000000009c037f776add7fffffffe0800984f1a8454883612280324040838040180000030009000000000000000180207a520000018000000000000000000000000000000000
B2[389] <= 640'hef0000f0cef020c09fff70fbffffffff2f85c2008c51bb1c12e330602422a900004c222b8f0194080000000000000001e0a527548040008000000000000000000000000000000000
B2[390] <= 640'h780000000000017c700000f7fe007180cb369fffdffffb07db4400440751406563279a082000034401aa4143b400000000000000000006093020827c0c86400000000000000000000000000000000
B2[391] <= 640'h6c00000000000053000000000180000004de83ff8fc84fff7bfa0670093ae529a2a70140000017b4c41c80a232000000000000000000020d51224ebca8bd008000000000000000000000000000000
B2[392] <= 640'h6c0000000000003c00000000000111003e673bebfbc01c17fbf006fa0032ec0000c2b160000000314680000000000000000000000000000ff9e7ee7cdc10000000000000000000000000000000000
B2[393] <= 640'h3c0000000000001b0000021c0f000ffe03ef8f4306302007fbc007e0000042d21946fe000000000000000400000000000000000000000007fbe7fe7c8000000000000000000000000000000000000
B2[394] <= 640'h1000000000000002700057fe17fe007fbf00f7a3f3a06ffc0fc007f800000b5ba4c900000000000000000000000000000000000000000007fff7fe7c0000000000000000000000000000000000000
B2[395] <= 640'h19e00000003ff5f801f000b2000003ffe0fc0073ffffd004e360000000000000000630000000000000000000000000007ff77f67c0000000000000000000000000000000000000
B2[396] <= 640'h6fc0000000000fef002fa6e80070780ff3e80f3fcfdbc0203002000000000000000000000000000000000000000000007c67f6780000000000000000000000000000000000000
B2[397] <= 640'h1610000000160067fe007977e4584803f3600f3fcfefeff5163b00000000000000000000000000000000000000000000fe67fe71c000000000000000000000000000000000000
B2[398] <= 640'h300000000000000d000000003ff00007f80274fa8840009be00704fff6df78360000000000000000000070000000000000000000000001ff57fe60c000000000000000000000000000000000000
B2[399] <= 640'h7a00080060fcfc0001fc8884b08400009ff05fcfffa2dccb632000000000000000000400000000000000000000003010347fe680010000000000000000000000000000000000
B2[400] <= 640'h2c60000000003fc0009fe7f3f8500df9fe07feffb60012b610000000000000000000000000000000000000000002007f33f4680000000000000000000000000000000000000
B2[401] <= 640'h1a3000000000007fff006ffdf0703ffffc073acfc60036b700000000000000000000000000000000000000000000017f33f4080000000000000000000000000000000000000
B2[402] <= 640'ha000000000000007f800006f83f0ffff80332dff7f306b700000000000000000000000000000000000000000000037b31f0000000000000000000000000000000000000000
B2[403] <= 640'h683000000000000000fc00fb83fc38ff801f3fff7ffae870000000000000000000000000000000000000000000003fb01f0000000000000000000000000000000000000000
B2[404] <= 640'h14001f000effff000003fe7d820e70ff00193ffffffa7860000000000000000000000000000000000000000000001f901f0200060000000000000000000000000000000000
B2[405] <= 640'h638030038000e7ff400003e6007f00e000807ff73f64800000000000000000000000000000000000000000000001200130203820000000000000000000000000000000000
B2[406] <= 640'h61c00000000007fff80001d807c008000007fc031c5900000000000000000000000000000000000000000000000600130007f00000000000000000000000000000000000
B2[407] <= 640'hdc0000000000000001c000f2300000000003fc00895900000000000000000000000000000000000000000000010fc01b00035a0000000000000000000000000000000000
B2[408] <= 640'h3680000000000000000100bef80680000001f8000a00000000000000000000000000000000000000000000000007601900026a0000000000000000000000000000000000
B2[409] <= 640'hc0800003c387fe00000003f200f000000189e00000000000000000000000000000000000000000000000000000020190003e00000000000000000000000000000000000
B2[410] <= 640'h34000003e0000f98e00000068030000001e3398c4000000000000000000000000000000000000000000000000003800000287c000000000000000000000000000000000
B2[411] <= 640'h1a00000000000000ecce00012fd00000006b6800000000000000000000000000000000000000000000000000002c000010205e000000000000000000000000000000000
B2[412] <= 640'h28070000000000000000c0fdc4070000014a30400000000000000000000000000000000000000000000000000640000102040000000000000000000000000000000000
B2[413] <= 640'hb0000000000000000000001340c000000cec0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[414] <= 640'h2800000001790700000000050000000001f40600000000000000000000000000000000000000000000000000000000000024000000000000000000000000000000000
B2[415] <= 640'h14004f9072000380407f8001800000000347804000000000000000000000000000000000000000000000000006000000009e000000000000000000000000000000000
B2[416] <= 640'h37e0e001000000000000000dec40000000b98000000000000000000000000000000000000000000000000006e0000000e6f800000000000000000000000000000000
B2[417] <= 640'h15f800000000000000000001823000000024a008180000000000000000000000000000000000000000000003000000007f1c00000000000000000000000000000000
B2[418] <= 640'h5210000000000000000000004000000000a5409000000000000000000000000000000000000000000000004c0000000000000000000000000000000000000000000
B2[419] <= 640'h3700000001ff83800000066140000000003a903c0000000000000000000000000000000000000000000000460000000000000000000000000000000000000000000
B2[420] <= 640'h5003fec3fc00000000000042000000000660c0a80000000000000000000000000000000000000000000007c0000000000000000000000000000000000000000000
B2[421] <= 640'h2be0f000000000000000000700000000003850be000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[422] <= 640'h15f80000000000000000000260000000000780d8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[423] <= 640'he83c0000000000000c000009000000000033d7f600000000000000000000000000000000000000000000200000000000000000000000000000000000000000000
B2[424] <= 640'hb0f8000001c00000000000640000700000df9e780000040000000000000000000000000000000000000000200000000000000000000000000000000000000000
B2[425] <= 640'h6400000000000000000007860000f1000015eb100000000000000000000000000000000000000040000000300000000000000000000000000000000000000000
B2[426] <= 640'ha00000000000000000000007c0173f30006be000000000000000000000000000000000000000000000003f00000000000000000000000000000000000000000
B2[427] <= 640'h40070000000000000000000007873ee0001b1000000000000000000000000000000000000000000000003800000000000006000000000000000000000000000
B2[428] <= 640'h349fec0000000000000000701ff3f19e100c400000000000000000000000000000000000000000800010007c000000000006000000000000000000000000000
B2[429] <= 640'h49bc00700000000000000c00ffc0e101806000000000000000000000000000000000000000000000038006c000000000000000000000000000000000000000
B2[430] <= 640'h1600003880000000000000023f87f82371040000000000000000000000000000000000000000000000020000000000f0000000000000000000000000000000
B2[431] <= 640'hd0000000000000000800e7f00fe18b3fc00000000000000000000000000000000000000000040000000000000000000000000000000000000000000000000
B2[432] <= 640'h148900000000000000000ffc59e27d00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000
B2[433] <= 640'h93f80000000000000000f802fcc00000000000000000000000000000000000000000000002e000000007c000000000000000000000000000000000000000
B2[434] <= 640'h74fe00000000000060000387030000000000000c000000000000000000000000000000000680000000ee8000000000000000000000000000000000000000
B2[435] <= 640'hc8000fffcc000004001f049e00020004000001c000000000000000000000000000000000700000000ff0c00000000000000000000000000000000000000
B2[436] <= 640'h33800c00000080000f8f80000006000c00000030000000000000000000000000000000006c0000000000000000000000000000000000000000000000000
B2[437] <= 640'h1c8000008000001fc7e000000002200c0000000000000000080000000000000000000000440000000000000000000000000000000000000000000000000
B2[438] <= 640'h3600007ec0007e7e8000000000020040fe00180000000004000000000000000000000007c0000000000000000000000000000000000000000000000000
B2[439] <= 640'h50000e000fc87800000000000000140163fff000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[440] <= 640'h14000013e3f000000000000000000003c8157000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[441] <= 640'h5800fe0b00000000000000000000047d38d8000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[442] <= 640'h173f7f200000000000000000000004fc3fb8000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[443] <= 640'h40180000000000000000000000004bc3020000000000000000000000000000000000000000000000000000000000000000000000000000000000000
B2[444] <= 640'h1fe000000000000000000000000009e1fc0000000000000000000000000000000000000000000000000001000000000000000000000000000000000
B2[445] <= 640'hac0000000000000000000000000000000000000000000000000000037000000000000000000000000000000000
B2[446] <= 640'h62880000000000000000000000000000000
B2[447] <= 640'h60ef313e0000000000000000000000000000000
B2[448] <= 640'h7e0000000060000000000000000000000000000000000000000000c000000000013f285d300000000000000000000000000000000
B2[449] <= 640'h7f0000000060006000000000000000000040000000000000000008b00000000002a08174c00000000000000000000000000000000
B2[450] <= 640'h5f0000000000002000000000000000000120000381900000000000480000000710a442c0000000000000000000000000000000000
B2[451] <= 640'h5e000000000000000000000000000000008c00000405000000000024000000009029c190000000000000000000000000000000000
B2[452] <= 640'h3c00700000000000000000000000000000000017c760002c00000000000000000000000f9cc0000000000000000000000000000000000
B2[453] <= 640'h3fc00400000000000000000000000000000000007dcc8001800000000003c8000000000000000000000000000000000000000000000000
B2[454] <= 640'h5dc00000000000000000000000000000000000077c3ba098f8000007ff3c21000000000000000000000000008000000000000000000000
B2[455] <= 640'h5fc0000000000000000000000000000030000003ffecf3ef24ffa0dbc076df800000000000000000000000000018000038800000000000
B2[456] <= 640'h79c000000000000000000000000000003180ec003e7f2bfe7f7f01980b021c00000000000000030010fffffe47fffe0020060200000000
B2[457] <= 640'h7e00000000400008010cf7c0000ff14001803140000a03e0303eeaa819fd3880000001e80013fffc9fffffff677fff0004020200000000
B2[458] <= 640'h1000000000000000000078000000000000363efa1ce0c31bf18000000e400016603f03ff43e50bf530c0000001fe01fffe7f9fffffffe1ffff2000030200000000
B2[459] <= 640'h38000000000000000000000000000000000e3ffe00c8870000000000000000100001fff1f35e0cc2207e003189fe01fffe7f9fffffffe1ffc70004020e06000000
B2[460] <= 640'h70000000000000000c000000000000000000000000000000377fdf3f9b9f95bfb8da74003189fe01fffe7effffffffe1ffff8006020f06000000
B2[461] <= 640'hc0000000000000f700000000000000080000000000000000000000000000003c8fffff70e30eef1febce41380dec01fffe7ffffffffff1ffffec00028f02000000
B2[462] <= 640'h180000000000001f700000000000000000000000001f9f800000000000000001f1fffc1fca0867f80e95770984ce401fffc7ffffffffff9fffffc00008703800300
B2[463] <= 640'h100000000000007ff00000000000000600000000001cc0c00000000000000001f8fff02309043c77e57ffc37d7ee480fffe7fffffffffd9ffe7fe00000783800160
B2[464] <= 640'h8000000e0000000000000007fe000000000000005011424ffc80000000000000000000001e007c2d1c00f0a73fdefb5c9ffeb7c0fffc7f87ffffff00ffc010000007f1000000
B2[465] <= 640'h300000000000000009c0e337e0000000000000007f0000000000000006258d8481800000000000000000000001e00f817e000c83bffed8e31d6fbb7c07ffc7b8ffffe7e00ffe1bc78040fff800000
B2[466] <= 640'h700000000000003ff2ef301000000000000000000c0000000000000000659084988000000000000000000000001f801c0000001f900dcee39db7e13807ffcfb9ffffeff00fff1fe38000ebd000000
B2[467] <= 640'h78e800006001ff803cf0d0fa80000000000000000000000000000000000110c4ec500000000000000000000000ffff00000000001f8b40c8cfe03000007f81f030c0300000010fc00000008000000
B2[468] <= 640'h1c0000033dc00fff49d5d7b6000000000000000000000000000000000011c0cec500000000000000000000001c073fe000000000160a32e008db000003fc1e000000000001000e8f20001c000000
B2[469] <= 640'h1c0003ffe2e427b0c000000000000000000000000000000000011460db740000000000000000000000fdfffc000000000073795c3ffeb80003ffeff03bfffffe03fff8b0ea0000c000000
B2[470] <= 640'hbf0c1ff8001cc2f060000000000000000000000000000000000010c00ddb58000000000000000000000f00ff000000c800008980a9df7a48061ffebf0ffffdfef8079803e0f00006000000
B2[471] <= 640'h1f00000001e123f0000073c9cfc0000000000000000000000000000000000010620d988d000000000000000000000c010f8000f9f6000002f2dffe7e98021fffef03fd78fe7c09ce4b2da40038180a00
B2[472] <= 640'h88c80000cdf840000002118f60000000000000000000000000000000000000106007913e00000000000000000000083f87007ff9ba00000007f3c3fff0020f5d9624f7e963ece1c0380e570733541e00
B2[473] <= 640'hfe7fc0032ec00000010001bf300000000000000000000000000000000000003040039797000200000000000000000c00c79f7ffbbe800000000fc67f54020c2770053f07e80fa0000e11bd0716bf0000
B2[474] <= 640'h33ef8017cc000000000093fb0000000000000000000000000000000000000304000919a00020000000000000000091f3f1f7ffff000000000000e1e5cc2000080003ff8700978030f013f030fe00000
B2[475] <= 640'hffffff6c000000000001b840000000000000000000000000000000000000006000508b000000f00000000000000bf1ff07e7ff800000000000007e00200000602ee0c03f88f8f1942ac6000c000000
B2[476] <= 640'h6ffffe01c000003803e9c000000000000000000000000000000000000000060005e8a220002f80000000000000c07e007b6f0000000000000000020400003700eff5e8101b70601cb6e0000000000
B2[477] <= 640'h1fff03fc40cc00003f8042980000000000000000000000000000000000000000100027bc14000c8400000000000003f80003ffc0000000000000000000000000b2c4ff5360555c071a7335004600000f
B2[478] <= 640'he3000fb031c000007c06acdc0000000000000000000000000000000000000800b00018801b000c8c00000000000000000000f8000000000000000000000000013380f8540fcaf1c79803e90059f50014
B2[479] <= 640'h2003fff01b610000780882500000000000000000000000000000000000000800400007e01e0304cb000000000000010000002000000000000000000000000000ffbfe0dd37007fe3e03da090beb40a1d
end
always @(posedge vga_clk) begin
B3[0] <= 640'h38030008800ffff1fffffefdfffffeffffffffffff0000000000000301e37efffffffbfffff3ffffff7cfee77ffffcc0ff9d1f7ff3e1f0fffffffffffffffffff7fffffffc3ffffffffff7fb
B3[1] <= 640'h38c000000001ff00ffffff9ffffffeffffffffffff0000000000000011e77ffffffeffffff7ffffffffffe7efefefec0ffdffffffbffe37bfffffffffffffffffffffffffe3fffffffffffff
B3[2] <= 640'h40e000000031ff00ff3fff1ffffffefffffffffffd000000000003009ce7ffffffffffffff7ffffffeffff7ef6fefec3ffffe7ffffffcf73fffffffffffffffffefffffffeffff7fffffffff
B3[3] <= 640'hc00700001871fd40ff7fff1fff7ffefffffffffffb0000000000030c9cc7ffffffff7ffffffffffffefffffffffffffffffff7ff7fffff71fffffffffffffff77fbdfffffeffffffffffffff
B3[4] <= 640'hc00780001031fcc07ffffc98fffffefffffffffffb0000000000c18e0107dfffff73e7ffffe7fffffffffffffffffffefffffeff1fffff73ffffffffffffffe7ffbdfffffffffffffefffff9
B3[5] <= 640'hc000000001fd807cfff8f8fffffffffffffffffd0000000000e0c0030f9ffffff3f7ffffffffffffffff3dfffffffcff7f3cffbefff8ffffffffffffffffffffbdff3fff7ffffefffffff9
B3[6] <= 640'hff00e031f898ffcffffeff7fffffff000000000000619f0f9fffffffffffdffe7ffffffffffdffffff58ff7f3ffffeffffffffffffffffffffffff99fffffffeffff7fffffff
B3[7] <= 640'h800000003000010000c0ff8078103f19ffcffffeff7fffffff00000003000c039e0fbfffff8ef9ff9f9f7fffffffffffbf7fff18ff7fcffffefffffffffffffffffefefffc99ffff7ffefefffeffff7f
B3[8] <= 640'hc000000000600000001e7007c0638fc70c37ce1ffffffffff000000000080e01fdfffffffffff99ffdf7ffffffffffffffffec7feffff7fffff7bfffff9fffffffffffedfef39ff3ffffb7fffffffef
B3[9] <= 640'h1fd00cc6000f0feffffe1ffffffffff00000000010007f8f0fffffffffffffffe7ffffffffffffdfffef7feffffffffffffffffffffffffffffffffeffeff3ffffbffffffffff
B3[10] <= 640'h80000000000000000000fc0081008100de7fe3f0ffffffffff0000800021070ffcffffffe7fffffff3fcfffffffffffffdfffef3cffffffffe73fffffffffffffffffff77fefceff3cf99fdfffffffff
B3[11] <= 640'h80000000200000000200fc0089008100defff378fffffffffff0008000200f0fff1ffffffffeff6673ffffffffffffff7ffffffffffffffffffbffffffffffffffffff73f19feeff18f89fcfffffffff
B3[12] <= 640'h848000000004000002007c000800000079c77cfcfffffffffff000c000000f1ffffffffffffeff667bc7fffffffffffffffffffeffffffffffffffff7fffffffffffff7bf31f38ff83f89dffffffffff
B3[13] <= 640'hcc8000000080000000007c0000000c007bc73cbefffffffffff00080000807ffffffffff7ffeff66ffe33ffffffffffffffffffeffffffffffdeffff73ffffffffffff3fe31f380007f899ffffffffff
B3[14] <= 640'hfc0000000000000000007c00000004003f03380cfffffffffff00031000000fffe1ffffefbf8ff99fef13ffffffffffffffffffffffffffffffffffff7ffffffffffff9f9f1cf80007f839fff7ffffff
B3[15] <= 640'hfe0000000000000000003000060004040c0cc000ff77ffff7ff82031000380fffffffffef1f8c3998c3f3fffffff7ffffffffffffffffffffffffffffffffffbff3fff8f1e1cec0013f87b77f77fffff
B3[16] <= 640'hf900000000000000001000000000000103e1fcfb7efff3fbfffeffe0000618077ffffff0982e613099ff9fff9ffeffff3fffffffff7efffffffffffffffffffffffff7f83c990c849f667fb7ffffffff
B3[17] <= 640'hf10000000000000000000000000000990000fc7fffc3effffffeff600004810f7fffffe09866203198ff9fffffffffff1fffffffffffffffffffffffffffffffffff7f0f3c991cff0366ffffffffffff
B3[18] <= 640'hf70000000000000000000000000000383c00c003c0838ffffff7fe20008081ffffffffc08047106166ff9fffffffffffff7fffffffffffffffffffffffffffffffff3fff7e9938cc73ffffffffffffff
B3[19] <= 640'h660000000000000000000000000000181e00c003003c1ffffff7ff00800018ffffffff008006003866ff9fffefffffffff7ffff9ffffffffffffffffffffffffffff3ff0ffff31807fdbffbfff7fffff
B3[20] <= 640'hfec080300000000000000000000000000380800309383ffffffef74300031cfffffdff03e406003c66ffffffcfffffff23fffffd3fffffffffffffffffffffffffff630fffff20fe049b3fbfffffffff
B3[21] <= 640'hfec000200000000000000000000000000386000118c17bfffffef763380383ffffffffc16604800c60006fffefffffff21ffffff3fffffffffffffffffffffffffffe307e76600848e9f3fffffffffff
B3[22] <= 640'hfff300800000000000000000000000200004000000010ffffffeffe23833c1ffffffff800000008000006fffffffffff3bfffffffffffffffffffffffffffffffffffbe0c3660000ffffffbfffffffff
B3[23] <= 640'hfff720830000000000010000000180000004000098030f7fffffff7cc371b81ffffffe000002008080006f7feeffffff3ffffffffffefffffffffffffffffffffffffc07c3668ecc31fcd9b6ffffffff
B3[24] <= 640'hffffcef0000003210cc00082000100002100008000000e7f7fffff3839feff3ffffffb00c08000006881fcff11fffe990f7ffffffffffffffffffeffffffffffffffffff38710001e7f9fffffffeffff
B3[25] <= 640'hffffdce0000000600c8100020618000000000000000001ffffffff7c393ffffffffff900800000000980cfff1bffff990c3fffffffffffffffffffffffffffffffffffff08300e00c7ffffff3fffffff
B3[26] <= 640'hfff7fef8e00000e0ce030012603ce000010000000000019efffeffdf113ffffffffff900000000000980037f0fffffb98cffffffffffffffffffffffffffffffffffdfff03008e08e77fffff7fffffff
B3[27] <= 640'hfffffffcf8000000f7c00012f07ccc00010000000000019fffffffce813ffffffffff800000000000000e1ff0f3ffff88cffffffffffffffffffffffffffffffffffcffc010c0000ff7fffffff9fffff
B3[28] <= 640'hffffffffff000307fff0ffb63ffff3000000000000000033ffffffc499fffffffffffc0000000000000001ff0f3fe7f88cffffffffffffffffffffffffffffffffffcef8808c00017ffe8f7eff9fffff
B3[29] <= 640'hffffffffff00c30fffffffbe7ffff00000000000000000637fffffc09dfffffffffffe0000000000000003fe87ff0370063ffffffffffffffffffffffffffffffffecff0c00c21013fffcf7effffffff
B3[30] <= 640'hfffffffffc00c3cffffffffffefff8000000000000000023fffffff39effffffffffe6000000000000000cfe803f0061003ffffffffffffffffffffffffffffffffecfe0100001013fdfceffffffffff
B3[31] <= 640'hfffffefffc101fff7fffe7ffffffff00000018000080000effffffff9effffffffffc4000000000000000ccf8000006101ffffffffffffffffffffffffffffffffffcfe01c000000f798ceff3f66ffff
B3[32] <= 640'he7bfbfffff998efbffffffdffffef8880000120100000a3f7feffffffeff7ffffff1c00000000000000040004770fc0004ffffff7fffe7fffbfffffffffffffffffffcc08219381df30163ffefffffff
B3[33] <= 640'hfffffffffff1ce3ffffffffffffff1810000100100000061ffffffffffffffffe30080000000000000000100f8308c0002ffffff7bffffffffffffdffffffffffffffcc0821880197cc0f7ff69ffffff
B3[34] <= 640'h3ffffffff3727f0ffffeffffffffe3010000100003000001ffffffffffffffffe1c08000030c0000000040001c31000002bffffffb3f7effffffffffffffffffffffe104801880007c78633f6dffffff
B3[35] <= 640'hff7ffffff3667ee7fffc9fffff3ffe01c000030003000003ffffffffffffffff38cc800000072008000000010e000000039effffff3f7eff6fffffffffffffffffffe10080000001dc0c00ff6dffffff
B3[36] <= 640'hff7fffffffe6feffffff9ffffffbff98c00003000000000f3fffffffffffffff3c00000000c001180000010100000000009fffffffffffffeefffffffffffffffffffc0032c30003cf037fff6dffffff
B3[37] <= 640'he7fffffffffeffffffe3ff7ffff3fffcc4008280000000081fffffffffffffff0300000081e10108000000000000f00000bffffffffcfffffeffffffffffffffffffbc6032c30c67c7c0eeffefffffff
B3[38] <= 640'h3ffffffffffffffffe166ffff3fbffccc00b0c0000099001fffffffffffffff83000000c30300890000c0000000200000bffffffffdffffffffffffffffffffffffff6030620c66f7c004ffcfffffff
B3[39] <= 640'h18ffffffffdffbffffe066effefbfefbcc0092c0030f9900fc7f7fffffffffff000000033f3800c00001340030000000013b7fff1ce7fffffbfffffffffffffeffffff00306480667f00feffcd1f3e7f
B3[40] <= 640'h3bfffbffffffffffff8019bb3f99effffcc1fe0f1ee1fe0080e7ffffffffffff800000003f67ffccc000000000004400817fdf3fc3987ee7ffffef7fffffbffffffffef0c0380698fff17f3e1cf063ff
B3[41] <= 640'h3bffffffffffffff7f8098bb07098ffff31cfffe1807fe0000e7ffffffffffff8000003cff7eefdf0000000000000000003f8f3f3e98ffeffffffffffffffffffffffe41c0f00f98fff1ffff1efb77ff
B3[42] <= 640'h3bfffffffffffe9f7f00009c03067ffff31cfffe383cf98107e7ffffffffffff0000003fe37fc7ff1c00000000000000001f0e1e1f98fffffffffeffffffffffffffff00c0f08f99ff78efff1f3f7fff
B3[43] <= 640'h3bfffffffffffefff800009c3066fbffff0cffff38fc71000fffffffffffffff00000123e3ff1ffefc00000000000000001f0f9c8399c3fff8ffffffffffffffffffffc0c0f00799ff30e7ef1f3fffff
B3[44] <= 640'h3bffffffff3ffffffc00000cc06627fffe861fe71f8e73003cfffffffffffffe000000e3ffdf3ef8c000000000000008000f7fc8c399c3ffffffffffbdffffffffffffc0ff3e039fff70ffff037fffff
B3[45] <= 640'h3bffffffbfffffe61c030000830003fffec31fe00f8f7f0038fffffffffffffe0000087e7ffe3e7fc700000000000000001f7fc03899ffffffffffffffffffffffffff00ff1f019ffff1ffff01ffffff
B3[46] <= 640'h3bffffff88feff660c0480200300807ffef1fffee1ceff0001fffffffffffffe00000c3efffeffffff00000000000000001f33ce1c99fffffffffffffffffffff7ffffc7ff1c619fffe3ffff01e3ffff
B3[47] <= 640'hfffffffffc3ffe66c00000203c800e3ffff1ff7ff0ff9f8001ffffffffffffff0000c3cfffffefff8080002000000000041f71df87d9ff7ffeff3efffffffffffcfffff8fff8739fffe3fffef3c3ffff
B3[48] <= 640'hffffffffffc4fe8cf8840000008400ff79de7ff3ff70310000ff77ffffffdffe000799ffffff7ffe0020108000008000000173dffd57cffffffffffffffff7efff7efff8e7c3883fff7efcfff7fcffff
B3[49] <= 640'hff7fffffffc03f873e100000000000ff6fffffffff71000000ff7fffffffffe70038ffffffffffff00001000000000003c007ffffffedfffffffffffffff7fffffe7fffc7e0f88fffffefeffffffffff
B3[50] <= 640'h7f7efffffff0ff071f1000000000013ffffffffdff730000003f7fffffffffe7003fffffff7ffffe000080000300000000007f7ffffeffffffffffffffff7efefffffffc7e7efbf7fffe1fffffffffff
B3[51] <= 640'h3e67fffffff1f938f08000004000009effffffffff010000007f7fffffffff3c000ffffffffffffe000001103800000000017fff7fc7ffffffffffffffffffffff7efffcc77efbf3ffdf1fffffffffff
B3[52] <= 640'h3ee7ffffff31f931f08000000000008ebdffffffff70800000ffffffffffff3c00ffbfffffffe7f6000000203800000100017fff7fc7ffffffffffffffffe7fffffcfffcc7fffbffffddefffffffffff
B3[53] <= 640'h3fe7ffffff1339c1e0000000000000033ffffffefff8800003fffffffffffff1003ebfffffdffeff000000000000000000009fcfff3cffffffffffffffffffff7ff9fffc9ce3fbffffdde7ffffffffff
B3[54] <= 640'hff7fffffffcf9981c3000000000000312ffffffefffc000003fffffffffffed1001fbffffffffefe002000008100000000018fefff7ffffffffffffffffffffffffffffc9cffdf7fffddffffffffffff
B3[55] <= 640'hef7effffffcf981ce0980000008001b147ff67effff83100007fffffffffce9800c3ff7fffef7f660020400000008000000387f3fff3fffffffffffffffffffffbbffff8cbfe9fffffddffcfffffffff
B3[56] <= 640'hc378dfffff3f6e0060000080c00000869ffffefffeff7000033ffffffffff3f10007ffff3fdf9f798000003100008000001cfff09fff7fffffffffffffffffffffffdffdc77f1cfffffeffffffffffff
B3[57] <= 640'h3ce3ffffffff6e00200600000000000389ffffffffe730003ffffffffffffb70001cffff7fff9ff88000000100000000000fffffdffffffffffffffffffffffffefffec1fffe9dfffffeffffffffffff
B3[58] <= 640'h3ce7ffffffff9801000000030000012081ff7fffffe311e13ffffffffffffe300008afe7ffff9380000000003000c10000073ffffffefffffffffffffffffffffffffcc0fffffffffffffffffffffffb
B3[59] <= 640'h3ccf7fffffff9801802000000800310001e7f7ffff7e1f00c3fffffffffffe000081fffefeff97c0000000001000008000073ffffffefffffffffffffffffffffffff8c07cffffffffffffffffffffff
B3[60] <= 640'h1f7fffffff98009803000001008c870067e7ffff7e1c00c3fffffffffffe000003fffedfff97f300000000000000800007e7fcfffffff3ffffffffffffffffffff7dc17effffffffffffffffffffff
B3[61] <= 640'h813c7ffffffffd001800000000008400001fe7ffeffec8803ffffffffffffe8000033fe7dfff37710000800400001800003fc33cffff7df3ffffffffffffffffffff1fc1fffffffffffffffffffffffe
B3[62] <= 640'h3cffffffffee01100000000300000002997377fff780807ffffffffffff88000083fffffff36600000000000001000001f877fffff5757ffffffffffffffffffffdec0ffffffffffffffffffffffff
B3[63] <= 640'h1cffffffffffe7c10006008000030000009831737eff0000ffffffffffff780c0001fffffefff6fe000000f080009000000f3ffff7ffe73ffffffbfffffffffff7ffdc003fe1f9fffffdff7fffffffff
B3[64] <= 640'hdffeffffffff7fc0000e208018008c06000001eeefff880107fffffcffffc0c00010ffff4ffff1f0008080070000c0000003feffffef7ffcfffffffffffffffeff7e9087cf7ecf7fffffffff3fffffff
B3[65] <= 640'hffffffffffffffc0f00e800800000c8600000006ffff880133ffffffffffc00626007ffffdffff0100000007000144000000fff03ffffffffffffffffffffff07f7709878effffffffffffffffffffff
B3[66] <= 640'hffffffffffffffe40004000f0000038200000000ffff8000fffffeffffff800e47007effffffff0100000007000124400000fff03fffffffffffffffffffffe07f67800e8ee3fffffffffffffffffffb
B3[67] <= 640'hfffffffffffffee6000000810000013000000006ffff80027fffffffffff803878807effffffffe000002007000060400001fff0ffffffffffffffffffffffe03f63f01c5ff4fbffffffffffffffffff
B3[68] <= 640'hffffffffffffff768000008000000012000000273fff80023fffffffffff800038886effbfffff060000e002000070000001fffcf8cfffffffffffffffffffe00f63175ffffcffffffffffffffffffcf
B3[69] <= 640'hfeffffffffffc7760000c11000000083000080223ffe40003fffffffffff80001d087effbf7ffc2e00000002000072000000fffdfcefffffffffffffffffffc00060669ffffeffffffffffffffffffde
B3[70] <= 640'hffffffffffffcf76000001190000009000004022fffe40003ffffffffffe00008b01fffbfef0f8e40000000000006e400000ffffffeffffffffffffffffffffc0060e48f7fffffffffffffffffffffff
B3[71] <= 640'hfffeffffffff3e7200011c3800011e1000006076ffe640007bfffffefffe000081039f38be8178e60040010000000f411101fffffffffff9fffffffffffbfffc0060278731fffefeffffffffffffff7b
B3[72] <= 640'hfdff7fffffffff0c008066c6800001000101060ef3fcc0007ffffffffefe000100c03b703f20ccf8000000008000719c0001ff7f3fffffffffffffffffffffdc30007bfc73fff3fffbffffffffffffff
B3[73] <= 640'hfffffffffffffcc0c4007cee00000000200000037ffe3c007ffffffffffe300000303b000020000e00000100000076600100ffff7fffe7dfffffffffffffffdc30007048d57fffffffffffffffffffff
B3[74] <= 640'hffffffdfffff7cc000007eff00000100000000137fce38007ffffffffff871e0033a208000000000000001800003ee61e3a47ffffbfff39fffff00fffffffffe030000008c10ffffdffffffffffffffc
B3[75] <= 640'hfffffffffffff81c8000e7ff80000100000c6103ffefc100fffffffffff07ff8001a0080000000c000001c800003ee41c18c7ffffffffcdfffffc0ffffffffff0600000004008ffffffffffffffffeff
B3[76] <= 640'hfffffffff3ffc01800000fffe0008000c00c6107ffffc100fffffffffff8defc000e00000000000600000c8000007f0c00083fffdffffcfcffff8003ffffffff8000000000007ffffbfffffffffffeff
B3[77] <= 640'hffff7ffffbffc1c01c003fffb8008000001c000fffff7c007ffffffffffcde7e0006000000000004000087c00000778cdc103fffcfffc3e8ff7e0003ffffffff0000000000007fff7bffffffffffffff
B3[78] <= 640'hffffffffffffe0c038203fff3c0000000038000fffff7c007ffffffffffc7ffe000f0403000000e0000007f08000fec0c0011fffffffc38fff7e0001fffffffb000021b20000ffff7fffffffffffffff
B3[79] <= 640'hfffffffffffff8000060c1ff3c01000080318037f3ffff007ffffffffffd7bf000330000000004070000bff00c03fee0c0011ffbffff3e0fefe10001fff0ffff000033b70000fffffcfffffffffbffff
B3[80] <= 640'hffff7ffffff73c800361ffff5fc0600000070046c7ff7f007ffffffefffcc680000000001c000718000619c40019ff9c7c8087bfffffc6c1fe0c00003f997ffc8000c3ff0000f7ffe3f6ffffdffffce7
B3[81] <= 640'hfffffffffffff00800607fffff000000001e000406ffffc13ffffffefff0f000000080001e000798000011c6003fe7c776000fffffffc7c1fe8000003719fffe00007fff0000ffffff76fffffffcceef
B3[82] <= 640'hffffffffffffc0180060ffffff860c00003e008000ffffe01fffffff7ff0180000000001e3e00ff8000002c2003fe7c1e6001cffdfffc71fe780000473207fff00003fff8000ffffff67fffffffe8773
B3[83] <= 640'hffffffffffffc0000380ffff5ff00800800f800100fffff00ffffffffff0000000000019e3301eff800026c2003ff81ce400087fffffff3fe7800006036600d700803fff80017f7ffe66ffffffff027b
B3[84] <= 640'hfffffffffbf7fc800180ffffdff0800000cf800001fffff01ffffffffff000000008601973003fff000006c000e7fc1cdc00007f73ffff3ffe800000036600100000ffff80013e7fe0e0ffffffff08f8
B3[85] <= 640'hfffffffffff73c0001801fffbff0000000ff8000000fbff81ffffffffff0e0000008000131803fffe0100e6000e33c81188001ff737fff3ffe008020010000000007ffffc0001e7fe5e0ffffffff1cfb
B3[86] <= 640'hffffffffffff3c00cbc03ffffffb000001fc800000061ffc1ffffffffff8f0000008000000803ffffc011c3000620800000001ff8f7ffbc7fe00830300000000000ffffffc00047bf002ffffffff8323
B3[87] <= 640'hfffffffffbfe008001d8ffff63ff400001ff802000001f7c1fffff7ffffc700000c8800080013ffef0011c30002003000100009d8ee3fbc3ff830c0000000000000cfffffc80060ff807ffffffff8723
B3[88] <= 640'hff7fffffefccbf8107e4ffff0fff010011ff9800008efef83ffffffffff0f8000104000030007ffffd000681000000000000000ff6fffffffc4118e0000000000021fff3ff8001661800fffffeff0040
B3[89] <= 640'hffffffffffdcb38003c4ffffefffe00039ff810000047ff81fffffffff207c00800400000000ffffe780000000000000000000c026fdff73fc000f000000000000307fffff0000070000ffffffff00e0
B3[90] <= 640'hffffffeffffe92000061ffffc7fff0003fffe6000000fff10fffffffffe0e000080600000000ffff77c0000000800010000000070200fc01f0008771000000000000ffffffce00010000ffffffff2160
B3[91] <= 640'hfffffefffefe820000e1ff8f07ff20003fffe6000001ffe003ffffffffc0e400000000000001fff398c0090000c000108000000fc0000c21f1003df1000000000000effefffc03000001ffffffff31f1
B3[92] <= 640'hffff2f7ffee0be7801e1ff8e03ff01007fff6e00006378c003ffffffff0066000100e0000001ff71ffe0800080e00003c00000f881010c2141003ffd000000000001ffffffff380000007fffffff60e3
B3[93] <= 640'hffff2ffff7e0bef00101ff8f01ffe700fffffe0004f7f9811affffffff183f003e00f0000001ff79fff0000003ff00037800007801010e0760007fffe000000018007ffffffffc0000007fffffff2063
B3[94] <= 640'hffffe6ffffe1b7c00101fe8600fffe71ff71ffc406ff99000fffffffffe9b800800030000000ffe03ffc800003ff00ff7c00000710000e8e3000f7fff8000000300c7ffffffffe0000007fffffff0003
B3[95] <= 640'hbfffeefffef3b7e08190ff8401b9dc7dff017fee047f9080cffffffffdc41800001800000000ffe07f7e010000ff3ffef60000e0b8008e8e700737fbfe000080031cc3fbefffff9800007fffffff0001
B3[96] <= 640'hfe4ffef3e6cffefc0080ff04011ffb3f7cc01f30003f8006cffffffffff800000001001000009fdb1ffe900746ffffff7f00001e2021008f7907fffde0108c000088cef731ffb7d819005ffffeff0300
B3[97] <= 640'hffc7fffff7efffff0000ff06003fffffc3009f8100bf00028ffffcfffff907000100000000009fe01f7fbefe07fffffffe00040e0030009ff903ffff60010000000e8ff008ffbff839007ffeffff0000
B3[98] <= 640'hffffffffffffcff38000fe000030ffffc000ffc311fe00031ffffcff7ff70000010100000000fec11f3ffffe9ffff1fffe0006630030003ff103f9070003300000073ff08c7ffff871007efeffff0000
B3[99] <= 640'he7ffffff99ffeff30000f8000001ff7ff003ffc01fff0003ffffdfffffe30000180310000000ffdf1f07effff9ff0070ff800e731c20c03ff103ff279801180000ee7ef0803ffdf970009efefffe0800
B3[100] <= 640'he7ffffff9ff9fffb0001e0010807ffc47901ffc10ffd0003ffffdffffff80000002b7e00c09ffff807c3effff9fc003003e00c7f3fc3c07ff103ff6699000c80003cfff0003df97970000ffffff00100
B3[101] <= 640'h7fffffffbff9ff7e0001e0031807ffc00000ffe0cfe80101fffffcfffff800033effff3064bfff980710efe7fff8000007f0007f07c707e7f0037f7e10000c80813fffc00038717ff00007fffff08110
B3[102] <= 640'hffffffffeff9fe7a0001fc000007ffc00000f800ffe8011bffffe8fffff801037ffffff864bfff190600edc3ffc000000ff800ff83ff0767e00007ff20000000833ffd000000607df60033fffee28100
B3[103] <= 640'hff7bff7fc6fb8ef30001fc00e087ffe10083f804ff60011fffff0effffc01001e7ffffdfc3bfdff96603e00099c0000004fc00c7e7fcc077e040079b76e020000ffff0007000647df60071fefc0f0900
B3[104] <= 640'hffcfffffffff99708189fc000001fe711027fc19ff2001fffffff3fef6803883fffef1fcfeffe7c1630001806c800c1100fc01ff3ffff27fb20007fefc00000e0fff00840f00f0cdf3004ffffc3800c0
B3[105] <= 640'hfffffffc7fff8920800df800000ffff11027fc19ff800087fffff3feff8008b7ffff07fcbfffe7ff0708010041001c00007e00fffffff03f120001fffef000037ffc0000e000f1fbfb00effffec100c0
B3[106] <= 640'hffffffff7fffe620000ff800801fffec003fa01ffe80841ffffff3ffff10ccbf7fdfc4febfff7fdc0600000041003980003e803fff7ff2ff000000ffffff00e3fe00000001015ffffc006fffffc10080
B3[107] <= 640'hffffbfffc7ffe600006efc00801ffffc003be00ffc0000ffffffffffbf10febf7ec0c07fffff7fcc0000c000400019e6233e800ff773b7ecb000017fff1fccf3fc00000000c3cffd780069ffff380280
B3[108] <= 640'hfffffe7ee7ff6e000064fc00881fffff001be007ff000107ffff7f7f9801fffde080001f7ff331c0000fe00040001de7701f8007fff3bf06b000017ffffeffff7000600000ffcffcf18069ff0f180380
B3[109] <= 640'hff7ffe4e7fff0c0000c538000003f7f30003e007ffc001037bff7fff9001fffcc000800f7df10080003fc00010019df3fe0f80077ffff600020000ffffeffffb600fe00000c7ff9cf1007dff07c10380
B3[110] <= 640'hffffffff1eff808000493c002013fff10007e007ffc0000331ffffff121bffff0000000e4101010001fcf8001003b9ddff6fc000fffff2f0830000fffffffffe003fe00400ffffc071004fffc7c103c0
B3[111] <= 640'hfffffffc03ff802000097e7089ff66f0207f0127fe38000300ffffff361fffcd000e20000104010001eefc80423ffb5dfee7f000fffef73f83008737fffefdbe83ff400401ffcf8138010dffc3380300
B3[112] <= 640'hfffbff7099ffc020100327edefc881f140673203f9f8000162fefbdd1e83ff7c0000000000000c0637fb61012071f9f3cfc3cc009efe73862080c2fbfffefffe83ffc001001d7f180000ffff3f980000
B3[113] <= 640'hfffffffc11ffc012080007ff7fc0087b206730017dfd800003ffffff3c0fff600000800100010c2ffdbff800001ffff3ef87ff90fefff4f6200003ffff36fefc87ff000103fcf80080003bfffe800000
B3[114] <= 640'hfffeffce33ff019704000ff7ff80001f0cc336817cffc00001fffe7f7801ff600001c0037bf88eefbcbffc00081f86ffef07fff01ffffea2000003bfff337c3807ff381ff3fc002000003bffff810000
B3[115] <= 640'hfffeffcc63ff019f06000ff3ff00341fc081bec07ced060009fffc7ffc06ffe80713803bffec8fefbcbff8000cff02ffcf077ffe1f3f1f03000003ffe01303700ffff01ffbe800000000fffcff810000
B3[116] <= 640'h1ffffff887ff8c9604009fb3e2003c19dc89fffc6f3f6400097f306ece0ffffc00b9003fffe3ffffff3fd83c07ff177f0fc37fff797ff103000003fff08003f01fffc03f7fc0c0000008fffdff000001
B3[117] <= 640'h7effff300eff9cb600001fb68000e301fc01fff86f3ffc0088ff204ecfc3ff4c0499403ffb02ffffbf33f81e07fe807f0fc17ffe73fff122000003fec00018601effdc3f7fc0000000001fffff600000
B3[118] <= 640'hfcffff0006ff87b200001bb20011fb80cfc1fff80cbfff6000ff0067fff0ff780f89001ff003ffe7a002fc0e67fc0c7e7e81fffe07ff1b82000003efc00010001ffff92f99c0000000008fffff608000
B3[119] <= 640'hcf9fd80087ff0332401c19b30061fef90fc7fffd29bbffe004f8cc737f707f710c8f040fc018f0e7e0787c1e66fb8cf9460038fe00ffb88610010339fc1001009fffc0099900000000008f7ffce08000
B3[120] <= 640'hfcfefc00827f867900033e9200707ee00fffc1f9e0c0ffe0001c747fe7e07e880130003f809063e164c0d91e9ef81c39e64272fea2339800010000f03fc680821ffec0391986000600460ffffffcd000
B3[121] <= 640'h1cff3e0000ff8000000067900020e3f306bf1700d8007ff014c7667f7ef03ff80100100f801103e001fcf83f9ff888386e4002ff82339000000001001ffe0084fffc933b1980006600e603ffff8c0000
B3[122] <= 640'h1e0f3c0480ff90100c016330000003f006b8bfdfaa0060301cc3747ffefc1ff8080110078023803003fc783fbff000780e0903ff403280000000010003fe03c47ffc13f10000004000e703ffff8e0600
B3[123] <= 640'hc600c006c1fcd0000c202032000000000781fbf06cffc1003f74f47ffffcdf380801107f0021000003ff3f0fbff880f80e0f037f609201000000000f02e3f3013fc003f000010100200203ffff006000
B3[124] <= 640'h80000306c1f8c980771c2037181c010f0020bfe6e300031fffffffff7ffe8f000000367c0cff70007fff3f0deff9d0e802e8167fec0200000000000f0001fb19ffc003f000010003308fefffff706000
B3[125] <= 640'h680f87f8073c0081781c0800000107fee28011c3fff1ffffffffe0fc00000fff81dfff800677e3ffbffc1c3e0006d10fcfc03c0000000801e8106fff07fc003fc00010039009fcfffff710000
B3[126] <= 640'h8e90fc3c307fc31c0681000100b001767f28000cffff19fefffffe83f90030fff9ffe79c1067fe3ffbffe003a8005f00e037c200000000003fdd863f3c00808fe0000000f9069fcfffff701900
B3[127] <= 640'h188f1fffe6f3ef30001168ff8fe3881753920388177e1911ffc7ffb83cbe1013fb4fee01ef07fcf3ff9ffe37e9d00fc0080a3c180000000003f9c00317cc1823fc0008003b987998fffff8e1980
B3[128] <= 640'h8000839cf11e3d5effdfff64037ff57bdce0f9fcf0663379cc06cfff7ce7c07df608bfc37c003f9866c61f7ffd90d4bf00c000013061e5000c1e000fff00079e990f3f990c000107e00486ff79802000
B3[129] <= 640'h1cffd81f003efdffffff7e0003f6f5fffd61f1ff320630ff0f04fff78047c00ff21ffde1f8000f9864fc3ffbfdd9ffefe1000103707ffe04009f0003f802869e800ffe190000000f010c03fffb800000
B3[130] <= 640'h3fff1e3fa167fdfbfff83f8021fcfe9f79f1fe7ff60010fffe807d718147f80f601fbfe0f8000fe124303fff3df1ffcff80001c7fc3bbc0600c300e37002001f80ff3e1801000038030021ffff800080
B3[131] <= 640'hffff1ff7f16f3ff9fff8338470ff7c103339ffff7e00017ffc807ff21c0ff87760ff3f01fc00078100203bfcbdd07b4df88001e7ff9b0ceecdff00614082021b00ffcf98f0009000008101ffff800080
B3[132] <= 640'hfaffff67307f1f9cefce03c07ffb180000097effbfc001ff7fc04fe63fffe0f3eb7fe9017c00060c00203b7ffdd0fa08f8e07fe6ffc0006ffdf980308100001bc779c30170001100008104ff3c800000
B3[133] <= 640'h8e3ff33e307f879cc0cf00e0dff190000081fec7ffc4e3fbfffccfeefff9c0f31f7f48003e001e0c0000837fffffee81e378feffffc1003ffdb8880080000019fff9fc810000000100100cff3c801000
B3[134] <= 640'h84fff7fcb09fdd6400cf9e20fed1f001101cf9007f80ff12f8ff6ffefffb03307fe2480c1f003e1f02fefff0bfffc001e37be2ffff71f00037f9010000000001fffffcc000000100002002fffe801000
B3[135] <= 640'hfc803eff338fbf66007fcf00ff9df00180c081009c5a8039ffff7ffeff7f03117860c0801f00fe1fc7f1ffe01bff980df8e201fffc769f0483fff12000010001fff9f304c4330400814831ffcf801000
B3[136] <= 640'h78797bffbc26fc20111983387fe6f8010c73801600210117fffff9f3ff8c6c00208c3c1c8fffe63fbbfff3e09ff7c106f17e01fff6501fffe1fff1000004000377fff180ee61000018000f7ff9e00000
B3[137] <= 640'h61070ff3fc87ffc0011807c17ff71803c0f00036003cc0023fffffdfe3807fc1ed0df8c787ffe13ffbfff7e01fff010ff93801fffe00011fe07ffff00040000077ffbf06de0f0000000002fff9e08000
B3[138] <= 640'he1008fb26006c18080000c83d9fffc0fc0cec73e0007c74033ffff03f0007e01fc1ff3e6c79fa07fffcfffc01f9e011f7810009fdc1c800fe000f3f08000000031ffbf071e4c0000200000fff9e0c000
B3[139] <= 640'hf9418b3ee00000620000800099ffec1e8f8ffe3e0017fc68317f191838001e00fc3ffffec79f00fd7f0ffec00f7e00ff38f0001ffd18800f628033fcc00000000f3fe1071ecc0003000007ffff1f8000
B3[140] <= 640'h7c021b9ef8e280e20f80800199ff061ffcfcfe9e7016e47f00ff111030001600fc1ffeffc3fe81d87bc09ec00fff00fe007c007f7f0886fe37fc07ffc00000030bfc61861ccf0006000007ff7fff0400
B3[141] <= 640'hcc0031c0fcc007fc1c9800001bffec0f9ef9c1867003ffffe03000800101f307ed1fffffe1fc0f88f9c09ec007fce7fecf6c007f6e0377fe7ff003ffe000000300ff73c4997d000e0000037fffff0e00
B3[142] <= 640'h4c800080fe04073939980100037ff80f1ffffb0000069ffff00000000003f30fccf9737fe1d86f80f9001fc00778ffffef68007ffe034fff7f7a01fff800000046df7e8f99fd0026000000fffffc8c00
B3[143] <= 640'h7d881414ff8107b9f1810000003f190fefe7ff3000069fbff0004108008f6e8fece97303fd860b80390013c002f70ef30cf0011fe600071100fe98fff882000046ffc60f990f0043302000fffffcc000
B3[144] <= 640'hfe6100000760067fff26010c84800207bfffce08618526837d0002018300bb077cfe11733e03f88280088042417f8bcf065ac6be7d017e80889800ffd020000071ff8f00e60e18800683003ffff9630c
B3[145] <= 640'hfee0100003fc67df3c068080fc00008f1fff0edb608100007f80123f1022bbc7eff800313bfff18106800800003fffffc07f7fbe7c03c8c020000fff8920000071f89c00646efc007fe0000fffc33804
B3[146] <= 640'hfff8100899b80f8c1802c0c17c010082bfde7f7f003f00002c80923ffc00bfc7fff8000001ff800000000400181ffffbe1f973fc7c03c00000000fff9f20000077f8cc002060c7617ffe2003ffc338c0
B3[147] <= 640'hddff1000d9f20188810000017b010003ff1c799f80f3600066c117fefc00bf87fff8800000f180c0013c9180b804f9f00ef9f2f87e30c00040017fffdf20c100cff8c003007007f3ffff6401fffce1e1
B3[148] <= 640'hffff3307dff380c0010021000e0008011c0c4dddf9e7e401f78017cfff10fd00ff989f0000f1800ffe11f9821100b0000c0102001f3be000cc83e0fffec400000e000000009effdfffff6601ff7ee7f1
B3[149] <= 640'hff7ff0c3fffe01e1000020001c800003bc00cddffbffc501ff80b60ffe10ed00b800dfc30033080ffffff9b701001004000108000f83e103ffe3f0fffecf000806001c00009f7fffffffee0dffff7e71
B3[150] <= 640'h803ff2f76ebe0700000060000ee00103fc00cc1ffffecc013ffcbffefe11cd000105e4c00009005ff87efffff08c810020000d8801c1f001fffff9fffec7c0000000180000191fff190ffc01fffffc30
B3[151] <= 640'h8031ff7f669fe0000100c00007f8010338000c7cffff7811e3f81fff7f9fc98100086419069c804ebf6f9ffefe8f1bf0c600099900fff8003fffffff7fcf80000000c1000031ffcc39017c013fffc008
B3[152] <= 640'h89ff3ffff6d810010011002770000f7810411b73f47c84deffe6ffff1f410100836d8080fb610ffe86dffbe707e3ff00c83b8fc03fe0007ffffffffcf3e0000800800004ffff0001017f807ffffeff
B3[153] <= 640'h13ffffffef81000000000037f400ff8900007413fe20ffeffefffffe7f80606007c800ffe607fce029fffe70ffedf0f40fdf03edfe0003fffffffffffe00000000000001fff000101ff807ffffff8
B3[154] <= 640'h1001f3fffedfe100018010007ff4801f9908000c0bf6007fcff6ffffff1fc0700007c01077ee07fce029efffffffaffff69fe73668461c0819ffffffffccc03000000000007fe000000fe01fffeeffc
B3[155] <= 640'h8800fffefe16602000001000fff4801f13e800080fd7c03ffff47ffff78bc0601016801016ee07fde92cfff7edefffffffdff73e23c20fc000ffefffffce800000000000007fe400000de013fffff1f
B3[156] <= 640'h18c001ff8741660203000088067d481ff3be000100fc7c017bffffffff799ffec00040000006e27ffff6cfff78840fffffff7ff1e7fc001e01005f3fffc570c00000000000077f400081f6801ffffe1f
B3[157] <= 640'h981001e3808660383c0001d0379ec1ff0d30000017d4f807bfffffffee39f7fe00c40008007837fffb67ffe810001fffff7dfff7f640003c1601f3bffcf710000000000000f7f000081f6c07ffffeff
B3[158] <= 640'h9b27000400006f83fffc010506ffec0ff0d30004017fef86737ffffffff2077fff3c4000c103837ffeb27ffe8030707ffff31dfffdf3010700603feffffff80300000000001ffe8000017f01dffffffe
B3[159] <= 640'h18f0800080087f83fffc007a817fed0ff83ee01e80fffe92e17ffff6fffc337ffef34c187374877ffcf267e400707007cf82193fdfdf813e3d761ffffffef8000000000087fffc8000017f600c7fffff
B3[160] <= 640'hcf8402100073f83fffe000000be7187c001703c001fffa88ffdffffffbee1eeffe0f8b83fff1ffc66e79fc80200f03fc9801c7eeeffc0ffcfc318fefffec01800011000003fd80e0000ffe0077fbbff
B3[161] <= 640'h87f8400801061983ffff8000016ffe87c810f1e3800ffda8007ffe7fff7f7ceefffde739ff1f1f1ff7f98ff93700f03f3b8000ffbedfc0dffefc0197ffff80000000010000fff80000003f00007ff9ff
B3[162] <= 640'hc7b84c0801221083ffffc000004ffe07e018e3c18007ffe801ffff7fffff3cfffffffff9ffc77f0fbb3901f016c0f03f7f8003ff77ffc1fff8f80107ffff80800000010800fff80000009f80803ff97f
B3[163] <= 640'h6e1b6c0110000081ffffe100600ffe076001c3c08007ffea03fdffffffffcfff7fffffffffff7fc099190170008071f9f3c01ff97eff013ef3e080037bff888080000000003ffc8000008edc003fff7c
B3[164] <= 640'h7e83fd0100000000ffffe000607fff07600003000007ffea206d79fffeffe3bbffffffdfff7ffc069888017c000021e97fe03ffbfe7e487fefc0c803f9fff800800000c100fffc0000008f0cc33ffffc
B3[165] <= 640'h6781cd80810000007eff980000e7f902e01800000007ffeb3049ffff3f7ffb99ffffffdfff7ffc04fccc01fe4c30010fffe07fffffe00c831e004011fffffe240000c20000fff40000001fc4033ffffc
B3[166] <= 640'he391fd80010000277eff8e008001b802c1000030000fff297000ffbf7f7dfc01fffffffffff7ffc06c64007f6ff801bfff603fff7d00000338010010fffffe640000c0300339e41000003bf8073ffffe
B3[167] <= 640'h62bffd1c18800087ffff840098781006c900002130e77e19fc81f73fe6f9fe70dffffffbfee7f80004a6001feffe19ff3f060fffe1001e8021c000501dfcffeee000010003ff06000000c2e3803ffffe
B3[168] <= 640'h9c6fffc000643007ffbfff60c1006400e0000031ff7fffccf101ffbfccfff9fcffffaffecfbfee0140000081feffff7fec00efee60001f80208198019ffff7fe8000000407fff600000001e1c03ffff8
B3[169] <= 640'h83fdffc000fe080efff3fc2306002400e300001bfffffecdf08070dfffc0fffcff7ffd7f8f72f00901000003dfc7fee14c007fee00003fc300119c801fffff3f800000000ffff600000007ff08039ffc
B3[170] <= 640'ha3cdffcc1ef88edefff3fc2202010400730301ff7fefffcdfc06ffdfefe07fffffdffdefffd7f148000001010f87b2c04c003dfc0011ffff8018c4800b7fffdfc00000000fffff00000007fe08038fc1
B3[171] <= 640'h770fffee1ef98effff39fff0e0000604717f81ff7ffffffdfc073fffeffcfe3fffbffde7ff9763400300090003f09004040039c0003bfffffc9fe480005ffffcc00000003fffff00000000fe800c07f0
B3[172] <= 640'h764ffff203fffffefe9cfffe34000200787ed93f7ffff9fcf003fefffdfcfe3f7fffd9ff6efbf0c01000010871f880040003fbc0000ffffffedf660e005efff8c00000003fffff00000000fec00003f8
B3[173] <= 640'hf2fdff6303ffff7ffec46ffe3c000000fce7d9ff7ffffffc7006e7fffdfc3ffffbfff93feffaf8400000010c7f7980000003e780180fffffffff767f800cffffc00000007ffffd800000007f300303fc
B3[174] <= 640'h8279ff7003ffff6fffc807fe700000009e679ffffffffffdf01fcfff7dec1ffffffffc1fbcbf7b4002000009ff7b010800006780000fffffffffb8a28004ffffc00000607fffffc00000037f300103fe
B3[175] <= 640'h9a61ff7e33ffffffef3838fc638004009e779fffbf7ff7e9f81f3eff7fefff7e89efe77f7cbbf80880004001ffff018080006990803e7fffffefff000004ffffc00c006607fffff000a407ffe3803ff3
B3[176] <= 640'hf973ff7f36f9ff33ff40027f731c02000b9863ff3dcdff77f81fffff7fff7f7ffffff9ffb7cf20008000080fe73c00c100036fc00204fffefffcee800e81ffffd90104990e7f87ff300007ffff800379
B3[177] <= 640'hbf79fc7f67f8f0f1fd0000e773cc00037f0f70cee04dff0df80effffffedffbfffffff1fb78760000100003fffff00000001ff002000ffffffffff000081fffffdc006bf0cfffffe2012cfffff0083ff
B3[178] <= 640'h1d383ceee7789df1fd0000e7e7c400007fc620cec1006fc1c00fffffffebffffffeffffff20000001800803ffff800000001ffe02003ffffc0c37f000000fffffcce67ff82fffffc0002cfffdf0087ff
B3[179] <= 640'h988001ce27f09f1fff00003fffc79000ffe68009010002e1c03fffffffedffdffffefffff0c000003800013ffffc00000000fff80001ffff00007f000000ffffffffffffebfffffc0012fffffff01cbf
B3[180] <= 640'h8180808f67e0800ff7000018fefef1e3dc6f80812600037a803fff7fffecfedffffefffff2c00000f000003fff3f0000000073fcc000ffff0004fcc000003ffffffffffefffffff800bffffffd4003ff
B3[181] <= 640'h8100789fe3e0880ef0000001fefe1bf39cfe0101e6800749007fffff7ffcfffefbdfffffb70000016300003fffff4001000603fde0407ec70082dc0000003f3ffffffffbffffffc00016fffffce003ff
B3[182] <= 640'hc1001099e7e01b04e0000001fffe9b709bf80101c09000c0803ffffcfffdfffeffdffe7f360001216300000ffff8400000e60fff6c4000800000980000003ffff9fe7600ffffffe00102fffffce001ff
B3[183] <= 640'hf83003b93cf00001f8000018fcfefbf1d2db40a181160001803fff6fff7bffff5ffffaffb0070121600000047f1e5018c0e39fff7d60000800a0100000003fff81016000cf9ffffc01bfffffc74000ef
B3[184] <= 640'he0010086c6f0000cf20800001df9f7fc98e7422684f8000102f9df67f7cf7f3fef7fffcff230860f9c406023779f00000698fffffe1c00800000700001003f8300000121303cffc09876ffdee78000ff
B3[185] <= 640'h1c06fc000cf0000000197feff81fff00e385f8e398007b7feffdc07ff8feffffff7c00103c9f4000033fcf000202bdffffff1f01180030200000037f9200002ff00111ffc099e7ffffff8018ff
B3[186] <= 640'h100001c00ff0000b0000000093ffcec1fff40e30fffe380004fffdff9e0fffefecfffbffc0030f89f4080007ec78020e3ffffcfff87811e7c7000000003ffb000003fff18003ffc1fdffffbfc00187f
B3[187] <= 640'h100008100f30700b0000000011b3fce00fbc0060ffffff9006fffdbf9014fffffdffe9fff0012fc9d41800c7cfe80e061fffc8ffffeffe6fe00000000ffff9000003fffc00007f89bfdfffbfc00093f
B3[188] <= 640'h8000008100f18000b000000000193ffe03f9c0864fdfffff906ff1fbf800cf7cfffefefeff001fff3848080c1ffc800730ffffe3ffff3fe6ffff000001ffff8000006ffde3c0033bfbfdfffdff00033f
B3[189] <= 640'hc3000000038c1e0f0000000000077fe033d4d064ffffff8907bff7fe000e779fffffffbee011fff3840000e173c800610f7ff630fff7ffff8ff0000033fff80000007ffffe00003b9dffffed800033f
B3[190] <= 640'he200000003e87e1f00c01000004e7ff001ccf7cd779ff7f907fffffe0c0e607ffffffffe6013efff1404000f0be0344007fff0307ffffff3cff060001ffff80000007ffffff803339e7ffff980001ff
B3[191] <= 640'he0008000263ff0e1f00c800000046eff60c7eff8f7bf7ef3915dfffa200002c0fef7ffce7f8032ffe1401801018f000c003fffe00201fc593eff060718ffffb000000fefdffe8071397efffffc0000ff
B3[192] <= 640'hf00404000f07fff3f801200000001f738101fee1ffff7fff7c3f7ffca0801cc107fc38200f604cdf0088060303082084b031f49000e138ff797fe3fed2ffffc8000001fffee3c0882e0fcffc000081ff
B3[193] <= 640'hb00606000f0ff93afc0000010000317381c00001ffffefffe7fffff9830031f06ffff83887661c1f0008008f021900800031fc180c00007fffffffffffffffc8000001fffee20000c01f7e7fe00033ff
B3[194] <= 640'hb002c7fcff83ffbefe000080200030e763c00003cffe6fffe7ffff71377173fceffffe1c83ee0d39420a309ebe5d0001807bff381e010007ff7fe7fffffffffdcc0001387ffc0000181ffffe00003b7f
B3[195] <= 640'h9000c7ffff81ff7ffc8000c0c00003cf76007003fffffffffffffff83e7973fecefee60007fe01306003789ffefd0001ce7fdfe10f980007bffffeff7ffffffffc0000307f4c8000009f7efc0001837f
B3[196] <= 640'hcce7ffff71fff43c0000008100061f7680c3e3f3ff3efffffffffc329f7ffffffee6801fff018060309c9ffffd00309e3fdee01fd8800399cf3c70397fd9feff00800033c400200007fe9fc001c4ff
B3[197] <= 640'ha08fffffffe027ec1f0000000000001ffec1c77ff3e77fffffffff9fb38ffffffbfee6c003ff88060036dffffdbe8030873fff8001c1c0019b8ef9e081ff993effc1f200000000000007ffce0080fcff
B3[198] <= 640'hf71bfffe87f200400f70006000000003fcffff7f73f7f9fffeff3fffb7f7fffffffef90003ff8c06001ffffffffe00008b3fff880367fc80011ce18080038106fffff600000080000007ffc800007fff
B3[199] <= 640'hfd7e9fff03fe20000f000c01000006035f1fffff33ff9ffffe6712ff3ef3ff7fffef9100137cf0200086ffffffef0001bc9f9f98037e3bfc003100c018018102ffffffc000200020061fff8e000172ff
B3[200] <= 640'hfe7c03e021ff0318077000000000003f967f73fff0f3ffff929863fcfb7cffffffff7e0c23df70010003ff7bfffb4007c4e7ffe20fff9f7e00000000000060023effffde20000000001fff018406ffff
B3[201] <= 640'hff000160007f923903e000000000003fdeffb3fef70fff3f9f9063feffffffffffffe30477ffe000003ffffbfffe6007efffff2607ffbfff00038000988000001fff7fff00004000000ffe000000fffc
B3[202] <= 640'hc1100000003ffeff03e1000000002007dc7e330ce0dedeffb30000ffffffffffcffee300ffffe002007fdbf37ffe8000ffff7ff803fffffff020000080000000023ffffff8004800003fff800000ffff
B3[203] <= 640'h37c00201fffff01e1000000093007f33cb080c0fefffff00000ffffffffffdffe6080fffffe060f7e81017ffe9000fb3ffffcc07ffee7c4e0604000000000007ffffffe0f7d00007ee7800100ffcf
B3[204] <= 640'hc3f800200fcd07c0f000000001303ff13cf000003f7ffff00000ffff7fffff7fff7680fefbfe661ffed8007dff8101f03eff9f801fffe0c7000e4080000180007f3ffffff8fdf0007fe700c00cffff
B3[205] <= 640'hfff8607003c00380b000041901783ffc3fe600007f7fffbe00000feffefffe7effe300fce1fefffffc98187c3fc15ff8fffff90006b7f403c480000000008000307fffffffff9330ecff00c00dff7f
B3[206] <= 640'hffffffffc0000180f800033ffffffffc3fe60000fffff77e0000040ffeffff7f9c0000fcc07fffff798080003ff6bffefffff800063b7e01e0c000001800840039fbfffeffbffb7bfef8006009ff77
B3[207] <= 640'h3ffcfffffff00201c07e8000bffffffffc3ce000008fcfff7e08000037ffffffff1c00001c0466fefee1810000767e3ffffffe99034619362004040001000006003f3fffffffbff9fff7d1806319ffff
B3[208] <= 640'hfff97ffffffc3ec1c4ff01007fff6fffff7c7027077eff7ff807a4839fef7ffffc00000042903df0ff000400007ffefffeffff400087ff998303c6008100f0c0800173fffffffbeffcfeffc089c07fff
B3[209] <= 640'hfff9ffffffff7fc0e40fe3007ffffffff83f8000833fe7fff82002001ffffffcff800000400013f97c000000001ffcffffffffe400ffff8d8be007000080c1100000737fffffffcffffffb081bfcefff
B3[210] <= 640'hfffffffffe3fe7c87c1fffc1ffffe33ffe7e0260013fcffffd8002001f73fffeff810000380003387800000c71037ffffbfffffe0070ffc63d06071800800300c000633ffffff7ffffeffc080ffcc7ff
B3[211] <= 640'hfffff3ffdc7ffffc3c03ffc3ffff00001cff060001ffffcfff8080007ff7ff7ffc000001980000383800043fffc03fff810007fe01005fe63900000000000081c000637fffffffffffffff869ffc7fff
B3[212] <= 640'hfffff3fc01fffff83c01ffffffff000038ff000009fffff0ff01c000ffffffe67c0000079800203800003f3fffe010fe000001fec0010f7073e000010000000007000063dffffeffffffef065ef17fff
B3[213] <= 640'hfffeefcc0107dbf83f017ffffffe000038ff40000dfffe307f0110007fb7ffe4070000039800003080003fffffff033c0000003fe8010f7941c00003e620180000000047ffffefffff7fe00bf3f1ffff
B3[214] <= 640'hff67fe8000049fff0f000b7fe018068000ff400069fffc0307f178007ff57e0f030000017e00010080001ffff3ff0008003ff801ff000c7944000003eee0180000000023fbffefffffffe80bb873efff
B3[215] <= 640'he0675e80081000ff87e7803cc0012686001f50026ffff80007dfff017fff7e98000000017e000800001c1fffc4fe000009fffe003ff1000004000623ffe081380000007039ce7effffbe8812d17b1fff
B3[216] <= 640'he4007f003c00809fc3ff80046001cff8007f41263bffec80007ffffbffffff86000000000f000000000ffff8839fe0001ffffffc0ff2000000001803e0e083300000000180efec7dbb89c1464df8ff0f
B3[217] <= 640'hfe803e001cc0000f807ff0000003fff8803f00363fff400000fffffffffffe07000000000f000000001f7fc00003f800ffe0fffe07fe800000008007ffffe70000000100003eed9ffff9802ab0eb7fe7
B3[218] <= 640'hfb817c031c00001ff03ff80108fffefc803e0c36ffff0000007fffffffff7e000000000007000007001fff800000ffffff0003ff80eff880000081dffffff7c400010300043ca38ffef9188fd3297b35
B3[219] <= 640'hf7d9c0019f00181ffc1bf9182effcffe80ff4ce7fffc830e003fffffffffff800000000003c0003f00ffff0000001ffffe00001ff04ffe07a00003fffffffffc0000008000836399fe7b0072f5887bbf
B3[220] <= 640'hfffffc00bff81803fe017fd806ffcfff007e6dfffffc830c011e0ffffffeff8000000000c3e0003e03fffe0000000ffe00000003fc0dff7fa0002eafbffffff800000000000161f1fb780065e1ef3fa3
B3[221] <= 640'h7e7c3c00fffc1820ffc06fdf47ff00ff001e6fefffb80180808c03b9dffffc0001000000e1c0003ffffffc000000000000000000fc017ffff8003ee78fff7fe300000008803c30e57ff08013c8ab0787
B3[222] <= 640'h4e188000ffff1c2003e007ffe7f9003f403f4fefff8002f8000100110eff3800010000002000003fffe7ff000042000000011000fc017fffff0067ffcfffffff00000000803c00857fe601809a68cf59
B3[223] <= 640'hc6800c84fffffc0001fc007fffff303f60ffcc7cff800ef900010000dc7e800030000000201803ffffc3ffc000e0000000007f003f31ffffff8047ffc7ffff3c0000008100030c180e07082959356f97
B3[224] <= 640'h890002b9ffff3800007f00007ffff1ff01fffff018003c00000000005c6f98003041000000c003ffffc1ffc0000120007e03ff803ff07ffbfe003ffffffff9e0000000000000114ed10590b00199046e
B3[225] <= 640'h980003fffffff000007fe00000fff1ff00ffffc00000ef8000000000083e98003000100007300fffff807fc000002000ff013f803ffc3ffffef007ffc7fffb0000000000000010de18e190ab88a22c61
B3[226] <= 640'h103bffffff0000007f80000e971ff00ffff000003fff000000000003c600000001c0060180f7ffe007fc000003100fc803fd81ffe0ffffe200081c37ffe00000000000000058a3d0124a1a8dbaf40
B3[227] <= 640'h6008ffffffff3180000fe8000c021fe01fffc00000ffffc000000000000600000001800e000060ffc003fc000007900ff801fd80ffe07fffff800c383ffff0000000000000004f93ef861794c5dd675
B3[228] <= 640'h21cbfffffffff600000fe80004700fe81fff0000078e7fc00000000000000000000000000000687fe00338000007000ff0003000ffe077ffff800c308fffe00000000000000041613a86bf7dec94001
B3[229] <= 640'h81e3fffffffffff88007e80001c14ff01ffe000007fffff00000000000000000000000000000fc7ff00018000007004ff0100000ffe07fbfffa02e33effff00000040000000052442f04ae581627471
B3[230] <= 640'h281e3ffffffffffffc001f88001c1dff007f0000003e3dff80000000000000000000000000001fffff0001c00000008fff0000001ffc07fffffc0aaa3efffff800000000000001403b780fd28d3a0ee1
B3[231] <= 640'h66cf3feffffffbfffe001f8e00183fff007e0008c17fc7ffe00400c0002066010000000000006f7cfc000000000001ffffc000001ffe07fffff8022a83fffff800003800000000ca79b8099ee68e6860
B3[232] <= 640'h2f3ffffffffffefffe001f80c00033ffe07c001980fb1fffc08400c0000000312000080000001fffffc000ffe000003fffe000003ffe03fffee8002007bffff80000000000200122f20acabe9b382953
B3[233] <= 640'hffffffffffffff1ffe000fc8600001fff0380003effc1ffffc0e080000033c310000000000001fe0fcc001ffe600003efff000003ffc03fffee8000103fffffc000000000080137442903ce043335fe4
B3[234] <= 640'hffffffffffffe3073c0005fffc80101ffc000003fffc3ffffe1e1f0000077e710000000000039f78fcf801fffe8000fce4c000001ffc03fffee00003a8fffffe0000028000813135b2b372e90021e8e4
B3[235] <= 640'hffffffffffffc11f200001fffe80000ffc000e87fffe1ffffff83f3f008eff7be00000000001fffffcf8000ffe8007fcfdc000001ffc03ffffe00003fcffffff0000c3800000bf0c0a3234933137e025
B3[236] <= 640'hffffffffffffffff000007ffff80001f7e001effceffffffffe13fffc080ffffff0001000003ffffffff001fffc10001ff0000003ff803fff18000013efffffc0000c7000a006bd16480a1248479ec3e
B3[237] <= 640'hfffffefffffffffc201007ffffc0000f7f003ffffffffffffffffffffffcffffff0033c01c07ffe1ffff000ffbf90001ff0000003ffc0ffff38000003ffffffe0001100000813b4a52eb6483190b9b78
B3[238] <= 640'hffffdcf93ffffcf0002007fffff00003ff403fdfffffffffffffffffffffffffff60ffc00883fff3ffffc31ffff90003fd0000003ffc0fffe100000007fffffc0000100000019648ae11e2889c41b129
B3[239] <= 640'hfffe80000fffff000001effffcf00003ff780f8f9effffffffeffffffaffffffffff7ffc83c37fffff7efffffdfd8007e00000017ffc0fffe100001083fffffc00000000000206c51a9b89a3083cd1f0
B3[240] <= 640'hfffe0000000f17000007fffff3fc0001ff710ecf73fffffffffff77ffefffffffffffffe76fec7ffffff703ffffff00c00000001fff00fffff00000000ffff0072005873d11c7a046b403e14a1a2d9fd
B3[241] <= 640'hc7fc00000000000000effffffbfe0001fff30f8e77ffffffffff8727ffffffffffffffff7fffeffffffe7bfffffffc0000000001ffe00fffffc000001effff0050000050446c88a1a675f4d7353d570a
B3[242] <= 640'h3fffffffffff0000ffff37c687ffffffffff0f07ffffff7ffffffffffffffffffffefffffffffc0000000001ff0003fffff000003ff9ff601d80014046177b73069724c04ab65f56
B3[243] <= 640'hc13ffffffffffff8007fff338e867fffffffff1803ffc18e03ffffffffffffffffffffffffffffff0000000001ff0003fff7fc00067fffffa00f9063c1420b41fc4c89784e5b089df2
B3[244] <= 640'hc01ffffffffffff8007fff73fe841fffffffff7801fe0004007ffffffffffebf3ffffffffffcffff0000000001ff0000ffefff00003fffff800990682013d047c718ed3e24144a75b4
B3[245] <= 640'h3c07ffffffaebea8003fffffff800bffffffc3f000f80000003ffffff1fffeff7effffff1ff81fffc000000023ff000000efffc007ffffff800cd45f4413c8a1422263164b0c3b7212
B3[246] <= 640'h3edffff83f86be00001fffffff0000ffff79c37800f00008001fe7ff4047ff8330fffffe8ef01ffffc000003ffffc00000fffff803ffffffff52d4565423c911b13c297c2b504ab8f6
B3[247] <= 640'h7fff7e02f821c0004ffffffff0000fec000810000e000000007e7fe0007ff83f01ffffe84411ffffc000003ffffc00000fcfffc77ffffffff56dc5c4da3f11ecccd39976ac6910f69
B3[248] <= 640'he0033001003c07fffbf81e03c00000ffffffffc01ff80000018000000000000ff3f00007ff318000fbffe007ffffff0000037fff80000ffffffffffffffffd5855a089a04f9dafaca93f22ac03e57d
B3[249] <= 640'hce3007800000fc0fff6038080000001fffffffff01fff000000100000000000007ffe00007ffe38000037fc057ffffff000000fbffc0000fffffffffffffffffebbcde4061e3ba3f9307cddc081ca4f8
B3[250] <= 640'hff3f7fe100007cfffea020000020001fffffffff07fb00ff800000000000000000ffc00003fffb8000003fe017ffffff000000f7ffc00003fffffff00407d59f2e6127b5c00ee5c828b0c0c078c80055
B3[251] <= 640'hfffffff0000000fffef830000020007fffffffffffe001fff000000380000000001f000000e7ff703ce87fe017ffffff00000007ffc00000fffff0000000000653328d67c8b2b4491a7260a022a0082c
B3[252] <= 640'hffffffff8000037fffff70000020007fffffffffff0003fff800003f80000000fe0000000080ffffffffff003fffffff00000003ffe00000ffffc00038000002e33fec962bd844a325e864cb4e71b677
B3[253] <= 640'hffffff7fec00003ffffef8000000007fffffffffdc0007fffc8000ffc0000007ff000000000007ffffffff00ffa87ffe00000000fff8300000ff00007c0000905deb7dfb2224f890d6207f36301d0238
B3[254] <= 640'hffffffff7ff000fffffc80000000007fff7fffff881307ffffc000ffe0000003ffc0000000003fffffffff80fff8fffc000000007ffff80000fe0bfffefeebb040789c0c6d9bfc590603a12700c494e6
B3[255] <= 640'hfef7fffffbfffffffffc00000000007ffe7fffffde010fffffc000fff000000bffe1008000003fffffdffffffffffff800ff28001ffff80000003ffffff8e7bc55b5c76288906d669bcf25309c7349b7
B3[256] <= 640'hfff07bffb803fffffff800800030005ffeffffffff00c1ffff6001fff80000ffffffff8fa8ea03fffffffffffffcfff0007f08801c7fc40000003ffffffc1980e4fc8c15ea4e8aaf9b0a8ca805c0fef3
B3[257] <= 640'h800373fc9919fffffffc800001f8000fffffffffffe07bfffe6003fff80000ffffffffffffff0003ffffc7ff7fffbff000ff08071fffe0000003fffffff8016b291cdb3ad00f6865018625b82321fc93
B3[258] <= 640'hc003317e81007fc7ffff800007ff00003fffff80fff03ffffee00ffffc00ffffffffffffffff00000057dfff3fff1ff001ff001ffff82400023fffffffe06088b3930888af17268247129e18c142c4c7
B3[259] <= 640'hc000793ff8803bc3fffffc061fffb00003ffe3007ff81fffffe01ffffe7fffffffffffffffff80000000ffff01fc27e107ff003ffe000ef0003bffffffe000245933ccbc7bf519c28410430b9518091b
B3[260] <= 640'hc000fffffc000083f03fffff03fffff8003f000003fc03ffffe0fffffffffffff3ffffffffffe8ffaffaf3f00000790107ff007fec013fff0001ffffffe0000130ba7b89d1036007840347511910c004
B3[261] <= 640'he0007ffffc010001f81cffff83ffffff0000000000dc03ffffd1ffffffffffffe7ffffffffffffffffff380000007ffb017f007fc4007fff0000ffffffff0620e623d15af481b60746b186510424f54c
B3[262] <= 640'hf800061fde03fce03ffffffff3ffffffff000000001c01ffffd97ffffffffffffffffff1ffffffffffff81001f27ffff007f001fff00010c0001ffffffffc41ffaeb828c99db21534136035f721f00bf
B3[263] <= 640'hf800047f9f8fffff1fffffffffff011fff3c0fff801fc0ffffd93fffffffffffff7ffff8ffe7fffffffff0007effffff803f0003ffc00000017bfffffffee16dbe3c99896e5f4437c1dec54017282236
B3[264] <= 640'hff8000ffffe1ffff87fffffffff800017fffffff700071fffffffffffffffffffffffffffffcfffffd7ff73f0ffffffe003f8000003fffffffff803fffffe910e115b91889fb1bb26946274c8226c11e
B3[265] <= 640'hffc000fffffc3fff81fffffffff800001ffffffffb00207ffffffffffffffffffffffffffff00700e00ffffffffffffe013fc00078000000ffff00007fffa0b3aeb83b045920f0024a100ce2680e610b
B3[266] <= 640'h3ff8c0ffffffc0c8003fffffe0000118001fffffffff007f7fffffffffffffe3ffffffffff0000000001ffffbefffffe401fc09bffff81fe000000003fffff589fdbc30ee18b6031c8e087800c81a1ea
B3[267] <= 640'h3fffff80fff80000001fffc00003000007ffffffff877e3fffffffffffffc07fffffffff0000000001ffff03fffffcf3fffc3ffffffffe00000000c17c21bd49825905bf8fc2b186887134e539be00
B3[268] <= 640'hf80fffff001ffff103001fff8000030c80007effffffffee3fffffffffffff801fffffffff007f800000ffff83fffffd73feffffffffffff0ff800000000b65a8857892eae95c488e16847567aa02135
B3[269] <= 640'hff801fff000ff1fffff8fff8000000ff800000ffffffffc43fffffffffffff000ffffffffe00ff800000ffffe7fffff9cffc1fffffffffffffffbf188000f396b8cb4f5480e29736e73a9a262b9d40f4
B3[270] <= 640'hffe003ff030e003fffffff30000003ffc0000000ffffff003fffffffffffff0003fffffffc00ffe000008003ff3ffff89fe0001fffffffffffffffff80002d69b7c5cfa534baf2a12c4411670a082508
B3[271] <= 640'hfff803ffff8e007bffffff00000007ffe30000007ffef9003ffffffffffffd0003fffffffc00f8f000000000fe3ffffe7f800003ffffffffffffffff000099d6805062e219e49a324b39aa33e0113044
B3[272] <= 640'hfff03ffffff8000cfffc0000000000fff8000000fffff0001fffffffffffffc01ffffffffff8f80000000000037c21fdf0000000fffffffffffffffffe80fd6f3ad7e4507b2abae15678861d584ed40c
B3[273] <= 640'hfff01fffff3800003c000000000300fff8c000007ffff0003fffffffffffffe03ffffffffff8f8000000000001ff9ff00000000000ffffffffffffffffc0a06ec7729e4ee44644da5e12e06fe5f30aa1
B3[274] <= 640'hfff80ffffe000000180000000000001fe08000001ffff806ffffffffffffffe078fffffffff8ff8000000000000f83f00000000000ffffffffffffffff70d8e36365951a0c1fb27707e0042cc7043056
B3[275] <= 640'hfff81ffff8380000000000000000001fe0e000000fff3f07fffffffffffcfffff8fffffffff8fc0000000000000011f00000000000ffffffffffffffff61bd19a60675dc78e59a38367576e4569202b8
B3[276] <= 640'hc700fffffff80000000000000000001fe0e0000003ff1ffffffffffffffefffffffffffffffef80000000000000039e000000000000fffffffff00ffff433db9b480f49d476f0800df2ea798d79907ee
B3[277] <= 640'h7fffffff00000000000000000001fe000000001fb1ffffffffffffffffffffffffffffffef00000000000000003c0000000000001ffffffff007fff43b4f5570404930542f90e67b3a2f9f049b7ce
B3[278] <= 640'h7fffffcc0700000000000000000000000000000000713fffffff7fffffffffffffffffffff7effe00000000000000100780000000000ffffffff00002f83a629a9ce49436338e90422cf2897bb8333a9
B3[279] <= 640'hfffffe000000000000000000000000000000000000201ffffc7f3fffffffffffffffffffff3fffe00000000000000000fc0000000000fffffffe000007dce89e519e110b5224a19ab260c044d04fac20
B3[280] <= 640'hfffffe000000000000000000000000000000000001c00fffff3e0cefffffffffffffffffffffffe0e000000000000001ff80000000e0ffffff0000008cd4ea48ea09604a499af029a49395418f0257c3
B3[281] <= 640'hf007fc0000000000000000000000000000000000010007ffff1e0effffffffffffffffffffffffe0c000000000005807ff8000000000ffffff0000008c4d28f1e28000015c25a865c101176f27a10a55
B3[282] <= 640'hfc0000000000000000000000000000000000000007fffc1f0fffffffffffffffffffffffffffffe00000e001f81fffc000000000ffffffff0000004a5bc1198e0800a81040b771a033c29bef060d
B3[283] <= 640'h3c8000000000000000000000000000000000000000fffc0f07fffffffffffffffffffffffffffce1c000f01ffefefff800000000fffffffe000000ec128a0fb2b1978b86551b36c5432dbbe2a904
B3[284] <= 640'h8000000000000000000000000000000000000000fff80e00fffffffffffffffffffffffffff8e1ffe0f89ffffcfffc7f00fffffffffff0000000e8698eda40f88ee8b36179c41d7650ac244179
B3[285] <= 640'hffff8e00fffffffffffffffffffffffffff0e1fff1f991fffffffcfffffffffffffff80000004b2045645344d00760454081243a51e13059bc
B3[286] <= 640'hffffffce0effffffffffffffffffffffffffe0e1fff9ffe03ffffffffffffffdfffffff8000000668a49daf224049fab1498b570e6c450e0e0f7
B3[287] <= 640'hffff3ffe1effffff1f3ffffffffffffffffff5f5fffdffe41ffffffffffffffffffffffc000000319ae1659520123a1b718e620186e93e061c6b
B3[288] <= 640'h737fff73033f8fffffffaafffffffffffffffffffffffff7fffffffffffffffffffffff0000080291b1089a3361c069a5dac70508e6598245faf
B3[289] <= 640'h717ffff807ffffffffff0fffffffffffffffffffffffff03fefffffffffffffffffffff8000000784344f2bfcb8c5b73a47f0166856a43366a08
B3[290] <= 640'h30007ffff7ffffffffff80001ffffffffffffffffffffffffffeffffffffffffffffffffffc0000001b323020870b04c0312095221991a685cb0745d
B3[291] <= 640'h78017bffe39fffffffff80003ffffffffffffffffffffffffffeff1faffeeabf00ffea800000000000a732c6102e8e44656fce4900b6425219b00d79
B3[292] <= 640'h7cffffffc1feffffffff80073ffffffffffffffffffffffffff0ff0f0000000000f0000000000000005bd3914dcd0f300a51c49fc24d00f99900214a
B3[293] <= 640'h7fffffffe3ffffffffffc0ff7ffffffffffffffffffffffffff1ff8000000000000000000000000023067290326f6c183a8b08da459c024538b010ec
B3[294] <= 640'h7fffffffe00fffffffffc03f8f7ffffffffffffffffffffffff3fff00000000000000007f00007ff7fa68092777be3194d4702fe44e37ed0635827b2
B3[295] <= 640'h1ffffffefc701fffffffc0ff007ffffffffffffffffffffffff1ffe0000070e000001fffffffffffff8cde03f19967c1bada74b183b986394641c861
B3[296] <= 640'h7fffffffe0030fffffff166677fffffffc1fffffffffffffffe1ffe000033ffe00007ffdbffffffffe71b0099b499e0440f85baac3738d7578a80e22
B3[297] <= 640'hffffffffa0230bffffffe26ffffffffffffffffffffffffffffffee00117ffffffffff7eb6b7fff0002b9f62f000019936086954019bac7f3179645c
B3[298] <= 640'h7fffffff80000aabffffb37fffffffffffffffffffffff38fffef8e0115fffffffffc060e2320000004f768618d4dea28e304413830d7cfefe2c9e66
B3[299] <= 640'h13ffffffe00010000ffff987fbfffffffffffffffffc000002020000077ffffbffffe001c220000000008859a1274e242fe83b822c7808d56c0996e50
B3[300] <= 640'h17fffff0000038000ffff90f3fffffffffffffffff000000000000000fffffa2bf8800407c24000c0105292bb2494a3c45371272706e6964c0c490715
B3[301] <= 640'h7fffff3eff730000ffffa271f73ffffffffffffff8000000001cf055ffffc00000001fc3c0085ff455238e321047000c5133bf18428a0f664039aa1c
B3[302] <= 640'hffffe30f80030000ffff76d9fbffffffffffffffe000000000f7ffffffff00000000ff48a40cffffffd49890017020ae022ac88e2181156920041924
B3[303] <= 640'hffffe30ba92300811ffff34f83d7fffffffffffff000000182c3fffffffe00000000ff90ae92ff7fffbba50eb93a0d4d1829dfe420cd4c306285596c
B3[304] <= 640'h500000000000000000000000000000007fffff007ffffff89ffe22c3b77bffffffffffffbf000006e1e61fffffff410200077bb02566827ffe6c4a7d81430f4bcb4c57828282e51f16842d1e
B3[305] <= 640'h780000000000000000000000000000007fffff00fffffffe1fe4fdcffc5cfffffffffffffc0003ff01ee039effff6fb0201cfa7cde8a6007fc2d9ba0c0152144e8224368313ee0f8caa2355a
B3[306] <= 640'h788000000000000000000000000000001fffffc1ffffffc03fe6d65fbc5a07ffffffffffff000006000007fffffdcfb2001c4e032ae86fc1ffc093120e76024908786ccd6027ac5d00f5a745
B3[307] <= 640'hf8e000000000000000000000000000001ffffff0ffffc30067d27d9111020018ffffffffffc0000000fe07fffcf0374fb8fc1f3ff4542ff13ffd986446068ad5d580ff3c7264ac80cf81ea37
B3[308] <= 640'h7e0000ffffcc000000000000000000000000000ffffff0fff780001c4619bc402f800100a3fffffcc000e00000030180fc070ffe781e9465797dfb7494dbc44153162181949eda9094f7c7a5f88a72
B3[309] <= 640'h7e0001fffecc000000000000000000000000001ffffff0fe000000595da9c00117f80400000100ffff01880000f8de80009d3ffe3f090d236eb9c3e0da113b2c80a03aa814dce1923d3be644d0940a
B3[310] <= 640'hfffff8fffff0cc0000000000000000007f000000fffffff0f00000005cd3db1a010cf862000016007fffff03ffff4ed37f00051f9ffff2c1e1b37ffe450c1b41850aa814b3f00515c17bc43100b80cb8
B3[311] <= 640'hfffff8ffffc0cc000000000000000000ff000001fffffff8600000007c40b17d0003e771001ffff847c77cf003e67001c1dfdc84a3fff8077cd4133035e1c75f114c0c60494acd50f0a1f2de642030e1
B3[312] <= 640'hffffffffffe7fffffcffff0000000000ffffe003ffffff0100000003f88f0090033e6c750018c0f90afd4bc0e39dc03ce707e9d67fddfc0d767b940031840b4507a26660ef2639817094337800745628
B3[313] <= 640'hffffffffffffff1f000000ffff040303000000ffc0fffff180003c00f872fcd7ffe25e747e8b07f8fd737540000601ff7f95f3697f7fbd611b253fffb2b56e98a9a600ca3dcce3428199a1b782603480
B3[314] <= 640'hffffffffff7effffffffff00d0f0fe00feffffc0ff00003ffe0007e0fc0c0c41f8bed39af974cf0040030f0785c907ffff3a47967ffdbe078a9f67ffe8d820c58e408083cc15ca6848f4c8ddda40904e
B3[315] <= 640'hfffffffffffffefff00f00ffffff00000000c1000cf00f007fff003e001de741e6ec01b7482a00809f7c07f7839d04ffe300bac93fb7f4b9cc60cff16ba5a587797101c0eca320a4c1d402a57a9c4465
B3[316] <= 640'hffffffffffc180000000000000030fff07ffffff00ffff00fffffff7ff381840000ee3676c4bc1268f8f821fff35fe1fe09783c93fbef300bbe4f5f17206c9a8117c29fe1faf099d21eab591e3728534
B3[317] <= 640'h3c00003fff7800000000000000ffffffffffc000ffe00000fc00ffff000407983002f0017c015b69a382e9ff7ffbfe1ffc0801001fa4ca8f848551fc4166f04089c24c22182404d50a51a38a27ce2cc1
B3[318] <= 640'h7f300000008fffff00000000003ffe003000000ffffffffc00f3cfc8000f8f81000100cbd1cd63b8e9a384f7ffffcff386103a09b0fafe3e9c30f7ef2266399d0a116e6828e303c932f1a9a22ca465a
B3[319] <= 640'hc13ef8007ffcc0000000ffffffff7ffffffffffffeffff03e005ffff800000df0c70491f80b1d6772881ec607ff3fffe80600005c3397c58e857cb7fa56b0d2b5443ca0211c6d4680917bc8da9c60d1a
B3[320] <= 640'h3ffffffffff07fffffffeffffffffffffffffffe70100e000073fc0180000cfffffc11fc300dfdfe23f001168e071ff0000401c8670eab89fa06c171c05ac22e6728a0bd0263ca800b62f082ed02851
B3[321] <= 640'hbcffe1c0ffff03fffffffeffffffffffffffffff81000000000f7ffe1f1f03ffffff80f870008c807f1f02ffdaf000010000f0644c6a68a2e22f66134c68115e82ba363bd94e690940da53edd264001c
B3[322] <= 640'hfff00000000e3fffffff0ffc00003f07ff00fee3000000000000fffc07ff07fffffe07007863ffff7f001fbf3fac00000001e05869901e4a9cb66002429ce8f7ea802823a51116698110d448d7025681
B3[323] <= 640'hffffffffff1f1fffff1f1ff8000003030000f800000000000000fffc01f803ffffff0c8073f7ffffe7c0ff7df912018f8000c1ec253fc980ecec8a8f966166a816986c5804454635910302e7a0066a60
B3[324] <= 640'hffffffff000f07ff8007fffe00000000000000000000000000ce3ff800e003ffffff1f00cf7fff030780fffdffc200f100c0fbd8c36d9a73634587bb9c20e029a14a303024c1100a014607e268281854
B3[325] <= 640'hffff0000000003ff0000fffc00000000000000000000000001ff7ffc0000007fffff0fc0df7cffffff8000fff1fe3ff8000fe1d9bffc9404c20e5731168b3a78eb369c5032d435600206838a60605095
B3[326] <= 640'hfffffc8000007fff0000000000000000000000000000000001fffffff800003fffff17e00e1f86fffee2000f017b8088ffe01956ab2c8a5c77f8176a7712ae4620193f405409cc720105a664ee1e3204
B3[327] <= 640'hf1ffffffffffff0000000000000000000000000000000000ffffffff00001fffffffff8c007981c7d80708f0ff8080feff9f04250c86192875ab1fe2464290b04137406ec92419d98cbc75772a2c8a
B3[328] <= 640'h19fffec000f00000001ffffffffffffffffffbe0abfafae3f8e00000c0ff003effbc00c001fbc002f1808600fffc7ecc383f9c899919b8815073128c54d50d5c70c52236021040b28cb495ac6bce1d8c
B3[329] <= 640'h31ffff00ffffe0001f1f0007ef000000fffff8000000008000fffffc1ff00f7fff060000ffc0007d0ff0007f5f7f807607808c86e8245a070e6a87566c261c3980320a0c316750f690285e2a18f43380
B3[330] <= 640'h63ff8007000000ffe002ffe0c1800000fc3000f4e03f00000000ff00007c00fff8709fe0007fffff070fff7f000c00fcc7800241cc0491e51defcf297829d14daa3d2610822060b8d87a508319b21647
B3[331] <= 640'hb1380000008000f800ffe107f01c7fffffff80e03ff0001ffff8000f3ffffeffffffc0003c8700bf8fc0f300fff01ff8b9fe18448d8451b63c9b3ef8e04a0a00c14d3d0c432701e068603303b0204f04
B3[332] <= 640'h823f19ff8000c0fff8008000fe000000000001ffffff7f3ffffc001fff0000e000000000e0fffcf00007c0018ecc0f803c7f505bbca51acb09790c0fe9516981e04124b1d5d2249950de71e558b06c0c
B3[333] <= 640'h980cfffffffffffff00000800100000000000003f8001cff01000001fffffffe0000f807ffff70000f3e81c3de0003007fd12a97021bb59aeb028a6e624d39821a181209303520f0219025e87e004d
B3[334] <= 640'h3c01c0000000e07f00003f000f3c0000000000ffc00000c0001f03fffcfff0ffff60c3e007ffffd0008701ffc0ff0781001f0a0aa0b38681c08a0c6d477c50813104e10860442eb581b26c73914a0618
B3[335] <= 640'h7f6400c00000003f00877fffc3c1000077ff0e0f0000c004007ffffffffefffffe01480003f7e078003f00800003000040ff868708d89258122ebf2f2c122387110f50846809fb4a4024e2b86b0c56e4
B3[336] <= 640'h13ff9b03ff00ffff9fffffffffff00000000000000000000003cffff8fffffffff8003c00130e1fdc09ffff67fffefff0fb5b7751a913b15802ce5981645c78a44af480a208edc9d8800e0f143262850
B3[337] <= 640'hd3c01e31ffffffffffffffffffffe0000000000000000000003cffff0fffffffffc01ff8f000007cf87fc0001fffffff9c7f399281c74ec29654e45bd7e1ed860841bc04658260d1282130ba3f101270
B3[338] <= 640'h30f81e7fffffffffffffffffffffe000000000000000003007ffffffffffffffffffffff8000c3ffe8000603fffff9f0fb79d3e09de7426005ee483a529f40666003b8d737380b10066f81d25c82a18
B3[339] <= 640'hc1c1f032fff7ffffffffffffffffff000000000000000007ffffffffffffffffdffffffffc08000f3dffff007effefff38ee4c9c923b0590a004e9568ab7938110468480138490aa586bdb8d00e42ae2
B3[340] <= 640'h8dfffee3fffdfffffffffffffffffffc60007fe0e000007fffffffffffffffff0000f0fffc0a6000100fff0037200f7e0b4ffa83650e4883834c0a8b9b0208e84512bb61826c13224c050249816c5418
B3[341] <= 640'h5000fd07fffffffffffffffffffffffffc01fffcf000001fffffffffffffffff8000607ffc039000011800f80f783ffee3fa388b608f989b92527f6f636269c565a4c9e4b2257481047db2df48441a6d
B3[342] <= 640'h86007e73fffffffffffffffffffffffffffffffffdffd7ffffffffffffffffff03c0ffffffff5000039fff33546fe0f09f7dc764217308c48854628871b9e7a1246818611100114cc05ee3cf5234185a
B3[343] <= 640'hd6006737ffffffffffffffffffffffffffffffffffffffffffffffffffffffffbff9ffffffff0000039fff7c6020b46c6bc5199cb6404c8d504341103f01a615a04291d018f041a4041018083621070d
B3[344] <= 640'h9dc0ff98ffff9ffffffffffffffffffffffffffffffffffffeefffffffffffffad1ffaf9f53f4a06231ff37ee7a720dea962baae7727961c0cc66197af4c08b604b180810dc00f00940e20153d0b0120
B3[345] <= 640'h6ff8fe07fefeffffffffffffffffffffffffffffffffffffffe7ffffff73dcff9ff45bf5ff59857ef6c5393300e6f8cb8003e65fd603a288c6ae54fdc30993048997a3c0980592100c039622fb9c7809
B3[346] <= 640'h80f0ff0fffffffffffffffffffffffffffffffffffffffff0f817fff3ce693e1a37705ffbfa4abf7fc3a198cfc01e3fff7d335290abc2a5275d0e2c44e0a4750308fe8409001a05c811100b118880626
B3[347] <= 640'h36c07effff8fdfffffffffffffffffffffffffffffffffff07817fffff6790cff841420ab70a03b96f9946b8008ccffff6fa63d332630b7a44993029f4c4fc8b90e0c82c867009f01008c65178223160
B3[348] <= 640'hb981fffc00377ffffff03fffffffffffffffffffffffffff8e787ff1074de00244a997eef71d4b089f8f7e181f6a00400ea4c9e1aaccd0a41124540e628a80474344020802010580088e75461162127
B3[349] <= 640'h4d001fe73c0007ff001001ffffffffffffffffffffffff80f0e7873afb937ef2e8a78084306082ef7636008f03fccdf24230559c101408201a24e5319403855de202a7fc421893b10d88b0206d040080
B3[350] <= 640'h9000f7f3f000fe8000001ff00ff1fffffffffff0000ff0080e70005f1f8077975d641b1e4fc5d7f5131003ff1ff5817bfbaa45c361f2246b3034ba04259532f4601aa4c010001102c86201117120828
B3[351] <= 640'h120007fdff3f9fc0000007f800e000a0001f1fff0000000003800006071f63cfd2d3c221c7abaeeef8b383fffffe0ff80c3d13ca105082841b04318c86c8859371422004008000a01001083308201370
B3[352] <= 640'hd00007cffff3fffe70033f8600100001807a0ff0f70000008000003df2fe6a688f49e096865aadf6093220ff7a64e7993fa13009020d10973840852ddc85024c043b52087182a40044119000d023d87
B3[353] <= 640'h400001fffff811fffc00ff8001000e4033f03ff800001c042801007fff87f7bb7b51a982f494fea22856bc3ff9e0dfe9e821bc8d18536c9d8db0358fb40ce1926229818041b900410824104560c54bc
B3[354] <= 640'h10c00007ffff80031b7f9fe00e1c30c37e060300000003f008007fffffffbf231e819d768594db07f1ada93f7e1703c781a21c06612af360dc13f076c1e48218f16ac0d80304c4cb50868a8246102603
B3[355] <= 640'h11c2000317ffc3c3fc49c01f838f0f3f04000000ec3f03fe700f7fff00803f740e4107e145aec5dbd0b80f07fe79ff0783d94044e302106322f361c63c00d8ae0340a7f2260290880a60b10444002322
B3[356] <= 640'h15cf80000009ffff8518cbf801ef67ff2b7007c70fff07f980c3800100009e424c21c2903480952892ead3fc04b00002024f8c644168ce94481481540d60c845270a0058a200d0040900100ac0892526
B3[357] <= 640'h29ff900000008fd006c7f5ffffe1f300a1fc3f4673ff0fffe1e00000000031434611510460b8ebe24caa3dff8031cfe042729766d444a36e72dad9d9012b80208106a0ce0620e8d463403406a01a222c
B3[358] <= 640'h69fb3800000000df007fba6fff430fff8700b0184fff1fff3e3e00004021794fa30a410a969b2d65749ed5cf3f282ff8e256828013636e1e299a43063f00433c2f07c4c846024602300020102e041cb1
B3[359] <= 640'h9f0180000000086fe0206616c87fffff8c37cfc1ff81f27787f0000e08611d223c0c13a9816e3a7860b5a0c0b63affffc49ca0624e10c8196f6bec2a41b4216811404230086261c888c033108102497
B3[360] <= 640'h7790c072000100077ffffe0000ffff1d7e1f7e0118611980380c0c042080fb92dfd78757b7a4a93593eb9df86d505a1ffd38429624d7213d9589045e103816a53057e06b0065e10088d02700e844298f
B3[361] <= 640'h691f12996100001f07fffffe07e1ffeffd80fc07ff601af800460e6021f8fc12b0a093932580a81c84223100ffc4f71702d2182e241cb1346180b511e8c3521a1112200e80001980043022843e440540
B3[362] <= 640'h9393c210e48c001f007f0fffff81ffb0aeff00037f3cec3b800f060101fc779948062534c99ea473b9a971afba36fb80812f1a40159cf642259111ab91e8a03a29009201822190182c2284c412205809
B3[363] <= 640'h3595739cc0000002000001fffe00ff48a97f0001841f0ee3180e002546e60ffc8c58b055d2927e6953179f1f3b913d70e08948a88018438c7a121864f929c373498801108a80e4c02020c415100c1288
B3[364] <= 640'hc6704c3c809c0000000007ff7f11ff6f75fe00830000de3f030140047c7f079507fd20e2a852a811c700fa093bcb4bf9986933d832a095bb7114ba1709a9c365888c10da40116d092120585b18224244
B3[365] <= 640'h3cd383953103000000000fff7fffffd024fc003c000031fee1c0c4719e43b0d6cd494e9f0a849237d7128911022a65898ca8414c230e16c132385526f00626cc001400260011e341c2c60c049462806f
B3[366] <= 640'h59924afffaf3800000003ffeffffffa0de800004803c601ee026419390358092a005496385021006a08eb670172161796e6a4265026615fc98e101b4504624902c800356800010005c64808680001241
B3[367] <= 640'h37c005f95d58000000003ffcfffffff061c00000019fbc00018363c5090218c346db4124b488062d083ac33e3cd21a95e2c003002165607acc2170cb4904451eb049010030852e8814e65a48830608e1
B3[368] <= 640'h7a8980f805a43a0073ff1f08647f32000031061fff030c354765faa3a85dbf1199f0584cdb861309bf6322b78c0315042d2d009b01c33ee4999cc8a091e04c200830402cc80401000002dc2881
B3[369] <= 640'ha37eacdd3b7f20607ffff8f539983000300068cffff210c62b1a0fcf00f04db2c1091ec81263480afec4f4d6cf3bed82c030413f021012415cc664200b4a40228800003123808000031821048
B3[370] <= 640'h6f3e22ce2b931c2ffffff87f7cc805c001e20077ffffeaa1eccf98f8407c39d4c4009c69bc5889e7fe5463b10d5c2cac852104982a0e5c2c829a66309809114aa50084510000418300b6301c0
B3[371] <= 640'h4184dc3e22738419fffffff8926be2e7f3c0004f7fff8d02b4f5764b40ce58d001c2b88400a20b907fac7af05b3aa01e6c2285a8289812452ce9001c41484484042088240053005a2099440084
B3[372] <= 640'h90abd6dea02c8160003019b46d79c1980ff0ffffff83804210422f9323179a4c1de076c8000c20abeb029445c1009b010920c3022094034995140510022080ae202842000710d030008b01086
B3[373] <= 640'h87b563d729fea0c000001a77cfaf3f8170080ffe83cf01c9a03ac810e38b8b7964e185d381068087e20704668199c8032640069d1022c3298a0443c006022451008f712480600240004660190
B3[374] <= 640'h72efaf5c2f191180059a0dfba0003e0c386f8f09e20548c44e550cddca116544489012495858870e40d77b3b9d06000013d412090a00c81c222140271d98011c1b50120a612200000210688
B3[375] <= 640'h3eb8d1f9a5411c6ffffd5b0cd40003cccf9c0fc1f1f81929aa5909e81653b4405b9c4a050d6d4610488f5fda841804800412d40d9a23226c2c428262060124325c81b3c34125c000e304248
B3[376] <= 640'h1d230ed9ff8df74dff5ab00057300000cee77f187f9406448daa273186cf30c018005834030005d9edb03c01903020e26109c1c6061ca98738448b40e0071c021c118201c201500033f03ca
B3[377] <= 640'hf441cfe4be31381663ca000383008003fc004047960d2e649c62965ef8a99b03c56508f4314592da44527a1968614104a908420810f8b520061005b402d0cc8005805e1c920c00070f23ed
B3[378] <= 640'h100201c4a7f7e393900000002810000f0e7f100567f3da0f532be086491728845c9879190ade319a219801602062590087ec1186238443205c81ac32ac4013006818e18ca040000004028
B3[379] <= 640'h5efe009619a416570a40000d0313e0004602303e2bb3902723049aaec09b238c4243108894affcc2a14c8393308839401048369c5e24018518713dca41e1e68018c84184c1800c0000c22
B3[380] <= 640'h1957ef18668c91f76b40000c0ffffd80c7effff672934ff726758401688cc678b4479255c4b47d2d017d20833b090000000e2c36420887a10060c8203504c000000200030800000810ea2
B3[381] <= 640'hf534ffd0ff1b69df48000189fff1001f2ffdcf8a66b124070d79014526c88e47a8698850467fa44810e00e43035a0c1840100934feee1a4e1c00c4204401000000200004000000818c2a
B3[382] <= 640'h59fff80be4f9827040043863f3eeff7fce0ef75386cd1baa362f920869f004886ccc53035f7e084109270a460a3a2396c085017c64841631ac6462446401c0e212400c69200e0e1002a
B3[383] <= 640'h28b3ff96c3af56eaa1f5a4a9fff87fbff061fbf852020049c1685c2dd0f220ca9e108202a1e09060400208068482c3eca0c0039149910089154a40e8092411f00100167820000800029
B3[384] <= 640'hb8ff3fe0805807009f021c7d978e07ffc102b2d8f1f2708cf81160882dc1132591419144063261020c7b80c000f83ffe3f01d0ec64b36040c004380000c00700000019800000000000
B3[385] <= 640'h1d0fe3fffc000f90ed69d4686a3807ff5ffe831184a23454519fc2a868e8c0422480d9cd1459300e220e000000fffffc3fb88c980d9126140247000000000000000009800000000000
B3[386] <= 640'h2af00e001cff7f07f1ccff66b5fff8ffedfdce052cf4eba210198535b853344264000033063e231a2200100001ffffff7ff8060b08258e1d8262030000000000000009800000000000
B3[387] <= 640'h71400007f003cfc163303c78553fc0fff880218b9c7e825d614073681648a231008c0ed802c000060a043cc081fffffffffc0041000008ca7480de0000000000000009000000000000
B3[388] <= 640'h3c90e000007f989c037f54f55e7b00fef727c8c19955188a00a11311ed2273a8818000a8000243028601ff0701833ffffe7dafa7ad020002350dfe0000000000000008000000000000
B3[389] <= 640'h380000000000f677f00f0cef1d8c89fff0fbff807fc3fd90216e41b325c8a90d2116c31634d00818818b63e0a0e2c03df8600801ffffe1c5e18bb778de37c7fff0000000000000000000000000000
B3[390] <= 640'h400000000080e3d8ff000f7967e71a0c60dc801dbf105b2fc99803bd32008714e66210e42001a0420848085ac9001effc000e03fffff9c06be73d8ff27b86fff0000000000000000020000000000
B3[391] <= 640'h12000000000007f338ff80600181f8000dd95a0380d7987f78257bca72c585cf063230a400001ac1a694c161040084bf80718f8feffffdd1c2cc95035642ba3fc0000000000000000020000000000
B3[392] <= 640'h9200000000000347c00e00c3b1e111243666a3eaf4402417fa4ff965fe7bb0140582d887000030d06c1004000001f1fe000860078fffff20f61857fb23eff9ff80000000000e10000000000000000
B3[393] <= 640'hc2000000000000212000021c0f0f0ffe03ec6a1300d86607fbbf981f7e75a0cf309cc402704e000080000a0fc413f818000c60078ffefb29cc1e47fb7ffff1ee00000000000380000000000000000
B3[394] <= 640'h6c0000000000001eb00857fe17fe0e7fbf3ccaff87b8ae63f43818c7fffc0a30a4cd4010606700000033bc070ffff800001c000782f83929c80a67fbffeff0e8000000000043c0000000000000000
B3[395] <= 640'h100000000000000ea63f800003ff5f801f000b91098863e1f039f93831faf059a400008e40f78000111cf80007fc2000003c00078028302818aaedbbfffff04000000000000080000000000000000
B3[396] <= 640'h3a7c3fbc7f008efef002fafce0999b80e0397f139cfd81ed08810300e60fff80087ffe1e001e00000083c000000083b6f9b98c987fef8f02800000000000000000000000000000
B3[397] <= 640'h70000000000001aa1010ffff167e67fe10749c11b01803035ff33fcded51e029247036007c0ffff7dfe1f071e00003f83c000000003f2f1998448e27f8f07e000000000001c0000000000000000
B3[398] <= 640'h8040000000000000073c00038c3ff03f87f83a56c8f0007c9bdfff04b8f25eb5cd3b7fce003c0734f010018870f8f81ff031c00000001f3efed8619f33fef87f00000000000180000000000000000
B3[399] <= 640'h80000000000000000018ef8080060fcfc1fc9fc888000000cc0940cdfcb1fa360b0d0db8f80038cfbffaa001b8f0fff80ff1e1c00000001c3e02f8f197ffeff87f80000000000010000000000000000
B3[400] <= 640'h1cc9e000000003fc0009fe7e3c0100dc9618e7a21b6cfe5c92fb00000100000000003f879fff0000000000000080dffaaedeb97ffefee7600000000001180000000000000000
B3[401] <= 640'h2e0fc7f00003807fff206ff308303f0fe38b360fc60c5148fff0000010000000080ff00fff80000000000000081ffe80cc0bf7fb7fcff000000000000180000000000000000
B3[402] <= 640'h1200efff83c0ffc07f801007807f0e06e70d3e1ff7f36340ffe0000000000000080ff00fff80000000000000001ffc844e0ffffb3fa3f000000000018000000000000000000
B3[403] <= 640'h1bf30000000000ef800fc00f2743c270470edf3ff71fb178ffc00000080000000807ffffff80000000000000071ffc04f20ffffbff31f300000000180000000000000000000
B3[404] <= 640'h61f81f000effff000f03fe797df66f00f8e6c7fce0e3879ffc00000000000000800000000000000000000000717fe06f20edbf89f21f7800000001c1000000000000000000
B3[405] <= 640'h7a47c30038000e7ff42600bddfbbcff1f875fbf88c0f37fffc00000000000000800000000000000000000000207fedffacedbc65fa1ff80000000080000000000000000000
B3[406] <= 640'hf2e3cf803003387fff8f0c187f83ff7f87df9f3fce526fffe0000200000000080000000000000000000000000ffb9f9aceff82ffc03fc0000000080000000000000000000
B3[407] <= 640'h145fdffc17f71f80001c078e9cffffffb693c63ff320efffe0000600000000000000000000000000000000004fe903924e7fc95fcc1fc0000000080000000000000000000
B3[408] <= 640'h5286f9fff900002f8e0100ac06797ffc07fe37ffe33ffff800000000000000000000000000000000000000001ff899e6cf9e25ccc7fc30000000c0000000000000000100
B3[409] <= 640'h370800003c387fe200ff803e9e30fff80e51e1ff673ffff800000000000000000000000000000000000000001fffd9a6ef9c9dcdfefc2000000000000000000000000000
B3[410] <= 640'hdf000003e0000f98e0000c047fcfff81fedcc642a03fff800000000000000000000000000000000000000001fffc57fef9d9229ffdcc100000000000000000000000000
B3[411] <= 640'h20f7e07103860000ecce030591afff00f8e29fc3c01fff800000000000000000000000000000000000000000ffd3c7fce8d98d8c7cc0000000000000000000000000000
B3[412] <= 640'h1c3f8fffc7f707ffc8e00c0ff1ff8f0082383c92c00fff800000000000000000000000000000000000000000ef9b87f86c56bfcc7c00000000000000000000000000000
B3[413] <= 640'h31e7fffff7e0070fdee00005b2f3f00004223c7b00fff8000000000000000000000000000000000000000080efec0fc7b7607c1c801000000000000000000000000000
B3[414] <= 640'h3fa03fe78017907000f0007f48fc700003e9102200fff8000000000000000000000000000000000000000000effc0fe392b1bc1c800000000000000000000000000000
B3[415] <= 640'he1224f9072000380407780fcdff2000004d80ea00ffff0000000000000000000000000000000000000000800f919fa187761dc7800000000000000000000000000000
B3[416] <= 640'he89ce141003e00008000380837a0000e3f23706ff37700008000000000000000000000000000000700060199110000871a062f000080000000000000000000000100
B3[417] <= 640'h670fe0007ff8ff0fc0ff6479c6000fc0c0801684ff0000800000000000000000000000000000000007003cfa0000ff80e3fa000000000000000000000000000100
B3[418] <= 640'h1f5effece3c1000000e0f8064786001fc1f36001763d000000000000000000000000000000000000000700383e0000fc7ffe00000000000000000000000000000100
B3[419] <= 640'h3c31f8001c1ff83800010066d702003ff07de202cb8100000000000000000000000000000000000000e340b95200003e27e000000000000000000000000000000000
B3[420] <= 640'h1e7e3dec3fc000000000064a12002fff819d56cc6800000000000000000000000000000000000001ce178fb3100000f878000000000000000000000000000000000
B3[421] <= 640'h4d18f0000001f0ffe0ff7f6d8067fff001d4594b000000000000000000000000000000000000003e913c3ef8000086043800000000000000000000000000000000
B3[422] <= 640'h2027ffff0001ff078000994dd067fff0208e8b2ec000000000000000000000000000000000001f3eb13e3ffe03c000003800000000000000000000000000000000
B3[423] <= 640'h72bc3fffffe0000000c0200a28ffffff0c14b9404000000000000000000000000000000000001f3e113fe5dfc3e01c810000000080000000000000000000000000
B3[424] <= 640'h1f1765c00001c0000000000f887fff8f640117b1b00000620000000000000000000000000000070e6fbccfbfd2690e800100000100000000000000000000000801
B3[425] <= 640'had7c000000001f07033f1875ffff0eff80e072ef00000600000000000000000000000000000f8fa1ff8fe7cff883000000000000000000000000000000000800
B3[426] <= 640'h1e407100c1017fc2000fffcec3fe8c0cf83a8aff00010600000000000000000000000000001f8fe1ff8ff4094d810000a00060c0000000000000000000000000
B3[427] <= 640'hd798feffff0c0c00000f0ff84668b11fe0614fc00010000000000000000000000000000001e8f397f8ffc73cd1c18002b8082c0000000000000000000000100
B3[428] <= 640'hc16013f3fff00000000ff789e00cc97658331fe00000000000000000000000000000000001c1ff5ffced6c23ddc7803f88382c0000000000000000000000000
B3[429] <= 640'h19a43f87000000cffffff33e0003fe1fd719fe1000000000003000000000000000000000c001ffcffc447eb3dc3fc07fe7ff400000000000000000000000000
B3[430] <= 640'h1e023ff18388000fffff07c00fdc37907934efbc0000000000003000000000000000000000c009fedff8f8dbefdc3fc0f0ffe1e00000000000000000000000000
B3[431] <= 640'h3e03521022030fffffc00800e80f311976d83f800000000000003000000000000000000001e808fbcdc1fb23bfd1cc03ffff88f00000000000000000000000800
B3[432] <= 640'hed76dff7fffff0000071970b39d98afffcc40edff00000000800c2008000000000000000087fc0083c07f6f878071ffc00000000000000000000000000000
B3[433] <= 640'h13586ffffbfc000037fff070672bcffffcc017d8f180000008000070000000000000000001d10000183f83cff8070ff800000000000000000000000000000
B3[434] <= 640'h9901fe00000001019ff3e37c02e87ffffc000032180000000000070000000000000000001970000003127f07c070f8000000000000000000000100000000
B3[435] <= 640'hf53fc0fffcc038c0bf718c761fc05fffbc3000630000000000000000180000000000000008f800000000b303c070e0000000000000000000000100000000
B3[436] <= 640'h3d7800c00308f7fcc0c6c7c9c6061fff3c32001c0000000000c000001800000000000000023c0000307e3c01e03800000000000000000000000100000000
B3[437] <= 640'h2580001f7fffff99261800000005dff3cf2000300000000074000000000000000000000093c000001260001e00c00000000000000000000000000000000
B3[438] <= 640'hda03e7813fe079797f000000007dffbef3ffe4000000000bc0000000000000000000001bb0000003ff0001e00c00000000000000000000000000000000
B3[439] <= 640'h39f7ff1f10f346780000000000fffebfab2188800000000400000000000000000000000230000000200000e00400020000000000000000000400000000
B3[440] <= 640'he787f013c3cfe000000000001ffffff428188000000000000000000000000000000000c1c00000c000000400202800000000000000000000400006000
B3[441] <= 640'h3ce07d92aa800000000000000fffffb02c70600000000000000000000000000000000071e00000000000080300200000000000000000000000000e000
B3[442] <= 640'he33efcd60000000000000000fffffb894064000000000000000000000000000000000600000000002000001880180000000000000000000000006000
B3[443] <= 640'hfdfd6000000000000003cc00fffffbeacf9d00000000000000000000000000000000000084000000018000e8a0000000000000000000000000000000
B3[444] <= 640'h3e0180000280000000008001fffffea01fb800000000000000000000000000000000000f040000000fe00f8cb0800000000000000000000000000000
B3[445] <= 640'hc00000ff00000000000061fffffe6dffe000000000000000000000000000000000001f00000000180005def2000000000000000000000000008000
B3[446] <= 640'h1c000000000000000000062fffffeb207000000080000000000000000000000000000000000000060000b877a000000000000000000000000000000
B3[447] <= 640'h60000063fffffe1800c000000800000000000000000000000001c00000000000eacd04a51a000000000000000000000000008000
B3[448] <= 640'h87800107179effe0178000000080038013b0000000000000e13c0931f000000ce68e0352f80000080004000000000210000006000
B3[449] <= 640'h401fec00307139eff8c0e000000000003003b900000102c0000601000a13000000e2058afcb380000000030000010000000000002001
B3[450] <= 640'h6de80018703f877c00000000000000000181c0004486f8000000008c07000e002212388bcd000ff00001c000000000000000000000
B3[451] <= 640'h81c00df00018701f037e000000000000000001e13800fb2fa90000000006c0000e00010fdcf6010003f80001c000180018801000000000
B3[452] <= 640'h1c200ee00018701f03fec000000000008000017e8395801a6c000001008300000000720f86b00000000000018000000000000000000000
B3[453] <= 640'h34fa00b000018701f83fec0400000000000000319a2d270663800000000cf040000000e833ff0000030000001c000030003000008000000
B3[454] <= 640'h29da800000018721f032000f800000000100003c8e3397f1f100000781d41a480070031001c8000007880000160188300ffe0ff7e000e00
B3[455] <= 640'hd7a01b000018721e0ca23030000000004800032140edeaa0c2f69eebddaaa20000000880000000007800037fffe7fe01c67effff041f00
B3[456] <= 640'h400000000000000000000f920000000087c9f9dfab6000008811b4bc92b93c1b73601c03f67598cf64e800200416009017cffef000001b8000180dff8fdfec70600
B3[457] <= 640'h3fdfc000000a07df283f6ea33061feb381a58d2001ffe8c1f2c4ea1c6ee378518000ffe160fec0003607fff00988000f87bfdfdfff10200
B3[458] <= 640'h2800000000000000000787fc000000677cc0c2cd941822ebeac0019c92000302603ee3ed447eeca8bd3ac1fffee91e00cd8861ffffc01e0000d83e7cfdff703300
B3[459] <= 640'h400000000000007800006be00300000f7c7540c1f757468c8000800687800330f801ffee03382cc063d903ce76edde00058060fffffe1e0038fc1b3df1f9f037c0
B3[460] <= 640'h1f800000000000d8f80000100000000d37c0681b4fc9c810000000660193001d77bdf3f15e3934e5569d348ce76cdfe6f7da182ffff7e1e00007e09bdf0f9f812c0
B3[461] <= 640'h3a000000000000f68c0000000000001947c1f803fe00100411000004000d000dc8c7cffe85c1e10e0ed01a6c7f2d2fe7ffd8403fffffe0c00001207c573fddc1f00
B3[462] <= 640'h61003c001ec000000000000ee8f80000200080004c7800000002760700000000000080002f137ecf4259e2087fbb24df67b35bee7e628e030000ff06000003808379fc5c1c60
B3[463] <= 640'hff8ffcff9e9000000000000860d00000011c8000c7c90100b003cd0a0c000000000020002b8ffe3002e8c22881a452f842811b697ee4ae03fffffe26781801c03ff97c7e0290
B3[464] <= 640'h180000000000000000df5e8efff13e00000000000049f100000000090000edca8dc1e30003fe00000000000000002e007d5dd3e1d7dac025cf6520074a2007422c79fffffcffec3feff93f0b0e8e13e0
B3[465] <= 640'h1f0400003c00020f03ff6391cc81f800000000000048ec00000c000900003bb7bf37e781000e000000000000000026f0f9d85c60394fff078e42a51a4a209f7e8b73fffe79ff7f1e42860a17007e13e0
B3[466] <= 640'haf0bffffffffa00ffc1f25123ebb700000000000004f3800000c00090000f9b6fc367401000000000000000000001e07fe27f000067a1faf6088558dac609f7a0b63ffcefcfc000e05c60e1142e71000
B3[467] <= 640'h1c08717ffff9ffe0187cb4701046000000000000004ff900004c000980009feeecb642c000e0000000000000000010000fc86000003e18beff534cfc93c27806ecfcf3fcff803fef43ff000797820000
B3[468] <= 640'he1fe3ff07fcddc010797154281c0000000000000000d800004c0009800082ceaa20b0ce000000000000000000000c073fc0f80000097277e0fe68b41b0f7c03e1ff0e0fbff03ee0fd73900783c01300
B3[469] <= 640'h78ffe7e03fec03fcffe12f8537a00000000000000008000004c0009800002ce34c2bf720000400000000000000017dffe20180180000bde10c17cde5b3fcf19c4fc40060f1d40879ef250f813000200
B3[470] <= 640'he87e00003410ce0780feff1c5d80000000000000000000000480009800002cfa6066af6000040000000000000001700f800003f3500077b1b2aa69f53792379a7f07ffd1e8719abf4130ff809f08e00
B3[471] <= 640'h24dfc000c2e0dd700fff82ed31b80000000000000008400000080009800002cd8907298b0000000000000000000014f90e40012615e0007dfd243e4d2365a37870fc7d783e033251ba3a6bc04ff69380
B3[472] <= 640'hb4b6c77966f840060ffdef2f5f000000000000000004000000200008800000abc21826a08c008020000000000000194e4751a007abfc0000f81c4df9c665b492895b97c961c4183fc9a99cb3a9978190
B3[473] <= 640'hf9403ffddb3300380efff97e6e0000000000000000000000002000088000001aaa0c29468f050030000000000000153eb720b085b560000003304a8b8005f3c0c63bdcfb23411ef8e76ac883bda0a386
B3[474] <= 640'h43bef8ce6d3380f0ffffe190ac0f000000000000000080000060000880000018a80f3ed1be0500f8000000000000131cbc86b981ef800000000032ee60a5fcff703fd869b6f618fcf4fe768deb180082
B3[475] <= 640'hecc007ff70c3e10fffff4517b0060000000000000000e0000020000880000033880fe5ba9e060108000000000000398dec9a0160780000000000078e1e87c1e384d36121c0741b31c39082c7f3820e7f
B3[476] <= 640'hc06ff7fbddcff2ffc7c8ce200000000000000000007f0000020000880000003b8000ed76f03058c00000000000005c61f8356ee000000000000007fdebec1394ab740a17ad1f0e5e031dee76d019dff
B3[477] <= 640'h6f00fc6c592cffffc07959460000000000000000000ff0000020000880001c0ca80068034503867a0000000000000c8660049920000000000000000109273812bf390f4cedabd3d9179ce3f280fe01de
B3[478] <= 640'h6cfff3b1eaa3ffff83f6d3a80500000000000000000ff0000020000e8000140808003b3e6a8347620000000000000fc000032780000000000000000000c7fc903a4504941fba0bc4560dd6b06a1f866b
B3[479] <= 640'h5ffc0174d052fff787ef3ce20fe0000000000000000ff000012c000e8000944199001b1ce58468a00000000000000ee000005200000000020000e000000fef99608f2c122ef6d11390e255685844826a
end
always @(posedge vga_clk) begin
G0[0] <= 640'h0
G0[1] <= 640'h0
G0[2] <= 640'h0
G0[3] <= 640'h0
G0[4] <= 640'h0
G0[5] <= 640'h0
G0[6] <= 640'h0
G0[7] <= 640'h0
G0[8] <= 640'h0
G0[9] <= 640'h0
G0[10] <= 640'h0
G0[11] <= 640'h0
G0[12] <= 640'h0
G0[13] <= 640'h0
G0[14] <= 640'h0
G0[15] <= 640'h0
G0[16] <= 640'h0
G0[17] <= 640'h0
G0[18] <= 640'h0
G0[19] <= 640'h0
G0[20] <= 640'h0
G0[21] <= 640'h0
G0[22] <= 640'h0
G0[23] <= 640'h0
G0[24] <= 640'h0
G0[25] <= 640'h0
G0[26] <= 640'h0
G0[27] <= 640'h0
G0[28] <= 640'h0
G0[29] <= 640'h0
G0[30] <= 640'h0
G0[31] <= 640'h0
G0[32] <= 640'h0
G0[33] <= 640'h0
G0[34] <= 640'h0
G0[35] <= 640'h0
G0[36] <= 640'h0
G0[37] <= 640'h0
G0[38] <= 640'h0
G0[39] <= 640'h0
G0[40] <= 640'h0
G0[41] <= 640'h0
G0[42] <= 640'h0
G0[43] <= 640'h0
G0[44] <= 640'h0
G0[45] <= 640'h0
G0[46] <= 640'h0
G0[47] <= 640'h0
G0[48] <= 640'h0
G0[49] <= 640'h0
G0[50] <= 640'h0
G0[51] <= 640'h0
G0[52] <= 640'h0
G0[53] <= 640'h0
G0[54] <= 640'h0
G0[55] <= 640'h0
G0[56] <= 640'h0
G0[57] <= 640'h0
G0[58] <= 640'h0
G0[59] <= 640'h0
G0[60] <= 640'h0
G0[61] <= 640'h0
G0[62] <= 640'h0
G0[63] <= 640'h0
G0[64] <= 640'h0
G0[65] <= 640'h0
G0[66] <= 640'h0
G0[67] <= 640'h0
G0[68] <= 640'h0
G0[69] <= 640'h0
G0[70] <= 640'h0
G0[71] <= 640'h0
G0[72] <= 640'h0
G0[73] <= 640'h0
G0[74] <= 640'h0
G0[75] <= 640'h0
G0[76] <= 640'h0
G0[77] <= 640'h0
G0[78] <= 640'h0
G0[79] <= 640'h0
G0[80] <= 640'h0
G0[81] <= 640'h0
G0[82] <= 640'h0
G0[83] <= 640'h0
G0[84] <= 640'h0
G0[85] <= 640'h0
G0[86] <= 640'h0
G0[87] <= 640'h0
G0[88] <= 640'h0
G0[89] <= 640'h0
G0[90] <= 640'h0
G0[91] <= 640'h0
G0[92] <= 640'h0
G0[93] <= 640'h0
G0[94] <= 640'h0
G0[95] <= 640'h0
G0[96] <= 640'h0
G0[97] <= 640'h0
G0[98] <= 640'h0
G0[99] <= 640'h0
G0[100] <= 640'h0
G0[101] <= 640'h0
G0[102] <= 640'h0
G0[103] <= 640'h0
G0[104] <= 640'h0
G0[105] <= 640'h0
G0[106] <= 640'h0
G0[107] <= 640'h0
G0[108] <= 640'h0
G0[109] <= 640'h0
G0[110] <= 640'h0
G0[111] <= 640'h0
G0[112] <= 640'h0
G0[113] <= 640'h0
G0[114] <= 640'h0
G0[115] <= 640'h0
G0[116] <= 640'h0
G0[117] <= 640'h0
G0[118] <= 640'h0
G0[119] <= 640'h0
G0[120] <= 640'h800000000000000000000000000000000000000000000000000000000000000000000000000000
G0[121] <= 640'h0
G0[122] <= 640'h180000000000000000000000000000000000000000000000000000000000000000000000000000
G0[123] <= 640'h0
G0[124] <= 640'h0
G0[125] <= 640'h382000001c0000000000000000000000000000000000000000000000000000000000000000000000000000
G0[126] <= 640'h11fee000000c0000000000000000000000000000000000000000000000000000000000000000000000000000
G0[127] <= 640'h11ffe00000800000000000000000000000000000000000000000000000000000000000000000000000000000
G0[128] <= 640'h133ffc00000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[129] <= 640'hffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[130] <= 640'h8ffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[131] <= 640'h8ffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[132] <= 640'h8133fff80000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[133] <= 640'h28033ffe80000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[134] <= 640'h2001fffe00000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[135] <= 640'heffe00000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[136] <= 640'h7ff800000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[137] <= 640'h773800000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[138] <= 640'h373000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[139] <= 640'h166000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[140] <= 640'h164000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[141] <= 640'h8c000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[142] <= 640'h88000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[143] <= 640'h0
G0[144] <= 640'h0
G0[145] <= 640'h0
G0[146] <= 640'h0
G0[147] <= 640'h0
G0[148] <= 640'h0
G0[149] <= 640'h0
G0[150] <= 640'h0
G0[151] <= 640'h0
G0[152] <= 640'h0
G0[153] <= 640'h0
G0[154] <= 640'h0
G0[155] <= 640'h0
G0[156] <= 640'h0
G0[157] <= 640'h0
G0[158] <= 640'h0
G0[159] <= 640'h0
G0[160] <= 640'h0
G0[161] <= 640'h0
G0[162] <= 640'h0
G0[163] <= 640'h0
G0[164] <= 640'h0
G0[165] <= 640'h0
G0[166] <= 640'h0
G0[167] <= 640'h0
G0[168] <= 640'h0
G0[169] <= 640'h0
G0[170] <= 640'h0
G0[171] <= 640'h0
G0[172] <= 640'h0
G0[173] <= 640'h0
G0[174] <= 640'h0
G0[175] <= 640'h0
G0[176] <= 640'h0
G0[177] <= 640'h0
G0[178] <= 640'h0
G0[179] <= 640'h0
G0[180] <= 640'h0
G0[181] <= 640'h0
G0[182] <= 640'h0
G0[183] <= 640'h0
G0[184] <= 640'h0
G0[185] <= 640'h0
G0[186] <= 640'h0
G0[187] <= 640'h0
G0[188] <= 640'h0
G0[189] <= 640'h0
G0[190] <= 640'h0
G0[191] <= 640'h0
G0[192] <= 640'h0
G0[193] <= 640'h0
G0[194] <= 640'h0
G0[195] <= 640'h0
G0[196] <= 640'h0
G0[197] <= 640'h0
G0[198] <= 640'h0
G0[199] <= 640'h0
G0[200] <= 640'h0
G0[201] <= 640'h0
G0[202] <= 640'h0
G0[203] <= 640'h0
G0[204] <= 640'h0
G0[205] <= 640'h0
G0[206] <= 640'h4802000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[207] <= 640'h3d97600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[208] <= 640'h698fffb000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[209] <= 640'h689ffffe00600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[210] <= 640'h1ffffff1030000000000000000000000000000000000000000000000000000000000000000000000cefc7f0000000000000000000000000000000000000000000000000000000000000000000000
G0[211] <= 640'h803fffffff47c000000000000000000000000000000000000000000000000000000000000000000001ff7ffff000000000000000000000000000000000000000000000000000000000000000000000
G0[212] <= 640'h811fffffffffe000000000000000000000000000000000000000000000000000000000000000000001fffffffe00001c3ff00000000000000000000000000000000000000000000000000000000000
G0[213] <= 640'h187fffffffff0000000000000000000000000000000000000000000000000000000000000000000007fffffff00001ffffc0000000000000000000000000000000000000000000000000000000000
G0[214] <= 640'h143fffffffff80000000000000000000000000000000000000000000000000000000000000000001effffffff00019fffffe000000000000000000000000000000000000000000000000000000000
G0[215] <= 640'h77ffffffffff8000000000000000000000000000000000000000000000000000000000000000003fffffffff0001ffffffff80000000000000000000000000000000000000000000000000000000
G0[216] <= 640'h3ffffffffffe800000000000000000000000000000000000000000000000000000000000000001fffffffffff0ffffffffffe0000000000000000000000000000000000000000000000000000000
G0[217] <= 640'h2c001fffffffffff000000000000000000000000000000000000000000000000000000000000000f07fffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000
G0[218] <= 640'h7f817ffffffffffff00000000000000000000000000000000000000000000000000000000001c73fffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000
G0[219] <= 640'hffd9fffffffffffff80000000000000000000000000000000000000000000000000000000000cfffffffffffffffffffffffffffffb00000000000000000000000000000000000000000000000000000
G0[220] <= 640'hfffffffffffffffffe0000000000000000000000000000000000000000000000000000000000dffffffffffffffffffffffffffffff20000000000000000000000000000000000000000000000000000
G0[221] <= 640'hffffffffffffffffffc000000000000000000000000000000000000000000000000000000000fffffffffffffffffffffffffffffffe8000000000000000000000000000000000000000000000000000
G0[222] <= 640'hfffffffffffffffffff000000000000000000000000000000000000000000000000000000001fffffffffffffffffffffffffffffffe8000000000000000000000000000000000000000000000000000
G0[223] <= 640'hffffffffffffffffffff00000000008000000000000000000000000000000000000006000001fffffffffffffffffffffffffffffffe0000000000000000000000000000000000000000000000000000
G0[224] <= 640'hfffffffffffffffffffffc0000000c00000000000000000000000000000000003060f3000004ffffffffffffffffffffffffffffffffc000000000000000000000000000000000000000000000000000
G0[225] <= 640'hffffffffffffffffffffff0000000e000000000000000000000000000000000030003e0000037fffffffffffffffffffffffffffffffe000000000000000000000000000000000000000000000000000
G0[226] <= 640'hffffffffffffffffffffffc300008e000000000000000000000000000000000030003ec00083fffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000
G0[227] <= 640'hffffffffffffffffffffffe7e300ff000000000000013c38000000000000000030183cc100c3fffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000
G0[228] <= 640'hffffffffffffffffffffffffff07ff000000000000007efc000000000000000011187cc1003ffffffffffffffffffffffffffffffffffc00000000000000000000000000000000000000000000000000
G0[229] <= 640'hffffffffffffffffffffffffffdfff00000000000011fffe00000000000000002380f7e3003ffffffffffffffffffffffffffffffffffc00000000000000000000000000000000000000000000000000
G0[230] <= 640'hffffffffffffffffffffffffffffffc000000000001ffffff10c0000006046070340fff7c01ffffffffffffffffffffffffffffffffffc00000000000000000000000000000000000000000000000000
G0[231] <= 640'hffffffffffffffffffffffffffffffe000000000003fffffffde03ff007ce6ff6366fffef887fffffffffffffffffffffffffffffffffc00000000000000000000000000000000000000000000000000
G0[232] <= 640'hfffffffffffffffffffffffffffffff80000000000ffffffffdffeff47fffffff9c7feff7ffffffffffffffffffffffffffffffffffffe00000000000000000000000000000000000000000000000000
G0[233] <= 640'hfffffffffffffffffffffffffffffff800000003c7fffffffffffffffffffffff943fffffffffffffffffffffffffffffffffffffffffe00000000000000000000000000000000202000000000000000
G0[234] <= 640'hfffffffffffffffffffffffffffffffe00000003ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000000000000000000000000000040000000801000000
G0[235] <= 640'hffffffffffffffffffffffffffffffff80000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000000000000000000000000000808010000000000000
G0[236] <= 640'hffffffffffffffffffffffffffffffffc00000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff84000000000000f8c000000000000000448000000000000000
G0[237] <= 640'hffffffffffffffffffffffffffffffffc00000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0400000000001ffcc000000000000000004200000000000000
G0[238] <= 640'hffffffffffffffffffffffffffffffffe00007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000001fffff000000000000000020040000000008000
G0[239] <= 640'hfffffffffffffffffffffffffffffffff00007dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000001fffffc00000000000000420040000000000000
G0[240] <= 640'hfffffffffffffffffffffffffffffffffe200fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff078000000004ffff7c50000000000000026000000000000000
G0[241] <= 640'hffffffffffffffffffffffffffffffffff710fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000001ffffffe50000000000020004008000000000000
G0[242] <= 640'hffffffffffffffffffffffffffffffffffff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000ffffffffd0000000000090100000000000201200
G0[243] <= 640'hffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000fffffffffe8000000000000000411000400000000
G0[244] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe78fffffffffa8000000000000200000002000000000
G0[245] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc100000000041130004001000040200
G0[246] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc901000000062110004000000000000
G0[247] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc900090000201180010000000000020
G0[248] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd451409000028008000100b120000000
G0[249] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffea920011000804600000001980040800
G0[250] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4cb00008208480101010000080540800
G0[251] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec431443a202000080020000040400000
G0[252] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee4d24421002000c00000000000010000
G0[253] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe90920420010000001001000c00200000
G0[254] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec2640482002000101002094602400000
G0[255] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa4244008001001001844000106440840
G0[256] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa60681088008801001008021090440800
G0[257] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb60481849400001081102000400010000
G0[258] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd30104410001200001006004002000000
G0[259] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe9810b400100800019040060200101300
G0[260] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe56015209108000608982440010040000
G0[261] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff76222d108491180018910490240088400
G0[262] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb1b3cf630c99090988001078808204008
G0[263] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddcf26c204d98208284008040009002100
G0[264] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedc7414db259bc188104090102001000000
G0[265] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefb9e4cd8b752e0c801219010d200024000
G0[266] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedbdf44e1b0d2c2c6a183b01251c0100030
G0[267] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffeb2568b4e6643219c320320ce0000600
G0[268] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe77e7717891ec1b22484300380610090400
G0[269] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef7f77f340dcd9bf444e020094210193810
G0[270] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7bdbb12418dcb8b206a0280d4000104008
G0[271] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4dfb9738d3887c1b634ba0319840424200
G0[272] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecf1f298d2d225b90061921930181a4230
G0[273] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff76fdb4f419b280c58863a2866808041308
G0[274] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb37f4b1c40b225466a72164866400199906
G0[275] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff336e25849a2c64301992182c2904108900
G0[276] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff73b7f8ce8191863fe1d8202413000928920
G0[277] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbd7ecce00b30c8331e40f0033170c23108
G0[278] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddfb3c46e4813925f11f63fa0c9a7045380c
G0[279] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebe3948c2033a76fccba3e2649609412000
G0[280] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff6a7ec604364d26cce4661a705cb432000
G0[281] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff79817cd20c8359c34c765d109c93b870e01
G0[282] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3df67e58c012925fa7371c48164f8c24808
G0[283] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcdf8ce3842d6fc37f13604e658598404400
G0[284] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee6cf22648967e2ff8167ce64d389a05620
G0[285] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef8c27783148093b7fe6ca4e42449b9e25184
G0[286] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefe6d9fe31c8d35f9bf24f685258932606900
G0[287] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7f359bc2460c6764bfba6693830016001030
G0[288] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffde9de3c6ccef4effbc272b9c7070000070
G0[289] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff77fc3de69f28cce0f4fde226c84a8c1f06400
G0[290] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbbffb9e6998489e9727da048e844a64310708
G0[291] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcdfbd9d8b6c48db73afce011c10426e11006c
G0[292] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe74c4cf81a4489f66dfe080bfa36796c03224
G0[293] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff686024cde0413caf0fddc365934397707258
G0[294] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa6b0f75c1f3017d9be7cb070f4bcf8b50c242
G0[295] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff33cb36110219e1cdf7ebc61e1bd3614818c0
G0[296] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb10f9b2813e0887e1fbedc3f839f723783868
G0[297] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9a389800c1994eece9e583f2dcee67187b2c
G0[298] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee5d051189093906ecce483d9fcdedad8f914
G0[299] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb0d60dac06033ff6e6778331f67d88c89900
G0[300] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecf038202c0c56e52fb3060e6ce393ce849a0
G0[301] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff12cf408c08cd93aef92210462007e78e190
G0[302] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffffffff18c4b3647189ce1cebcc20689b00f9383724
G0[303] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3ffffffffffffffffffffffffffffffffffffffffffffffff1fffffffffffbe614199415a80cc463e061d9cf12b598b26c
G0[304] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1ff87ffffffffffffffffffffffffffffffffffffffffffff5fffffffffffff62e08140220b9ee2ff2639ee3338bd83858
G0[305] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc01f807fffffffffffffffffffffffffffffffffffffffffffb1fffffffffff3c42131c92363b34e0cb9e13ff8952fe85842
G0[306] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe007f807ffffffffffffffffffffffffffffffffffffffffffff17ffbfffffec9f0991080206673d90e38617de885e7e4f84a
G0[307] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc01ff003fffffffffffffffffffffffffffffffffffffffffff921fa1ffffff6ff8416e04b040f69bfb6c20fbcf846ff0d884
G0[308] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff003f0003fffffffffffffffffffffffffffffffffffffffffff90dff7ffffff6ffbb087319861221d8f6d20f73f8e66f8c803
G0[309] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc03f00001fffffffffffffffffffffffffffffffffffffffffff98fff3ffffffb9ffb21c2d4a238cfd967d8189ff8f8dfc6061
G0[310] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbbf0c000fffffffffffffffffffffffffffffffffffffffffff9dffdbffffffffdf595c94e64333fbd93981f3fbb599fc2031
G0[311] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff90300007fffffffffffffffffffffffffffffffffe3fffffffb5ffffffffffdfff0ecdcc466267f39f1681ceff7218fc9830
G0[312] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff06e00007fffffffffffffffffffffffffffffffffc1fffffffb9bffbffffffb3e7ee4a6602e62ff697e4c19ffe5222fcc810
G0[313] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000e007ffffffffffffffffffffffffffff003fffffffdcfff3fffffcbbfb5da0c330e327bfdf32c0ffdcdb8f7ce0c6
G0[314] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe03000000c01ffffffffffffffffffffffffffff8007fffffffe9fff3fffffc9bf9f6d059b9e36f299b38e1ffd9ed2fbc80c6
G0[315] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe1fc03eff000fffdffffffffffffffffffffffff8fffffffffffdff7bffffffbdfff2637c89e18de79efceb6ef3ec33bcc244
G0[316] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff81c1e0007fffffffffffffffffffffffffffffffffffffff5ff3bffffff9cffda30dc48a0c9c718f9491df7a83cfe6220
G0[317] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcfff0003fe81fffbfffffffffffffffffffffffffffffffdfff3ffffff5efbfd30e7644201923df909d84fe67edc4040
G0[318] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80017c007f80fffc0ffffffffffffffffffffffffffdfbf2fffff70cf79e88e3b06081601bfea96edfaf3fcc4040
G0[319] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0007c000f007ff001ffffffffffffffffffffffffe4dbf7fffff76736ffd6239a08dbc093f6c16510613fc40600
G0[320] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc001800000000c0001fffffffffffffffffffffffe49d3777fffda33bbd0611c208db3423f641730d859ff81232
G0[321] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff07c000000000000000fffffffffffffffffffffff6f472d3fffe8e93e59e4cb02199fe08e7017a5eb19fec3099
G0[322] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7c600000000000000007ffffffffffffffffbffbaeeecf3fffe01ca63cd00d861000631db8138fffcce8c6049
G0[323] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000001ffffffffffff7feef5fba5ee7b3fffc20024874186c400c06323281333f45ce3416e0
G0[324] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000000000007ffffffffff97feffff9a94677bfff623901f111a1e6c0e76232e89677d6124d84830
G0[325] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc0000000000000000ffffffffff939c86b7cc4e669bfffe23994ffc3b88248c3e3674414b73cd07c47026
G0[326] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb1000000000000001fffffffff93b4c23bfe6ccd89fffe3375ef2e14c864c0371420c119fcd987043666
G0[327] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000007fffffff83f6891ff74c9b33dff7b32c11e58c663444124cd809125c9172fe46ec
G0[328] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000000000003fffffffff53ff9d9fbf3c1a7bdfdce1c968a1800312221262d209265fb919f85808
G0[329] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8fc000000000039fffffffdfdb199fdd3c4efbd6fceb5b9fc1b09c1a32276663c02d2f92f9d828c0
G0[330] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff001ffff3f03cfffffffcffb0edfe62451efd7fc43f3ccd0191e08120b156848697801606862d9
G0[331] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0bf60b6ff638df9b9ffe4db2674901db00810605cc4878386190e4569b
G0[332] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe43ef0b0bfb2d9799bffe5b66f1c0c4619299e2269dc83c3e7148d86625
G0[333] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe13ff0f9bfd3b8f993bdb235bc8d8ce11904c32363c01b136737a74640b
G0[334] <= 640'h1efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe8fed1707fe349b297779275d1a2c0fc3000c24213c80d36ef9fb266e32
G0[335] <= 640'h83fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec5e94b87bf3d36da55e85a679d9987f10c0620c07d884b3e71f90c6835
G0[336] <= 640'h447ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc27e2db4ff9393c4ce6b0686084e0e73c8c200244b988473eb9fb367876
G0[337] <= 640'h4400ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff27f8cd25cbab7a65ffb02949ac4027760620402cb188273ecbf2560a5a
G0[338] <= 640'hff803fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffabe485a58fb23cedb79039c4966001a303106204510837bce5bcc61a59
G0[339] <= 640'h4c3f80fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe83e408a3c6923c5d87941238cc3801874311082048487bfdf1d9c83263
G0[340] <= 640'h10013fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe42edaf4bd799797dcfda112a4488b1b1c0130c608048392471e4ee223c
G0[341] <= 640'hcc0017ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbc4827199b9a633dcb6a324c12683038021900108c443ca551e4a6283c
G0[342] <= 640'h79019fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefc9317f0df19a675dcff278cc0320503402180011ccc63e9bd1ce321c0c
G0[343] <= 640'he009ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed881205b0cfd9a6fcd04f04841340033898188820134823c08f19e321a4e
G0[344] <= 640'h2001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffff900026f0e30cfd4e4eed9ffc0811b20038c30080800120c61d307028103270
G0[345] <= 640'h1000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffff00fe003fff900024d0f937fc8c4dfd95d9310c8c9e81c1c9180010069615907030180829
G0[346] <= 640'h1000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9ffffffffe00007e000000300102509d1b2e8c9ded8cec1b218c20415c60882018100606083193080022
G0[347] <= 640'h11c9fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdff9c6ffff00001f000000000001233c195f855bb529ec596491f0000600c46010300010084070200904
G0[348] <= 640'h13cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8ffffff98d800000ff3e0007c00010060200001e7dc6c07b7533f2785e1ffee280200c0010301018000400261921
G0[349] <= 640'h101c067ffffffffffffffffffffffffffffffffffffffffffffffffff8c61ffff8b80fcfff80000000000000003fff9bffc00160002264e4037f773d87c3f0bb26b74b04c0800100008900001300029
G0[350] <= 640'h60000033f7ffffffffffffffffffffffffffffffffffffffffffffffe000007e393821f7ff000000000000000007ffffffe000a0000072141677273f871ea2ce70c3618020800800000000060341129
G0[351] <= 640'hc000023fc7fffffffffffffffffffffffffffffffffffffffffffffffc0000040900401f9f0020000000000000067fffffe0080100813216297f8d9f4b9ec24224611c4000000c0200000000004112b
G0[352] <= 640'h50000033ffffffffffffffffffffffffffffffffffffffffffffffffffe000200203462a9f006bf2000000000007ffffffc00808024119100b7983d7cb96873c9213340000121602001000480200900
G0[353] <= 640'hc0000003ffffffffffffffffffffffffffffffffffffffffffffffffffff980000028ffbff827ffe401bf8000063ffffffd000010291e11c8b7d0fefc69f26de0019818000005004680000026080900
G0[354] <= 640'hc00001000fffffffffffffffffffffffffffffffffffffffffffffffffffff1734c93f67f784fffe409fffffc9fffffffff0ca5120953630093d87e74c9e4bc2008cca00000008c2000000206000000
G0[355] <= 640'hc0000000000c7fcbffffffffffffffffffffffffffffffffffffffffffffffb6388b6ee7d184feff57fffffffffffffffff40a523209b2388bbe53d1c7be84e6309e1200100002c1200000044000100
G0[356] <= 640'hc000000000033fffbffffffffffff803fffffffffffffffffffffffffffffff7388258cfd9a4ffffd3ffffffff9ffffffffec4ca4facc94f05de5e78c71d12023121180000008080000000480b00024
G0[357] <= 640'hc000000000031ffffffffffffffc780c3fffffffffffffffffffffffffffffcb1880b8cfb127e3ff937fffffff9fffffffeff76e6564612f0ffd8cfcc69800001030000000000042200000040900200
G0[358] <= 640'hc00000000003003ff7ffffffffcffff91ffe001fffffffffffffffffffffffdc1812b8cfe196e7fe97bffffffffffffffffbf26c6c02a71219edcdf615b644a02000000000004000300200002400800
G0[359] <= 640'hc00000000000001040019bffe6650001f07fe003ffffffffffffffffffffffdb3806b096c0c6ffff05bffffffffffffffffff94cde48cb9b2ff3cdfd03ac03302000000000000009000000000000000
G0[360] <= 640'hc07e00000000000001c0000e08000a040000000ffffffffffffffffffff83fcc1841f1dae02afbff43bfffffff7fffffffffeda65c4e498f2df3c8fd879840420040000000000009000000000000000
G0[361] <= 640'hd3d3c48000000000000001d0000000fc0000007ffffffffffffffffffe70ffee4841b9dc8003e3ff27f7ffffff7ffffffffbe6e6599f364e3963c8be879020020000000000000008000000000000800
G0[362] <= 640'h8e00e10e00000000000000000000010a000000fef817fffffffffffff818ffd53027319dc042e3fe337fffffff7ffffffffffe02710e376b2ddbc8fe930403080000000000000080400000000400000
G0[363] <= 640'hec003e40000000000000000000000b022000038000fffffffffffdb9ff8f3dd999174bb9c112f2f9177ffffffffffffffffdf7a27a845d671cbdc2ff931820b80000000000000000000000000000000
G0[364] <= 640'h98001da800000000000000000000020280000001ffffffffffffffb1ff8ffe2c48075294c00082fc03ffffffffffffffffffbfc273007ea72cee43f1931c04500400000000000006000000000200000
G0[365] <= 640'he0000060000000000000000000000202800000003ffffffffffffbe0fe0ffa1005077d90614b93fc17fffffffefffffffffefec23740745328de436f9a2200c00000000000000000000000000000000
G0[366] <= 640'hc000003fc0000000000000000000020200000000100003fffffffb79fffffc100447ff33200ba0fc0bfffffffefffffffeff3fd226667c012cdf47bd9c3240c00000000201000000000000000000000
G0[367] <= 640'h7f80000000000000000002028000000000000003e7fffa1bffffff0854877041000800f443ffffffff7ffffffffdb7405a5b35200cbf8ebf994c244c0000000000000000000000000000800
G0[368] <= 640'h18e600000000000000000202000000000000000033fff30dfffffc00488441836848016247f8ffffff7ffffffffd92c20f31227a1a7f8bdf904004040000000800000000000000000000800
G0[369] <= 640'h19c0000000000000000b02000000000000000003ffe205fdfffc082a9201a0808c413019dc7fffffffffffffff9ec904209f5e027e414f040210100000000000000000000000000100000
G0[370] <= 640'h7e042200000000000203100000000000000003ffc107fdffdc880d120580800c01b81b7dffffffefffffffef8d0002149ca30a7cc6af9e2420480000000300000000000000000000000
G0[371] <= 640'h21f80000000000000b00c00800000000000001ffc202f9fe9c400498c500401401a449fd7fffffbffffffe619000209b9cd31e4dcfc79860041c0001900000000000000000000000000
G0[372] <= 640'hcff180000000007e00600000000000000000ffc205f0ecc80080929020a010400049fd7fffffbffffdbe101380008f084b1e4b09979c0602300000921000000000000000000020000
G0[373] <= 640'h20ee00000000100001c00000780000001c3ff8407fccc88006096a060c0100120099c7ffff797ffddfe7003200026190916574c33960bc0800000400000000000000000000000000
G0[374] <= 640'h3c6000000100000800000000700003fffc04967cc8000002062260d0000860037cffffffdffffbdf2001000002558986274d39b621e0380000000000000000000000000000000
G0[375] <= 640'h139c000001000008000000000007fffff8020464c800000000804000100960487d7fffffefffff9c31000000c04001160b420d943880300000000000000000000000000000000
G0[376] <= 640'h6c000010000080000006007e811fff0420c71c800000011088800200000083e7ffffff7bfed9400008000118c8492508096807800000000100000000000000000000000000
G0[377] <= 640'h3dc001000008000000003ffc1fe600c00800c0040000080000300000040c7e7fffffe7ffff040000000000c0801224c31f124000000000001000000000000000000000000
G0[378] <= 640'h23c08c0001000000001fefc1fe600001840c002000009c000001000120cecfffffff7ffff00000000000764008c734e84000000180000000000000000000000000000000
G0[379] <= 640'h3e08000100000001fc00000003000080240000000030400000800300dd6ffffffb7ffff80000000000024001cf00800024800000000000000000000000000000000000
G0[380] <= 640'h1b7c000100000003f8000000018020002000800220b10800008010004c4ffffefd7ff79800000000000060010040005924000000000000000000000000000000000000
G0[381] <= 640'h180001000000ffe1000000020060003000801020220000c080000108dfffff7d3ffed000000000000000000070205004000000000200000000000000000000000000
G0[382] <= 640'h187c000c0c0000000020000400000000000420004404006410007ffff8e3fff4000000000000000003208001000000000000000000000000000000000000000
G0[383] <= 640'h1cfe08080000010800300004000000000049018010000000000003fffe72f070000000000000000013900000000000000000000000000000000000000000000
G0[384] <= 640'hf8780000000010008900400000000010000800030000000010001ffff32e0d0000000000000000008880000000000000000000000000000000000000000000
G0[385] <= 640'he4000000000013180004000000800000020000000004000001ffff808000000000000000000000440400000000000000000000000000000000000000000
G0[386] <= 640'h30200000000000180000000000000000100000000000000001ffff010000000000000000000000000000000000000000000000000000000000000000000
G0[387] <= 640'he00000000000e8000000000000000000000020000000000803d00000010000000000000000000000000000000000000000000000000000000000000000
G0[388] <= 640'h32000000001f80010000000000000326000000000000000000001004120000000000000000000000000000000000000000000000000000000000000000
G0[389] <= 640'hc00000000f0000000000000200002244000000000000000073e001c080000000000000000000000000000000000000000000000000000000000000000
G0[390] <= 640'h3000000ffc000000000000000000230400000000000000000080208000000000000000000000000000000000000000000000000000000000000000000
G0[391] <= 640'h1c00003000000000000000400008008000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000
G0[392] <= 640'h374003000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[393] <= 640'h12cddf000000000000000000002008080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[394] <= 640'h80000000000000000000000c010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[395] <= 640'h0
G0[396] <= 640'h0
G0[397] <= 640'h0
G0[398] <= 640'h0
G0[399] <= 640'h0
G0[400] <= 640'h0
G0[401] <= 640'h0
G0[402] <= 640'h0
G0[403] <= 640'h0
G0[404] <= 640'h0
G0[405] <= 640'h0
G0[406] <= 640'h0
G0[407] <= 640'h0
G0[408] <= 640'h0
G0[409] <= 640'h0
G0[410] <= 640'h0
G0[411] <= 640'h0
G0[412] <= 640'h0
G0[413] <= 640'h0
G0[414] <= 640'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[415] <= 640'h60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[416] <= 640'h8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[417] <= 640'h3000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[418] <= 640'h800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[419] <= 640'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[420] <= 640'h40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[421] <= 640'h0
G0[422] <= 640'h0
G0[423] <= 640'h0
G0[424] <= 640'h0
G0[425] <= 640'h0
G0[426] <= 640'h8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[427] <= 640'h0
G0[428] <= 640'h0
G0[429] <= 640'h1f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G0[430] <= 640'h0
G0[431] <= 640'h0
G0[432] <= 640'h0
G0[433] <= 640'h0
G0[434] <= 640'h0
G0[435] <= 640'h0
G0[436] <= 640'h0
G0[437] <= 640'h0
G0[438] <= 640'h0
G0[439] <= 640'h0
G0[440] <= 640'h0
G0[441] <= 640'h0
G0[442] <= 640'h0
G0[443] <= 640'h0
G0[444] <= 640'h0
G0[445] <= 640'h0
G0[446] <= 640'h0
G0[447] <= 640'h0
G0[448] <= 640'h0
G0[449] <= 640'h0
G0[450] <= 640'h0
G0[451] <= 640'h0
G0[452] <= 640'h0
G0[453] <= 640'h0
G0[454] <= 640'h0
G0[455] <= 640'h0
G0[456] <= 640'h0
G0[457] <= 640'h0
G0[458] <= 640'h0
G0[459] <= 640'h6000000000000000000000000000000000000000000000000000000
G0[460] <= 640'h0
G0[461] <= 640'h0
G0[462] <= 640'h0
G0[463] <= 640'h0
G0[464] <= 640'h0
G0[465] <= 640'h10000000000000000000000000000000000000000000000000
G0[466] <= 640'h12010000000000000000000000000000000000000000000
G0[467] <= 640'h0
G0[468] <= 640'h0
G0[469] <= 640'h88000000000000000000000000000000000000000000000
G0[470] <= 640'h0
G0[471] <= 640'h0
G0[472] <= 640'h0
G0[473] <= 640'h0
G0[474] <= 640'h0
G0[475] <= 640'h0
G0[476] <= 640'h0
G0[477] <= 640'h0
G0[478] <= 640'h0
G0[479] <= 640'h0
end
always @(posedge vga_clk) begin
G1[0] <= 640'h0
G1[1] <= 640'h0
G1[2] <= 640'h0
G1[3] <= 640'h0
G1[4] <= 640'h0
G1[5] <= 640'h0
G1[6] <= 640'h0
G1[7] <= 640'h0
G1[8] <= 640'h0
G1[9] <= 640'h0
G1[10] <= 640'h0
G1[11] <= 640'h0
G1[12] <= 640'h0
G1[13] <= 640'h0
G1[14] <= 640'h0
G1[15] <= 640'h0
G1[16] <= 640'h0
G1[17] <= 640'h0
G1[18] <= 640'h0
G1[19] <= 640'h0
G1[20] <= 640'h0
G1[21] <= 640'h0
G1[22] <= 640'h0
G1[23] <= 640'h0
G1[24] <= 640'h0
G1[25] <= 640'h0
G1[26] <= 640'h0
G1[27] <= 640'h0
G1[28] <= 640'h0
G1[29] <= 640'h0
G1[30] <= 640'h0
G1[31] <= 640'h0
G1[32] <= 640'h0
G1[33] <= 640'h0
G1[34] <= 640'h0
G1[35] <= 640'h0
G1[36] <= 640'h0
G1[37] <= 640'h0
G1[38] <= 640'h0
G1[39] <= 640'h81000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[40] <= 640'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[41] <= 640'h0
G1[42] <= 640'h0
G1[43] <= 640'h40010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[44] <= 640'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[45] <= 640'h1800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[46] <= 640'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[47] <= 640'h800008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[48] <= 640'hc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[49] <= 640'h4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[50] <= 640'h4000000000000000000000000000000000000000000000000000000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[51] <= 640'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[52] <= 640'h800000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[53] <= 640'h4000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[54] <= 640'h4120000100008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[55] <= 640'h1920100101208000000000000000000000000000000000000001000000060000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[56] <= 640'h800400c31101803000000000000000000000000000000000000000008c70801000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[57] <= 640'h800700008018010000000000000000000000000000000000000000000000800000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[58] <= 640'h10000100018210400000000000000000000000000000000000000180100800000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[59] <= 640'h16010200c003b8400000000000000000000000000000000000000018300000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[60] <= 640'h103000018008ee0f8000000000000000000000000000000000000012000026000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[61] <= 640'h2000080008c6000000000000000000000000000000000000000182000026000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[62] <= 640'he0001803000c0300660000000000000000000000000000000000000000322000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[63] <= 640'hc60600c000831f0098668488010000000000000000000000000000000303327e00000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[64] <= 640'hef8c8000cde066300600000000000000000000000000000000800b200007000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[65] <= 640'hec08f000c9ea666004011000000000000000000000000000000001303000100000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[66] <= 640'h84078f008c0fb6c60f80190000000000000000000000000000000012c0010000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[67] <= 640'h1fc03cd9381f333ec60480000000000000000000000000000000040010c030e000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[68] <= 640'hf0f0f138e0713ef3809800000000000000000000000000000004000707300600000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[69] <= 640'h71c39130f071f3fbc8d88000000000000000000000000000000400060f302e00000100000000000000000000000000000000000000000000000000000000000000000000000000
G1[70] <= 640'h33c339f0e17fb3fbfef0800000000000000000000000000101000090c0306400000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[71] <= 640'h333c79f0033f38df0fe60000000000000000000000000080010d00960178e600400000000000000000000000000000000000000000000000000000000000000000000000000000
G1[72] <= 640'h80c166cef8001b3c9c73f100040000000000000000000000008000201f10def800000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[73] <= 640'hf077eff7fc1f10087fff900800000000000000000000000000030000030780e00000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[74] <= 640'hc077eff7fe1030081ff748c80000000000000000000000001101080000131c000000000000000000020000000000000000000000000000000000000000000000000000000000000
G1[75] <= 640'hc060ffffffe10bc030fee49c00000000000000000000000000000080010131c000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[76] <= 640'h763dffffff0f8f83bffe670000000000000000000000000000000010000310600000100000000000000000000000000000000000000000000000000000000000000000000000000
G1[77] <= 640'h1c673ffffffffd3043ffff700000000000000000000000000000060000003fc400000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[78] <= 640'h3c67ffffffff9fc1e1ffcfc080000000000000000000000000000fc000003fe000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[79] <= 640'h27ec1fffff79fc73fff81800c000000000000000001210000010f07010c1fcfc0008000000000000000000000000000000000000000000000000000000000000000000000000000
G1[80] <= 640'h367ffffdffef9ffe7fff8101040800000000000000000000010308001000fbf00000000000000000000000000000000000008000000000000000000000000000000000000000000
G1[81] <= 640'h3862ffffffff7ffffffffe8199000000000000000000000000100f8000001fff00000000000000000000000000000000000000800000000000000000000000000000000000000000
G1[82] <= 640'h811870ffffffff3f7f7fffffc08f00000000000000000000000080000000003fffe0000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[83] <= 640'h3f0ffff7ffffe7f7ffffffc8e00000000000000000000000080804000033fffff000000000000000000000000000000000008000000000000000000000000000000000000000000
G1[84] <= 640'h10c1c3fffffffffe7ffffffffe9c00000000000000000000000000074000037fffe0800000000000000000000000000000000018000000000000000000000000000000000000000000
G1[85] <= 640'h3dcf3fffffffffffffffffe79c800000000000000000008000020200003cfffff08000000000000000000000000000000000c0700000000000000080000000000000000000000000
G1[86] <= 640'h1fdf3ffffffffffffffffff3ff98e000000000000000600000020000003fffffff8000000000000000000000000000000000c3030000000000000080000000000000000000000000
G1[87] <= 640'h81fcffffffffff7fffffff78fb99e4c00000000000003001010200800003ffffff44000000000000000000000000000000011c000000000000001000000000000000000000000000
G1[88] <= 640'hffeeffffffffefffffffffff7e7103800000000000001800000107000c1ffffffcc08000000000000000000000000000000118700000000000000e1c000000000000000000000000
G1[89] <= 640'h1fefffffffffffffffffffff76f3c0000000000000000400c30100f0493fffffefc0010000000000000000000000000000000f39c000000000001c00000000000000000000000000
G1[90] <= 640'h103f7ffffffffffffffffffff7eff8100000000000000e000000000f0693ffffff7c0000000c0001c00000000000000000000837fc0000000000000c3000000000000000000000000
G1[91] <= 640'h103f3ffffffffffffffffffffffff8180000000000001e0001c0000f06d7ffffff8e160811fe0003fc000000000000000000038ff000000008000c1c3008000000000000000000000
G1[92] <= 640'h10033f3fffffffffffffffffffffffef0800000000000006600100000f84cfffffffff102000fe00033e00000010000000000003ffff00000000000e100808000000000000000000000
G1[93] <= 640'h337ffffffffffffffffffffffffe80000000000000013f00000000f8cc7ffffffff100180fe300277c00000000000000000077fff800000038003c00c00600000000000000000000
G1[94] <= 640'h33bfffffffffffffffffffffffff00000000000000019830c3070000cd3ffffffffff000ffff00fffe00000000000000000063fffc0000007800309f7c0e00000000000000000000
G1[95] <= 640'hf33ffffffffffffffffffffffffe7000000000000000019100007c031ed3ffffffffe9900e3ff3ffeff00000000000000000007ffff000000031c018e7c0cc0100000000000000000
G1[96] <= 640'h1000000000000038fffffffffffffffffffffffffcc80000000000000003f77600c7086ff7e9ffffffcb2c766feffff7f000000000000000001bffffec00000100080ffcf0c18000100000000000000
G1[97] <= 640'hfffffffffffffffffffffffff4c0000000000000000f838708f78c67e7effffffffbefe07fffffffe000000000000000000b9fffcc00000000000ffff0019000000000000000000
G1[98] <= 640'hc0fffffffffffffffffffffffff4c0100000000000000f83060fffee07c7ffffffffffffe9ffffffffe000000000000000001f90ff9600000000003ff738001000000000000000000
G1[99] <= 640'hc0effffffffffffffffffffffff4c00000000000000003f30e3ffff70e7fffffffffefffff9ffffffffc00000000000000001f967f9600000000003ff7fc0c2800000000000000000
G1[100] <= 640'h6f0ffffffffffffffffffffffffcd0000000000000000f907e7ffff71e7fffffffffffffff9ffffffffe00000000000000001ff6fbf660100380003ffffc7c6800000000000000000
G1[101] <= 640'h7e1ffffffffffffffffffffffffe9c0000000000000003fef7ffffff8fefffffffffffffffffffffffff000000000000000016f7fffe72102e33ce1ffffc7cc800000000000000000
G1[102] <= 640'h6e7fffffffffffffffffffffffff8c4000000000000001ffffffffffffefffffffffffffffffffffffff8000000000000000007ff7fff0026e73fffffffff9c900000000000000000
G1[103] <= 640'h10ec7fffffffffffffffffffffffff88400000000000002f9fff7ffffffe7fffffffffffffffffffffffffc0000000000000000039ffffe00e67fffffffffff99900000000000000000
G1[104] <= 640'h608f7ffffffffffffffffffffffffffc8000000000000007fff7fffffffefffffffffffffffffffffffffffc000000000000000003ffffffb91fffffff7ffff30e300000000000000000
G1[105] <= 640'hdf7ffffffffffffffffffffffffff30000000000000006fffffffffffffffffffffffffffffffffffffffc000000000000000001ffffffd8fffffffffffcff80100000000000000000
G1[106] <= 640'h119f4f7ffffffffffffffffffffffff30100000000000000fefffffffffffffffffffffffffffffffffffffc800000000000000001fffffffcf3fffffffffcfff0000000000000000000
G1[107] <= 640'h117fcffffffffffffffffffffffffffe0000000000000007fffffffffffffffffffffffffffffffffffffffe8000000000000000017fff7fffffffffffffff1cf0000000000000000000
G1[108] <= 640'h81ffcdfffffffffffffffffffffffffe88c0000000000007ffffffffffffffffffffffffffffffffffffffff8000000000000000017fffffffffffffffffff3c78000000000000000000
G1[109] <= 640'h17fcdffffffffffffffffffffffffffdcf800000000001fffffffffffffffffffffffffffffffffffffffff800000000000000001ffffffffffffffffffff7c3c000000000000000000
G1[110] <= 640'h8000337ffdffffffffffffffffffffffffffff8800000000001fffffffffffffffffffffffffffffffffffffffff800000000000000001fffffffffffffffffffffe00000000000000000000
G1[111] <= 640'h3000377ffdffffffffffffffffffffffffff7f9c00000000001ffffffffffffffffffffffffffffffffffffffffff8810000000000000f7ffffffffffffffffffefc00010000000000000000
G1[112] <= 640'h86000007ffeffffffffffffffffffffffffffffefc08000020000fffffffffffffffffffffffffffffffffffffffff84000000000000000effffffffffffffe7feffe000000000000000000000
G1[113] <= 640'h1000007fffffffffffffffffffffffffffffffff400000000003fffffffffffffffffffffffffffffffffffffffffce800000000000000ffffffffffffffffffffc0000000000000000000000
G1[114] <= 640'h3104000ffffbffffffffffffffffffffffffffffe660000000003ffffffffffffffffffffffffffffffffffffffffffff000000000000007ffffffffffffffffe7ec0000000000000000000000
G1[115] <= 640'h3100003ffff9ffffffffffffffffffffffffffffe760000080001fffffffffffffffffffffffffffffffffffffffff7ffd80000000000003ffffffffffffffffe3040000000000000000000000
G1[116] <= 640'h300003ffffbfffffffffffffffffffffffffffffe40000000001fffffffffffffffffffffffffffffffffffffffff7fff00000000000003ffffffffffffffffec000000000000000000000000
G1[117] <= 640'h8730003ffffffffffffffffffffffffffffffffffe00008000000fffffffffffffffffffffffffffffffffffffffff7fff00000000000003ffffffffffffffffdc000000000000000000000000
G1[118] <= 640'h10000def0003ffffffffffffffffffffffffffffffffffe010000000007fffffffffffffffffffffffffffffffffffffffffffec0000000000003fffffffffffffffef8000000000000000000000000
G1[119] <= 640'h3fec0003fffffffffffffffffffffffffffffffffff910000000007fffffffffffffffffffffffffffffffffffffffffffe0000000000000739fffffffffffffff0800000000000000000000000
G1[120] <= 640'h19ff0803fffffffffffffffffffffffffffffffffff00010000001fffffffffffffffffffffff7fffffffffffffffffffffc8000000000000f03ffffffffffffbe0000000000000000000000000
G1[121] <= 640'h810081fff9007efdfffffffffffffffffffffffffffffffcc0000000800fffffffffffffffffffffffffffffffffffffffffffffc8000000000003000bfffffffffffde0000000000000000000000000
G1[122] <= 640'h8001fff90067cff3ffffffffffffffffffffffffffffffc00001000103ffffffffffffffffffffffe7ffffffffffffffffffffec0000000000030003e3ff7ffffffc80000000000000000000000000
G1[123] <= 640'h800cfff8007ffffffffffffffffffffffffffffffffc3fc08001000003ffffffffffffffffffffffffffffffffffffffffffffec0000000000000000c1fffffffffc00000000000000000000000000
G1[124] <= 640'h3900f87ff8007f7ffffffffffffffffffffffffffffffc80000000000001fffffffffffffffffffffffffffffffffffffffffffffe400000000000000000fffffffff300000000000000000000000000
G1[125] <= 640'hc101c0dffd003ffffefffffffffffffffffffffffffce180000000000001ffffffffffffffc7dfffffe3ffffffffffffffffffffffe800000000000000061f3ffffff000000000000000000000000000
G1[126] <= 640'h800387dffd001ffffffffffffffffffffffffffffffff3000000000000007fffffffffffee011ffffff3ffffffffffffffffffffffe80100000000000006113fffff6000000000000000000000000000
G1[127] <= 640'he0ff8dff803ffcfffffffffffffffffffffffffffff7c080000000000007fffffffffffee001fffff7fffffffffffffffffffffffefc100000000000000003fffff4000000000000000000000000000
G1[128] <= 640'hc799fb9efee436fbffffffffffffffffffffffffffffcc800000000000017ffffffffffecc003ffffffffffffffffffffffffffffff9e40068000000000004077ff9c000000000000000000000000000
G1[129] <= 640'h1cfff91fbf4c27ffffffffffffffffffffffffffffffff180000000000007ffffffffffff0000fffffffffffffffffffffffffffffff660000000000000000073ff00000000000000000000000000000
G1[130] <= 640'h3fff9f7ff29ca7feffffffffffffffffffffffffffffff180000000000007fffffffffff70000ffffffffffffffffffffffffffffffffc00000000000000000178000000000000000000000000000000
G1[131] <= 640'hfffffffffa9816fffffffffffffffffffffffffffffffec00000000000007fffffffffff700007fffffffffffffffffffffffffffffffce44000000000000000fd000000000000000000000000000000
G1[132] <= 640'hffffffffff8106fffffffffffffffffffffffffffffffe030000000000067fffffffff7ecc0007ffffffffffffffffffffffffffffffffe6cc0080000000000000800000000000000000000000000000
G1[133] <= 640'hffffffffff8187fffffffffffffffffffffffffffffffc0e000000800006fffffffffd7fcc0017ffffffffffffffffffffffffffffffffffdc0080000000000000000000000000000000000000000000
G1[134] <= 640'hffffffffff6287fffffffffffffffffffffffffffffff8fc000000000086fffffffffdffe0001ffffffffffffffffffffffffffffffffffffc0000000000000000000000000000000000000000000000
G1[135] <= 640'hffffffffff749ffffffffffffffffffffffffffffffdffef0000000000c6fffffffffffff1001ffffffffffffffffffffffffffffffffffffdc181200000000000000000000000000008000000000000
G1[136] <= 640'hffffffffffdb7ffffffffffffffffffffffffffffffffeed200011e17077fffffffffffff8007fffffffffffffffffffffffffffffffffffffce71000000000002000000004000000000000000000000
G1[137] <= 640'hfffffffffff97ffffffffffffffffffffffffffffffffffdf80011703e7ffffffffffffff88c7fffffffffffffffffffffffffffffffffffffff3f700000000000000000000000000000000000000000
G1[138] <= 640'hfffffffffff9ff7ffffffffffffffffffffffffffffffffffc00fbfe8ffffffffffffffffc8cfffffffffffffffffffffffffffffffffffffffffff00000000000000000000000002000000000000000
G1[139] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffdec4eeffc7fffffffffffffffe99fffffffffffffffffffffffffffffffffffffffffff8c000000000000000000000000000000000000000
G1[140] <= 640'hfffffffffffdffffffffffffffffffffffffffffffffffffff00feffcffffffffffffffffe9bfffffffffffffffffffffffffffffffffffffffffffec000000000000000000000000200000000000000
G1[141] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffcfff7ffeffffffffffffffff73fffffffffffffffffffffffffffffffffffffffffffee000000000802000000000000000000000000000
G1[142] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff77fffffffffffffffffffffffffffffffffffffffffffef800000000000000000000000000000000000000
G1[143] <= 640'hfffffffffffeffffffffffffffffffffffffffffffffffffffff9ff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff880000000000000000100003001000000000000
G1[144] <= 640'hfffffffffffeffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000000000600800001010000000000
G1[145] <= 640'hfffffffffffefffffffffffffffffffffffffffffffffffffffdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000000000000000e0e10680000000000000
G1[146] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff89000000000000000000007367c0000000000000
G1[147] <= 640'hffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf0000000000000000000373773f240000000000
G1[148] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffe800100000000000000008f73ff060000000000
G1[149] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffece010800000000000000dfffff0e8000000000
G1[150] <= 640'hfffffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff73ffffffec7800000000000000003ffffffdc0000000000
G1[151] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7fdffff7fcf8000000000000000f3fffffffc0080000000
G1[152] <= 640'he7ddffffffffffeffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffefff1300000000000001ffffffffb8000000000
G1[153] <= 640'h7e9fffffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc600000000000000cffffffffe8800000000
G1[154] <= 640'h7cff7fffffffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe8e00000000000000dffffffffe0800000000
G1[155] <= 640'he77f7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe1ec00000000000001ffffffffe0000000000
G1[156] <= 640'he33f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff79e00000000000003fffffffe6c000000000
G1[157] <= 640'he67cfffffffffffdfcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff73c00000000000003fffffffe6c000000000
G1[158] <= 640'h64d87ffffffffffc313ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb00000000000000fffffffeff0000000000
G1[159] <= 640'he70f3feffffffffc03e7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff00000000000000ffffffffff6400000000
G1[160] <= 640'hf307bfdffffffffc001bffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9c780000000003fffffffffff000000000
G1[161] <= 640'h7807fffffefffffc00017fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff88180000000071fffffffff700f0000000
G1[162] <= 640'h3847fffffefffffe00197fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1000000000023ffffffffffdc00000000
G1[163] <= 640'h91e4b3ffffffffff0039ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7c00000000003ff7ffffffefc00000000
G1[164] <= 640'h817cb7ffffffffff00397ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec000000000e0ffffffffff0ee0000000
G1[165] <= 640'h987ef77ffefeffffe000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec000000000ffffffffffffce00000000
G1[166] <= 640'h1c6ff77ffeffffffc001f3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee0000000013ffffffffffff80f000000
G1[167] <= 640'h9d4023e3e7ff7fff80017fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffff0000100017efffffffffee380000000
G1[168] <= 640'h63901cffffdfcffc20087fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe204000003e7ffffffffffc1c0000000
G1[169] <= 640'h7c02007fff9fffffe00107fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000007fffffffffffffe1c000000
G1[170] <= 640'h5c32c033f36ff3ff030107fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc4000040ffffffffffffffc0c000000
G1[171] <= 640'h88f0c339e367733c07003efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000006fffffffffffffffc83800000
G1[172] <= 640'h89b01f9fff40011c6000389ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000167fffffffffffffff8c1000000
G1[173] <= 640'hd021f9efe4084c6408003bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00377fffffffffffffff330180000
G1[174] <= 640'h7d861cdffed884c3068001bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc8fffffffffffffffeffff30000000
G1[175] <= 640'h659e00f3ff9900000010001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffff1ffffefffffffffddf7cfc03800000
G1[176] <= 640'h27ce3cddffe011000000007fdfffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffff7fffffffffffffffffffffffffffffffffffffeef9feeefffffdfffff081800000
G1[177] <= 640'he7cfefdffc000000000000e7dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7e08000000
G1[178] <= 640'he7ffffbffc00002000000067ff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3ffffff08000000
G1[179] <= 640'hffffff7fff0000000000003cfb7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffcff7effffe81300000
G1[180] <= 640'h7fffffffff00000600000018937ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdff3fff4dfffec0000000
G1[181] <= 640'h7effffffbe800004000000000373ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffeedff7fbc601000
G1[182] <= 640'h7fffffffff000100000000010907fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffefdff3f98600000
G1[183] <= 640'h2ffffeefff000000000000189817fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec3cf68ff6683000000
G1[184] <= 640'h3fffffffff80000080000000186ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefc6799008cc7010000
G1[185] <= 640'hffffffffffc00000800000000007fcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffe7183c0046000000
G1[186] <= 640'hffffffffffe00000000000000001f8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7f63c083104000000
G1[187] <= 640'hffffffffffe000000000000000113fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff606187108000000
G1[188] <= 640'hfffffffffff000001000000000193fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee46fee0dc000000
G1[189] <= 640'hfffffffffff0810030000000000067fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeef60fcc080000000
G1[190] <= 640'hfffffffffffc0360b0000000000067ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff8808400000000
G1[191] <= 640'hfffffffffffec060f000000000046efffffffffff7ffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef81c00198000000
G1[192] <= 640'hffffffffffff3bf3f800000000043f73ffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1fe783000001800
G1[193] <= 640'hfffffffffffff93ab800000000003b73ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7e030020000000
G1[194] <= 640'hffffffffffffffbebc000000000078e7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff67810000000000
G1[195] <= 640'hfffffffffffffffffc80000000001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ef88000000000
G1[196] <= 640'hfffffffffffffff7fc00000018010fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7c0c0480000000
G1[197] <= 640'hffffffffffffffffff00000000800c3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7c008400800000
G1[198] <= 640'hffffffffffffffffff70000081800e3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefec0c000800000
G1[199] <= 640'hffffffffffffffffff00600801810f37ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff7000400000000
G1[200] <= 640'hffffffffffffffffff30010006600c3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7effffffffffffffffffffffffffffffffffffe6e60190800000
G1[201] <= 640'hffffffffffffffffffe1c00106e6f8fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff07e0000000000
G1[202] <= 640'hffffffffffffffffffe70004c7fff8fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9660000000000
G1[203] <= 640'hffffffffffffffffffff0f08ff9f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbc3f000000000
G1[204] <= 640'hfffffffffffffffffff9200c3f9f7fffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe73010000000
G1[205] <= 640'hfffffffffffffffffff8f01f7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff0013000000
G1[206] <= 640'hfffb7fdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef80000000080
G1[207] <= 640'hfffc2689fffffffffffffffffffffffffffffef3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7c10098000000
G1[208] <= 640'hfff9670004ffffffffffffffffffffffffffe7d8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffee34114000000
G1[209] <= 640'hfff97600001ff9ffffffffffffffffffffff7fff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe6f01904000000
G1[210] <= 640'hffffe000000efcfffffffffffffffffffffffddfffffffffffffffffffffffffffffffffffffffffffff310380ffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7f81984000000
G1[211] <= 640'hff7fc0000000b83ffffffffffffffffffffffdfffffffffffffffffffffffffffffffffffffffffffffe0080000fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f8100000000
G1[212] <= 640'hff7ee0000000001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000001ffffe3c00ffffffffffffffffffffffffffffffffffffffffffffffeff8003000000
G1[213] <= 640'hfffe78000000000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000ffffe00003fffffffffffffffffffffffffffffffffffffffffffffff67c00800000
G1[214] <= 640'hfffebc0000000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe100000000fffe6000001ffffffffffffffffffffffffffffffffffffffffffffffc7c80800000
G1[215] <= 640'hffff8800000000007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000fffe000000007ffffffffffffffffffffffffffffffffffffffffffffe6c80c00000
G1[216] <= 640'hffffc000000000017ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000f00000000001fffffffffffffffffffffffffffffffffffffffffffffb2845400a0
G1[217] <= 640'hd3ffe00000000000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0f800000000000000000000000fffffffffffffffffffffffffffffffffffffffffffff5244140000
G1[218] <= 640'h807e8000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe38c000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffff7244140040
G1[219] <= 640'h2600000000000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3000000000000000000000000000004ffffffffffffffffffffffffffffffffffffffffffda244150040
G1[220] <= 640'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2000000000000000000000000000000dfffffffffffffffffffffffffffffffffffbffffffa004908010
G1[221] <= 640'h3fffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000017ffffffffffffffffffffffffffffffffff3ffffffe100140010
G1[222] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000000000000000000000017ffffffffffffffffffffffffffffffffffbffffff7130160080
G1[223] <= 640'hc000000000ffffffffff7ffffffffffffffffffffffffffffffffffffff9fffffe00000000000000000000000000000001ffffffffffffffffffffffffffffffffffff7ffffff582360049
G1[224] <= 640'h39c0000000003fffffff3ffffffffffffffffffffffffffffffffffcf9f0cfffffb000000000000000000000000000000003fffffffffffffffffffffffffffffffffb97d6fffd09220b281
G1[225] <= 640'h7dc0000000000fffffff1ffffffffffffffffffffffffffffffffffcfffc1fffffc800000000000000000000000000000001ffffffffffffffffffffffffffffffffff759ffffd302649201
G1[226] <= 640'h7fe00000000003cffff71ffffffffffffffffffffffffffffffffffcfffc13fff7c000000000000000000000000000000000ffffffffffffffffffffffffffffffffed94dfffec3804cb0a0
G1[227] <= 640'hffe8000000000181cff00fffffffffffffec3c7ffffffffffffffffcfe7c33eff3c0000000000000000000000000000000007fffffffffffffffffffffffffffffffed4dd7feec1484c3c90
G1[228] <= 640'hfff00000000000000f800ffffffffffffff8103ffffffffffffffffeee7833effc00000000000000000000000000000000003fffffffffffffffffffffffffffffffeded3fffec10a042c90
G1[229] <= 640'h1fff000000000000002000ffffffffffffee0001ffffffffffffffffdc7f081cffc00000000000000000000000000000000003fffffffffffffffffffffffffffffffe4cd2fffe6092246ad0
G1[230] <= 640'h2ffff0000000000000000003fffffffffffe000000ef3ffffff9fb9f8fcbf00083fe00000000000000000000000000000000003ffffffffffffffffffffffffffffffff65916ffaf0c824ea40
G1[231] <= 640'hffffc000000000000000001fffffffffffc000000021fc00ff8319009c99000107780000000000000000000000000000000003fffffffffffffffffffffffffffffffff29a7ffa70c049a640
G1[232] <= 640'h17ffff0000400000000000007ffffffffff00000000200100b80000000638010080000000000000000000000000000000000001ffffffffffffffffffffffffffffffff79827ff6f080090658
G1[233] <= 640'h1fffff0000c00000000000007fffffffc38000000000000000000000006bc000000000000000000000000000000000000000001ffffffffffffffffffffffffffffffff0c446ff4d01120464c
G1[234] <= 640'h1e7ff00000000000000000001fffffffc00000000000000000000000000000000000000000000000000000000000000000000007fffffffffffffffffffffffffffffff2044dfe4605a204c24
G1[235] <= 640'he0000003fff8000000000000000000007ffffff800000000000000000000000000000000000000000000000000000000000000000000007fffffffffffffffffffffffffffffff19116ff62868218526
G1[236] <= 640'hf80000017cf03e8000000000000000003fffff0000000000000000000000000000000000000000000000000000000000000000000000007bffffffffffff073fffffffffffffef90133ff6242c232402
G1[237] <= 640'h7c8e00203cff7ce000000000000000003fffff000000000000000000000000000000000000000000000000000000000000000000000000fbffffffffffe0033fffffffffffffefce145df72001210900
G1[238] <= 640'hfc8c0000003fc00020000000000000001ffff8000000000000000000000000000000000000000000000000000000000000000000000000fffffffffffe00000fffffffffffffeec4c41ff71889014308
G1[239] <= 640'hff080000000fe10020000000000000000ffff8200000000000000000000000000000000000000000000000000000000100000000000000fffffffffffe000003ffffffffffff6ea0ce1dda188906c948
G1[240] <= 640'h100000000000000000000000000000001dff0000000000000000000000000000000000000000000000000000000000000000000000000f87ffffffffb000083afffffffffff2f700e5ffb10b004d92e
G1[241] <= 640'h8ef00000000000000000000000000000000000000000000000000000000000000000000000000000ffffffe0000001affffffffffd93380e01f31a400c5804
G1[242] <= 640'hc000000000000000000000000000000000000000000000000000000000000000000000000000000fffff000000002ffffffffffc238c4c7df18411164004
G1[243] <= 640'h80000000000000000000000000000000000000000000000000000000000000000000000000000000fff00000000017ffffffffffdbc41028f8a831788506
G1[244] <= 640'h18700000000057ffffffffffc7c22461f81798422420
G1[245] <= 640'h3efffbffffe2a201461780b4c023012
G1[246] <= 640'h36fef9ffffe018815a87c4bc446313b
G1[247] <= 640'h36fff2ffffc2a8010a1ffa3e4071989
G1[248] <= 640'h2baebf2ffff81de43060fe0002021031
G1[249] <= 640'h146dfeaefff3c381b147dd802c0ad010
G1[250] <= 640'hfc0000000000000000000000000000b34ffc77df3027610027ddbc76289052
G1[251] <= 640'hfe000000000000000000000000000139ceb8855f16f1941857bff40c802081
G1[252] <= 640'h1fe0000000000000000000000000001122daade7f13740c926fbe58e812b0e8
G1[253] <= 640'h3ff00000000000000000000000000016e6dfac7febb6245220a9d80b35ab0ec
G1[254] <= 640'h1f8000000000000000000000000000000000000000000000001fffff800000000000000000000000012899fb99ff912642a402148124119964
G1[255] <= 640'h1fc0000000000000000f0000000000000000000000000000003fffffc000000000000000000000000052d9bed1ffcf0e79028a2fe0b0324490
G1[256] <= 640'h1fe0000000000000003e80000000010000000000000000000007fffff00000000000000000000000059e87ca55ff474a0b88c131e80f28c480
G1[257] <= 640'h1ff8000000000000003fe0010700ffc0000000000000000107fffffffc0000000000000000000000049b254212bfe56207a09183f847602402
G1[258] <= 640'h3f7c00000060000006ffe007fffffff800000000000007e007fffffff0000000000000000000000002cd7f7b63ffc077cf910017b904239040
G1[259] <= 640'h380000000100000000000000000001fffc000030e000001ffff00ffffffffffffffc0000001ff807ffffffc000000000000000000000000147e143bbefb730c4408b907dc0068090
G1[260] <= 640'h3fe3000000001f0000000000000001ffff0000790000003ffff80fffffffffffffff04001ffffeffffffffc0000000000000000000000001a9baa916e94f9a4b44902bfe602bc320
G1[261] <= 640'h1fffc8000001ffe000000000000001ffff80007f0000007ffffc0fffffffffffffffc7fffffffffffffffffc440000000000000000000008955d2e16b4e4331240a0867819364258
G1[262] <= 640'h1fffe000007fffe00000000000001ffff8000fff00000ffffff7fffffffffffffffffffffffffffffffffffff8000000000000000000084e823000c162e60014131a03770112404
G1[263] <= 640'h1ffe054007ffff98000000000000fffe800fffff0007ffffffffffffffffffffffffffffffffffffffffffffc0000000001c00000000a23150352c264d5c10a6550bef023342bc
G1[264] <= 640'hffcc0ffffffff000000000001ffff0007fffff83fffffff3ffffffffffffffffffffffffffffffffffffff3817f1fffffff7e7f85a38bea080c603e55ac672e07c530326795
G1[265] <= 640'h73cfffffffffff000000000007fff0007fffffcffffffff3fffffffffffffffffffffffffffffffffffffffffffffffffffffff4504185123002d1f3c9a686a8b25813c2c01
G1[266] <= 640'h1cffffffffffffffffc000003fff0007fffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8105c82308056d3d2c5c184804a8002f7d80
G1[267] <= 640'hf800000000001fffffffffffffffffc007807fffc00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff90404c0411891c9bc6c885981b70043631b9
G1[268] <= 640'hbfff0000000000ffffffffffffffffffc00fff7fffe07fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff60a93c0e802f02f4d7c0ece80bf82ab32281
G1[269] <= 640'hfffffff0000007ffffffffffffffffffc6ffffffffe07ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff12899a0e8122266634121fb10a523a04828
G1[270] <= 640'hffffffff18001fffffffffffffffffffcffffffffff0ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb195fd2e398523c55e1b4cf4003af908b956
G1[271] <= 640'h2fffffffe7ffffffffffffffffffffffffffffffff0fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8f6e56895225d86e380c4198e25bc9804e4
G1[272] <= 640'h57ffffffffffffffffffffffffffffffffffffffffe07fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd447ef85d0123cda4df22f69a48de6421440
G1[273] <= 640'h7fffffffffffffffffffffffffffffffffffffffff07fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff93ad72d98a02137f2c3621144215a499ac34
G1[274] <= 640'hffffffffffffffffffffffffffffffffffffffffff8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddb64b04399b042b9208e6a250999d050618
G1[275] <= 640'hfffffffffffffffffffffffffffffffffffffffffff887ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcdfaf55af8815493cef0274349d61b8946a6
G1[276] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffc07ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffaff0c88350ccc74c3460a4652e1b758c16c0
G1[277] <= 640'h17ffffffffffffffffffffffffffffffffffffffffffefc07ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb1ea1c910cd00637c222e487e208cc8508d2
G1[278] <= 640'hffffffffffffffffffffffffffffffffffffffffffff87c1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3a25f3c8124b02430b80615301a18b4289ed
G1[279] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffff03c1effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9b636fb470c940299b1c92592810c202582c
G1[280] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffff1c0cc7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4e99580784189c6db5a3a790504e14844592
G1[281] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffff1c0eefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa3f6f2224ca5cb63c2a0c20d9626c4407070
G1[282] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffc0e07fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd7cb89b2b289cc3921432a6637eae17013714
G1[283] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffc0e03fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc9be99fa47991c01cb94ab68242f863e37b1e
G1[284] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffff0f00ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc854758f19ee6d81f605814a92e087a42294d
G1[285] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffff8f00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdb5bb6770ee914b780719d5cb489342229e08
G1[286] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff0effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed7e6b7282a601ae3173fcc37ae21ccc909087
G1[287] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefd79ef9f3ac442cb9d1793121642c2930eb41
G1[288] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffff7b7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff74ea26fb66200c0f610441057432a8bd4788f
G1[289] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffff8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ba66d07f608410df037b72792cd563201cb4a
G1[290] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3e70310f52c454884918fd03d332e80973808c
G1[291] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffe79fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9da87d8930c60c0614586102f3e2811973f762
G1[292] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8fae9ae25f6a30643d0d5f037030892909451a
G1[293] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc29ec6f9679710b65bcfaa85bb20fd088083b2
G1[294] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd736d6061e20d8c8cc6fbdc4e2321054a07731
G1[295] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa0fd07ebcbfd48db76733d01a7e47f8ab083a0
G1[296] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5bf638df98219619ee973e49fe54b64a0c684
G1[297] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbc4747e19dbd80710c1dfee6846d1732208f54
G1[298] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffff6f5aae2ca44a89ef8536ef26898f3227201eb2
G1[299] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe17fffffffff4d67290660bed1800b7a6566cb2f86dd316678
G1[300] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0e17fffff7fffa798b5e4840f809daf2576a6463f56005d971c
G1[301] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffe0213fffff1fffc04ed58046e1014ee513bce3af1d6d08444600
G1[302] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3fffffffffffffffffffffffffffffffffffffffffffff00231bf3f447fc20f7ac543aa68d332a341a6307752b66ade816
G1[303] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddffe0fffffffffffffffffffffffffffffffffffffffff000f1bf300c000141982098a788b127bbd22b286883b4bb55507
G1[304] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3ef8783fffffffffffffffffffffffffffffffffffffffc900a099141800082085175cb794364d57883d1f5371e09d86505
G1[305] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfef7f81ffffffffffffffffffffffffffffffffffffffff805e0ac3fff8800c398a64962a276dec1b4131a0f9ead34cb51b
G1[306] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdff8f7f83fffffffffffffffffffffffffffffffffffffffffe9e9644000001360f182cedb301ae30edd4e3ebf4ff3b308c04
G1[307] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3fe00ffdfffffffffffffffffffffffffffffffffffffffffe46de05e000022f10b8400039a63a70485b9725da409c0f0ac3b
G1[308] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff78ffc0fffc5ffffffffffffffffffffffffffffffffffb01f00007ea00879c023b00c46287a9662d3a8d993b1e6d9c1d9d0d8f4
G1[309] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffc03fc0ffffe1fffffffffffffffffffffffffff3fffc000063f0fffd8e0c79c3c77694594bb8c4007b43cd90207cf3f550b81ca8
G1[310] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffff800440f3fff1ffdfffffffffffffffffffffe00000dff81fffffff602e647fffc7903099a9c4c280c9dc1c1440bcd702e04c3481
G1[311] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffd8006fcffff8380fffffffffffe7000007fffffffffffdc0ffffff5a9e40ffffe32200d39a46c6c107edb2b1f1f5325e3704a081
G1[312] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff000f91ffff8fe03fff0c000080001ffffffffffffff03e0ffffff56de44ffff92e5fb032dad70e247a5fc40b2bc83fb55600a64
G1[313] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff804001fffff1ff80c0007fffffff1fffffffffffff0ffc0ffffffab0fadffffdbcfe4a435b731a05f50a0e6432cefc840bc2218
G1[314] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffff800001fcffffff3fe08e0fffffffffffffffffffffffe7ff8fffffffdcdf2dffffefe9de05c3a318c1a47f8e78c0c665d9977c108b
G1[315] <= 640'hfffffffffffffffffffffffffffffffffffffffffffff000000000000001e03fc100fff00021ffff7ffffffffff3ffffffe7003ffffdfe809eb5bfffee43c825c380dc90e23d3348405f630d694e1042
G1[316] <= 640'hfffffffffffffffffffffffffffffffff000000000000000001007ff00000007e3e1fff800007ff967ffffffffffffffffe07ffffffcfe4c3ad53fffd8439a6d796e6ce146beb7e66ae62746d9d4e146
G1[317] <= 640'hfffffffffffff00007fffffff8000000000000ffffffffffffffff1c000000003000fffc017e068463fc0ffffffffffffffffffffffefe52b23f7fffe8a0c52b19722e25ce5cb9fc806de28f2346a8a1
G1[318] <= 640'hfffffffffffffffffffffffffffffffff8800000000000007ffe83ff807f00e3f07ffffffffffffffffffffeef02b7076fffecf348efd41734e2422fb9fd48cd08411112c6d3
G1[319] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffcc0000000000001fff83fff0ff800ffe3ffffffffffffffffffff6499d348021fffa98e96f2031d0c09329bb1aa9ffae37b27ecb0a
G1[320] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000003ffe7ffffffff3fffe00fffffffffffffffbff24c3bfac34bfffa4c3452b81bc0121e98bc2b819d73313794d9f8
G1[321] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000f83fffffffffffffff00ffffffffffffef0fd24b333faf7fffd9615c9e44836002d10837c2c01a3d5e45986134
G1[322] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000000839ffffffffffffffff9fffffffffffe784dd1b773c578fffdfdbe2f5e7b1386031e9321660397645556436c8
G1[323] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000000001ffffffffffffffffe3ffffffffffbf85d8ba5be909edafc7cb27942b80982c0671272f4821f8eb2f087890
G1[324] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000000000007fffffffffffffff87ffffffffffb85841e6d6a8387248925669ca8a524241989537440228a82efe490c4
G1[325] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000000003ffffffffffffffff01ffffffffde63fb5a32acc94e25017973bf8056144cd25e334a814ce622a4b808d3
G1[326] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000004effffffffffffffe003ffffffcccb3ed7425f327605d1e88914dc2b4034161a0ef18104121760da1081
G1[327] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffc0000000000000000000001ffffffffffffff83fffffe5d2d74e1283dededa58867e6c20e25e3322a4f01abc8beaf6c20582807
G1[328] <= 640'h10fff0f7f07ffffffffffffffffffffffffffffffffffffffffffff00000000000000007fffffffffffffffc00c067ffead90233f704fe777a2b13626175ddd3914075d402bc092301303ec0c86
G1[329] <= 640'h1000000000000000000000000000000000000000000000000000000000000000000000000703ffffffffffc60fffffe0b64ac73aa633035bb4846a5a232e30806155004d0c826d42949e81096
G1[330] <= 640'h7fffffffffffffffffff00000000000000000000000000000000ff8000ff60000000000000000000000ffe0000c0fc307ffffea39434379d5fae716c46ea99cbab33ac121a267be59033a59ae0943687
G1[331] <= 640'h10000000000000000007ffffffffffffffffffffffffffffff9000000000000000000000000000900000000000000001ffffef5c9f61b9b4f016d71060209868e4e252c13236b258025433260083834
G1[332] <= 640'h3fc00000000000000000000000000000000000000000000000000000003fffffffffffffffff80000100017007bfff1fffff3f90f5ff775ae956c103204981a38b47325030441201221fe6bc68696a
G1[333] <= 640'hfe01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7ffef7fefffffffffffd6fc1256721cf7077cc2472647666148312888051b7c001e29dde323a55
G1[334] <= 640'he1003fffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffff960d9aebb253b76f7888e7832f75d25e0986028df7f01963816f26c301d
G1[335] <= 640'h7c0041ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3ffffffffffffffffffb94ace9639402a2d2deb172d84230c6932846418bb82c004ccbfefb676fa
G1[336] <= 640'hbb8000003fff7c3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe300fe6fffffffffffff9b70fd45a487b26bf15def859fde4127b8c2461a7d98c02cf45371bc4808
G1[337] <= 640'hbbff0000007ff83fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff01fff7fffffffffffff890e513ee6d1d048c2047c4e502b874a80c608645d80c5784f53ca67dac
G1[338] <= 640'hff007fc0003ce3fcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5905f92a52b08f6718c9b74379284d0658cd220989af0c6143d2d98822fe
G1[339] <= 640'hb3c07f00083fc3fc1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcd7dff0f15b7b84be8f2db6d97422483208022c885d318012223a106089c
G1[340] <= 640'hfeffec0000cfffff0fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8db9500811293206a268c16b95f255121e238800336ac86dcff33384332d
G1[341] <= 640'h33ffe80001837eff07ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff03ffffffffff8f03f7cc8cf18d7fea7fa5613be14590d124236767a0ca059aaf6af43a53
G1[342] <= 640'h86fe60000301ffff01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fffffffffff81fffffff8fed5b6c2d09c0e8457ba70010373b048234bc3311200800008602290f1285e
G1[343] <= 640'h11ff6000000fffe1c2ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1fffffffffe3007fe0f3f00167da99a620424c847cffdf4da623904a15c218c008c1040a311121c13921
G1[344] <= 640'h5ffe000000088e000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5ffffffffc0000000000386edfc819cd374298ad1f001b770c35df03c0500cc3081690260d1f13ea190b
G1[345] <= 640'h2fff0000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4dfffffffc00ff01ffc0006fa67b215a6c2fccfa6aeaae2af3e0511ab87091218010560e2716db843740
G1[346] <= 640'hfff0000000000000ffffffffffffffffffffffffffffffffffffffffffffffffa7fffffffe6df9dffbf9ffff81ffffffcf0efda378a25549eb367752e0c6509e46a87198002848831589c48ec40f75
G1[347] <= 640'h2e360000000000000fffffffffffffffffffffffffffffffffffffffffffffffb41bffbfffdaf86390000ffffe0ffffffff26181847aab0c8a96f97328c9b4ea4a0aa30829438e01309802000063067
G1[348] <= 640'hc3000000000000007fffffffffffffffffffffffffffffffffffffff8000fff80970e0fffff27ffebf00c1fff83fffeff914d7136132fb134c85e60c4ee70104d44100c00c00422100c61031122c02
G1[349] <= 640'h2fe3f98000000000003fffffffffffffffffffffffffffffffffffc00739e03e075df0307158dfff6bbfffffffc000640030f00029c5f6253e210b3668992766e00c040c8580d3b1100a06046421b22
G1[350] <= 640'h9fffffcc080000000003ffffffffffffffffffffffffffffffffffc01fffff81c6c7de0800c9ffffdb9ffffffff8ff00001850413de2f7ebaac89c9868c17737a59680840100d186008100217000a20
G1[351] <= 640'hfffffdc0380000000003ffffffffffffffffffffffffffffffffffc003fffffbb6abbfe060f19fff4b9ffffffff9bfc30019b0e0330a9b499e825642260d1d359082e28830041a4740100242b661a10
G1[352] <= 640'hafffffcc000000000007399ffffffffffffffffffffffffffffffff0001fffde55c0b9d560f3940c6fbffffffff81e07003c9625140eeaafb39e5f6bc739cef20479de086182250528000251d165caf
G1[353] <= 640'h3ffffffc00000000000000f7efffffffeffffffffffffffffffffff8000067ff97ddf004083d9000aec407ffff9c1f1fffa73c9e3d464da9a5bb8149d9d4c99093691c8040138862041c12459241830
G1[354] <= 640'h3ffffefff00000000010c001efe7fffffffffffffffffffffffffff0000000e8cb16c499087b04fbff71600036001f9fff891487172ae09dafee889c86ef35ad123487c0604c56256c2810449880d19
G1[355] <= 640'h3ffffffffff3803400000000707f0003efffffffffffffc1ffff003000000049d75851192e6a21faa813f0000000ffffff09f58d0b94cc5715c6ce22991d1b2006404d4420012c0004298060ab400af
G1[356] <= 640'h3ffffffffffcc00040000000080007fc7fffffffffffff000000000000000008445ce730264f003c2c064000006fffffff006b5c3165b528bf7381bd90bead6501d28580102180c0303300053002100
G1[357] <= 640'h3ffffffffffce00000000000000387f3c7f0000fffffffec0000000000000034651355504a9c1cfc6c8cdc00007fffffff9a62c9073edefa100ecb7411ef438183ab9e200034818610320063944010c
G1[358] <= 640'h3ffffffffffcffc00800000000300006e001ffe0fffffffe9c00000000000023e1e544a0182338f9684cdffff19fffffff854dd3d2764eef1bcac48ac3902350127c48c02006644300010026c040180
G1[359] <= 640'h3fffffffffffffefbffe6400199afffe0f801ffc0dfffff4000000000000002405e145e93b782078fa4dffffff3fffffffb26eb26e50150b19ace24a1d19a0c431608c30000361008b0110002403c00
G1[360] <= 640'h3f81fffffffffffffe3ffff1f7fff5fbfffffff00f4f9c01000000000007c073e69a0ca50bc524783f57fffffedffffffe409658ceb016d81b27d51b07b9aab1083980c00003000c810000000521800
G1[361] <= 640'h2c2c3b7ffffffffffffffe2fffffff03ffffff8000008f0000000000018f0015b54650a348ac71f25b2fdffffefffffffef79a98c14a29d10ddbdb558a2641f901a2400006000084c30040009026400
G1[362] <= 640'h71001ef1fffffffffffffffffffffef5ffffff0107e800000000000007e7002a4fd0ebca09bd5c718fa7dffffbeffffff3d931fd8be3480518fdd2674c8a00b7310000000300400c800048413020000
G1[363] <= 640'h100001bffffffffffffffffffffff401dffffc7fff001000000002460070c220728bb54620ec8dfc22adfffff84ffffffc69af0dc70e2a8a29d6765804345744000004800100409e400000000241200
G1[364] <= 640'h70003257fffffffffffffffffffffc017ffffffe000000000000004e007001d2bdda8d7b057f75e9777dbffff867fffffe6cc6074cddc1321f35f90e9f20fa2c0000000801006008000008018440000
G1[365] <= 640'h100000dffffffffffffffffffffffc017fffffffc00000000000041f01f005ecb8c4926f80b5646beb6fbffff54dfffffccf35754ca72a808f6b83b2d1046c661500004c01003007000000000000000
G1[366] <= 640'ha00000603ffffffffffffffffffffd05ffffffffeffffc0000000486000203e8f1bb10e8d0fc1243f74efffff34bbffffffbd6001da703f0d6218b4a9a64291e0000000000020001020000040000200
G1[367] <= 640'h18000001c807ffffffffffffffffffd057ffffffffffffffc180005e4000ef8e588eaa42ef8d7f7ca3e5cbffff2e33ffffe6a1ab28d053ad4997f01dc8c3050a8080000020402c800120000000061000
G1[368] <= 640'h2519fffffffffffffffffd05ffffffffffffffffcc000cb28025afd937dbf8748597dcbd284f2ffff1a77ffb7b0efd31d00c998471cf503e0dab397a0c00d81404400004400000000041040
G1[369] <= 640'h663ffffffffffffffff405fffffffffffffffffc001dfa0a38dbd1447dd94779108a6e66b8ffffe321ffff7b4f55043935a0033d21eebe9e752da90400004e00000000000000000823800
G1[370] <= 640'h81fbddfffffffffffd06effffffffffffffffc003e380a083944f0bdf2411890ec66619e3fff8e137ffffd58e08d315a811d1dca6857085214900001404400000000800000000002000
G1[371] <= 640'hc0005e07fffffffffffff4013ff7fffffffffffffe00395d06096084d9b70adfa0a8cc5a325abfff9341fbfbff1e66cc014242298cf2027c9605c0200011cec300000003a04000000060000
G1[372] <= 640'h300e7fffffffff84009fffffffffffffffff002c5a0f5b37457c9deecd45ec8dfeb702bfffc3f673ca51eb7d786470472006b2e6699249804a00100c8000000006210000000040000
G1[373] <= 640'h1e000001111ffffffffef80023fffff87ffffffe3c0049980379450706095a17a104cedad67a8fffebfe662a1d8a38cd48d087f30aaaa39b98d4027e0006090000000000406000000000000
G1[374] <= 640'h3e0000000439ffffffe000007ffffffff8ffffc0003ca09837588c128d1c10d80bc97885cbd3ffff9c6dfdd78940aac52f00a71185ca2e5081e00060000000800000002007000000600000
G1[375] <= 640'h7fc000002c63fffffe000007fffffffffff80000078429bbb0048002df2c8cd92cd21627cef7fe79dd9fc86b0885a4403a9f9fa874ade7a8434049000002060000010000002000000000d
G1[376] <= 640'h187f000001013ffffe000007ffffff9ff817ee000f95618e70040032ea44523c18e9f467e4dffffeabff3bea30046404b843c6148f6f2bbe468000000388cb00000500000000000000008
G1[377] <= 640'h800fe000000623ffe800017ffffffffc003e019f01d9efd0b0a462013e9f8081873da73a4ffff3e7f3fa0da0e02700477a1648b4b0d22a06000180000c88800000000000000000000000
G1[378] <= 640'h80001fc00002543f680003ffffffffe0103e019fa4882b6080446104207292468db6831527fffbf2dff84f6208272044888149bc8811b024460c60008001c00000000000000000000000
G1[379] <= 640'h1ce0001fc0000141f40000fffffffe03fffffffc8d991e1a86b012448ce66d67043431c287ffec7de7f88633100280001485b82cf848194f7e1fe0000000000000000000000000000000
G1[380] <= 640'h33b80011f000004880000fffffffc07fffffffe48c166444010195000c167e54c6f3383e73ff077a5fae01180000000031581c42000a2123604c0001208000000000000000000000000
G1[381] <= 640'h1fc0001e0001000000ffffff001efffffffd8481bf000144e010c1d99607287f9a5c033ff83ee4a1ec8180000000000040228cd8ca2b0d04c2004400000000000000000000000000
G1[382] <= 640'h19003e0000e000000000783fff3f3ffffffffd4cf1981006845835ad1e08828068801cfe7ffdd56480b4000000000000000131d6f040611c0480200000000000000000000000000000
G1[383] <= 640'hc80004c400178000001301f7f7fffffef7ffcc6f0b800209618305e0792a0c27981900f5ffbda7eff608000000000000000909ee05024020080000000000000000000000000000000
G1[384] <= 640'hf000003860000000019487ffffffffefff76f88080620c9b0b8614bf54e106308189063ffbf81752700000000000000000517ce9900c000000000000000000000000000000000000
G1[385] <= 640'h306f8000000600fe0000011bffffffffffeca7c48a4f106445382274e0ce00020001804bbdbf61e7a0000000000000000002a9a9a8022120620000000000000000000000000000000
G1[386] <= 640'hf00ff8000000f000000004fdfffffffffffa7008c6140258db0322182160202000103322db8b120100000000000000000000000042604d0360000000000000000000000000000000
G1[387] <= 640'h3800fff0800003818980011fffffffffff17f508f01080718226036643042000000607242b4006028000000000000000000000000160000200000000000000000000000000000000
G1[388] <= 640'hfc0001cffff0018f89c484dffffffffe07006987014027940b001e426240580820c00023ae31b890000000000000000000000000000000200000000000000000000000000000000
G1[389] <= 640'h6fc00000003f80f00000013ffffffff0f80008010200119b19153280004040000081068c95b82500000000000000000000000000000000000000000000000000000000000000000
G1[390] <= 640'h30fff00000007c002604404ffffff002000000000002cbf949c4e3800000000000678ec173d50000000000000000000000000000000000000000000000000000000000000000000
G1[391] <= 640'h1c00ffecf80001f800090003ffffc030000000000000a151972622000000000000441cc1a0300000000000000000000000000000000000000000000000000000000000000000000
G1[392] <= 640'h7c00fcfe3f3f0007e0000048bffc000000000000000016002008e02000000000004000000000000000000000000000000000000000000000000000000000000000000000000000
G1[393] <= 640'hf8001000000f8000480002532200000000000000000009ec074940000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[394] <= 640'h1f80000000003f80003800437ff0000000000000000003f202c1c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[395] <= 640'hffc8000000007fc000f000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[396] <= 640'h3ffe780fff00071800900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[397] <= 640'h3c073ffbfc8ff8001fc0410000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[398] <= 640'hfc0010000001ff80013908010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[399] <= 640'h1f800000000011fdf00641800000000000000000001900000000000000000000000000000000000000000000000000003000000000000000000000000000000000000000000
G1[400] <= 640'hfffbe00103700083e0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[401] <= 640'h33ffff001ffe800007800000000000000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[402] <= 640'h300ffffffffffe00001f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[403] <= 640'hf0003fff8001fffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[404] <= 640'h3f000000000000fffe00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[405] <= 640'hffff800000000000ff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[406] <= 640'h1fffff07ffffc00002f800800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[407] <= 640'h3ffffffff7ffff9000030200000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[408] <= 640'h7ffffffcf0fffdf0000040000000000000000000000000000000000000000000000000000000000000000000000000001900000000000000000000000000000000000
G1[409] <= 640'hc001f000800007ffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[410] <= 640'h380000008020000000f841c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[411] <= 640'h1ffe87f87ffff0700000706000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[412] <= 640'h7fffffeffffffffff00000c18000000007800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[413] <= 640'h1e7ffffffff7fffffff880c00000000001e00600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[414] <= 640'h203bffe3000006801ffef3000000000002c0080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[415] <= 640'h3c000000000000000004c060000000000090000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[416] <= 640'hfeff9ee7ffffffce08c0018282000000034000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[417] <= 640'h3fffffff7fffffffffeff6e78000000000c800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[418] <= 640'h7fffffffffff837ffff9c7780000000003600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[419] <= 640'hfffffc0010000730000080000000000ec0180000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000
G1[420] <= 640'h1800f3fffe73ff667800000000001b0060000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[421] <= 640'h7f301f01fffffffffffff68000000000007e01c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[422] <= 640'h1ffffffff3fffffffff99ef000000000001f806000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[423] <= 640'h7fffffffffef811e3874eac000000000003f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[424] <= 640'h1effc63ffc00fefffefff87000000000000fc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[425] <= 640'h10f80fc837ffffffffffffc000000000003f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[426] <= 640'h771fff3ffffffffffffdf00000000000076000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[427] <= 640'h7ffffffffffff878fffffffff0000000001f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[428] <= 640'h3fffffffffe03ffffffffffffffff8000004000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[429] <= 640'hffffc0f7f003ffffffffff0ffffe0ff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[430] <= 640'h1001c0000fffffffffede7f7fffffc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[431] <= 640'h7fffffffffc00187fffe1fff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[432] <= 640'h3fffffffffff00007ffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[433] <= 640'hfffffffffc001077fffff780000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[434] <= 640'h3ffffc37c00f3fffffff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[435] <= 640'h37e000000fffffe77800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[436] <= 640'h1ec73ffffc800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[437] <= 640'hffffffcf00000000000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000
G1[438] <= 640'h1c3ffffff8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[439] <= 640'hfffee3000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[440] <= 640'h3e3000000000000000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[441] <= 640'hf00000000000000000000000000000000c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[442] <= 640'h30000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G1[443] <= 640'h0
G1[444] <= 640'h0
G1[445] <= 640'h4000000000000000000000000000000000
G1[446] <= 640'hc000000000000000000000000000000000
G1[447] <= 640'h0
G1[448] <= 640'h7f83c0000000000000000000000000000000000
G1[449] <= 640'h180000000000000000000000000000000602600000000000000000000000000000000000
G1[450] <= 640'h80000000000000000000000000000000103c00000000000000000000000000000000000
G1[451] <= 640'h80000000000000000000000000000000000000000000000000
G1[452] <= 640'h180000000000000000000000000000000000000000000000000000000000000
G1[453] <= 640'hc000080000000000000000000000000000000000000000000000000000000000000
G1[454] <= 640'h180000000000000000c000000000000000000000000000000000000000000000000
G1[455] <= 640'hf0000000300effffcf000000000000000000000000000000000000000000000000
G1[456] <= 640'h1c000038f3c0020040000000000000000000000000000000000000000000000000
G1[457] <= 640'h1000003cfffe00103700000a5000000000000000000000000000000000000000000000000
G1[458] <= 640'h6000300c00000000000000000000780000000003c0000a5800000000000000000000000000000000000000000000000
G1[459] <= 640'h9f30064800000000000000000000000000000000000000000000000
G1[460] <= 640'h3fffc64800000000000000000000000000000000000000000000000
G1[461] <= 640'h8000efffe5800000000000000000000000000000000000000000000000
G1[462] <= 640'hff8002fffff7eb6000000000000000000000000000000000000000000000
G1[463] <= 640'h1000000000000000000000000018c0001effff7ef7f00000000000000000000000000000000000000000000
G1[464] <= 640'h24008000000000000000000000000000000000200000007ffff7eb7f80000000000000000000000000000000000000000000
G1[465] <= 640'h7ffe3ef3fe0000000000000000000000000000000000000000000
G1[466] <= 640'hfff3ee1fee000000000000000000000000000000000000000000
G1[467] <= 640'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000
G1[468] <= 640'h4000100000000000000000000000000000000000000000040000000000000000000000000000000000000007f9deb3e7c00000000000000000000000000000000000000000
G1[469] <= 640'h464040000000000000000000000000000000000000000000700000000000000000000000000000000000000001dd73ffff80000000000000000000000000c00800000000000
G1[470] <= 640'h6660000000000000000000000000000000000000000000000cc00000000000000000000000000000000000000000099dfffc000000000000000000000007f800000000000000
G1[471] <= 640'h666000000000000000000000000000000000000000000000013c0000000000000000000000000000000000000000001fffff00000000000000000000003f71f0300000200000
G1[472] <= 640'h2400000000000000000000000000000000000000000000000184000000000000000000000000000000000000000000003fff000000180000000000408fffb0f17c0026000000
G1[473] <= 640'h3800000000600000000000000000000000000000000000000000000000010000000000000000000000007f8000000000000000000000ff810000006000000007f38e788000800010000000
G1[474] <= 640'h860000000000600000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000180000000000000000ef00c013000000000000000
G1[475] <= 640'h10004000000c001660000000000000000000000000000000000000000000000003800000000000000000000010000000000000000000000000000c000000000ff3ffff007ffe000100000000000
G1[476] <= 640'h380000020000030280cc00000000000000000000000000000000000000000000000008000000800000000000000000000000000000000000000000000000000007f3bff1168fc000040e0000000000
G1[477] <= 640'h20c00031f8900000000000000000000000000000000000000000000200000001c0001f0000000000000000000000000000000000000000000000000e13f8f9208fec000b0004400c0000000
G1[478] <= 640'h220e008380000000000000000000000000000000000000000000000020000000000001800000000000000000000000000000000000000000000000000125f8801ff0003c000000004f040004
G1[479] <= 640'he00000042207000300000100000000000000000000000000000000000000000000000000000001800000000000000000000000000000000000000000000000000000000ff000090000000000000e0400
end
always @(posedge vga_clk) begin
G2[0] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff0f733f1f783f11ff7effffff7ffffffffffffffffff7fffffeffffdfffffffffffffffffffff9ffffffffffffffcffffff7fe0fc8000
G2[1] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffdff0073cf0f3e7919fffffffffffffffffffffffffffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffff070f0100
G2[2] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffcffe033c3031ffc9cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffffffffffffffffffcff0870300
G2[3] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffec3fff03fc300ff8e9dfffffffffefffffffeffffffffffffffffffffffffffffffffffffffffffff7efffffffffffffffffffefedbe18700
G2[4] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffec3ffff1ffc00ffcf9bfffffffffeffffff7effffffffffffffffffffffffffffffffffffffffffff7efffffffffffffffffffe7f1ffcfbe0
G2[5] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffcffff8f7ffcffff93fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3993ef8e0
G2[6] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffdffff8efffcfef3dfffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffff7f81f7820
G2[7] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffff8ecfff3f37deffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7ffffffffffffffffffc9fe10f03
G2[8] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffff8ffe73f000ffffcfffffffffffffffffffffffffffffffffffffefffefffffffffffffffff9fffffffffffffffffffffeffeefcff76c3c0
G2[9] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffeffe7ff0073fffffffefffffffffffffffffffffffffffffffffefffffffffffffffffffffffffffffffffffffffffffffffefffe7ec7c0
G2[10] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffceffffceff737f1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7eff80
G2[11] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffcfffffceff7b3f3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefe9c
G2[12] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7c0fffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffff7ffffefe1c
G2[13] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1e1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc
G2[14] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffff7fffff7f803fffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffdc
G2[15] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffff7fffff7f8073feffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffefffefbf7cc
G2[16] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffff9fffefff7ff9ffcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8f77f
G2[17] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffe7f7ffefffbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3ff7ff
G2[18] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffcffe7ffeffdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8ff
G2[19] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffcfff7fc3ffbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef8f1
G2[20] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffee777e3ff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffff8ffcf1
G2[21] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffef7f77c7fdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffcffeff
G2[22] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7fff
G2[23] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff7fffe7fffdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffff7f3f3f
G2[24] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc
G2[25] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[26] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffb7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf
G2[27] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[28] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[29] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[30] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[31] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7e
G2[32] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffff
G2[33] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[34] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[35] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[36] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[37] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[38] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[39] <= 640'hffffffffffffffffffff7effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[40] <= 640'hfffffffffffffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff
G2[41] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[42] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[43] <= 640'hffffffffffffffffffffbffefeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[44] <= 640'hfffffffffffffffffffffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[45] <= 640'hffffffffffffffffffffffffe7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fff
G2[46] <= 640'hffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[47] <= 640'hfffffffffffffffffff7ffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffff
G2[48] <= 640'hfffffffffffffffffff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[49] <= 640'hffffffffffffffffffbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[50] <= 640'hffffffffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[51] <= 640'hffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f
G2[52] <= 640'hfffffffffffffffffff7ffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f
G2[53] <= 640'hffffffffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[54] <= 640'hffffffffffffffffffbedffffeffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[55] <= 640'hffffffffffffffffffe6dfeffefedf7ffffffffffffffffffffffffffffffffffffffefffffff9ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[56] <= 640'hffffffffffffffff7ffbff3ceefe7fcfffffffffffffffffffffffffffffffffffffffff738f7fefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[57] <= 640'hffffffffffffffff7ff8ffff7fe7feffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[58] <= 640'hfffffffffffffffffeffffefffe7defbffffffffffffffffffffffffffffffffffffffe7feff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb
G2[59] <= 640'hfffffffffffffffffe9fefdff3ffc47bfffffffffffffffffffffffffffffffffffffffe7cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb
G2[60] <= 640'hfffffffffffffffffefcffffe7ff711f07fffffffffffffffffffffffffffffffffffffedffffd9ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[61] <= 640'hfffffffffffffffffffdffff7fff739fffffffffffffffffffffffffffffffffffffffe7dffffd9ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe
G2[62] <= 640'hffffffffffffffffff1fffe7fcfff3fcff99ffffffffffffffffffffffffffffffffffffffffcddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[63] <= 640'hffffffffffffffff39f9ff3fff7ce0ff67997b77feffffffff7ffffffffffffffffffffffcfccd81ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[64] <= 640'hfffffffffffffffffff10737fff321f99cff9ffffffffffffffffffffffffffffffff7ff4dffff8fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[65] <= 640'hfffffffffffffffffff13f70fff3615999ffbfeeffffffffffffffffffffffffffffffffecfcfffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[66] <= 640'hffffffffffffffffff7bf870ff73f04939f07fe6ffffffffffffffffffffffffffffffffed3ffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[67] <= 640'hffffffffffffffffe03fc326c7e0ccc139fb7ffffffffffffffffffffffffffffffffbffef3fcf1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[68] <= 640'hffffffffffffffffff0f0f0ec71f8ec10c7f67fffffffffffffffffffffffffffffffbfff8f8cff9ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf
G2[69] <= 640'hffffffffffffffffff8e3c6ecf0f8e0c0437277ffffffffffffffffffffffffffffffbfff9f0cfd1fffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[70] <= 640'hffffffffffffffffffcc3cc60f1e804c04010f7ffffffffffffffffffffffffffefeffff6f3fcf9bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[71] <= 640'hffffffffffffffffffccc3860ffcc0c720f019ffffffffffffffffffffffffff7ffef2ff69fe8719ffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7b
G2[72] <= 640'hffffffffffffffff7f3e993107ffe4c3638c0efffbffffffffffffffffffffffff7fffdfe0ef2107ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[73] <= 640'hfffffffffffffffff0f88100803e0eff780006ff7fffffffffffffffffffffffffffcfffffcf87f1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[74] <= 640'hfffffffffffffffff3f88100801efcff7e008b737ffffffffffffffffffffffffeefef7ffffece3fffffffffffffffffffdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[75] <= 640'hffffffffffffffff3f9f0000001ef43fcf011b63ffffffffffffffffffffffffffffff7ffefece3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[76] <= 640'hfffffffffffffffff89c2000000f0707c400198ffffffffffffffffffffffffffffffffeffffcef9fffffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[77] <= 640'hffffffffffffffffe398c000000002cfbc00008ffffffffffffffffffffffffffffff9ffffffc03bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[78] <= 640'hffffffffffffffffc39800000000603e1e00303f7ffffffffffffffffffffffffffff03fffffc01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[79] <= 640'hfffffffffffffffffd813e0000086038c0007e7ff3fffffffffffffffffedefffffef0f8fef3e0303fff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[80] <= 640'hfffffffffffffffffc98000020010600180007efefbf7fffffffffffffffffffffefcf7ffefff040fffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffff
G2[81] <= 640'hffffffffffffffffc79d0000000080000000017e66ffffffffffffffffffffffffeff07fffffe000ffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffff
G2[82] <= 640'hffffffffffffff7ee78f00000000c0808000003f70ffffffffffffffffffffffff7fffffffffc0001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
G2[83] <= 640'hfffffffffffffffffc0f0000800001808000000371ffffffffffffffffffffffff7f7fbffffcc00000fffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffff
G2[84] <= 640'hffffffffffffffef3e3c0000000001800000000163fffffffffffffffffffffffffff8bffffc80001f7fffffffffffffffffffffffffffffffffe7ffffffffffffffffffffffffffffffffffffffffff
G2[85] <= 640'hffffffffffffffffc230c0000000000000000018637fffffffffffffffffff7ffffdfdffffc300000f7fffffffffffffffffffffffffffffffff3f8fffffffffffffff7fffffffffffffffffffffffff
G2[86] <= 640'hffffffffffffffffe020c000000000000000000c00671fffffffffffffff9ffffffdffffffc00000007fffffffffffffffffffffffffffffffff3cfcffffffffffffff7fffffffffffffffffffffffff
G2[87] <= 640'hffffffffffffffff7e030000000000800000008704661b3fffffffffffffcffefefdff7ffffc000000bbfffffffffffffffffffffffffffffffee3ffffffffffffffefffffffffffffffffffffffffff
G2[88] <= 640'hffffffffffffffff001100000000100000000000818efc7fffffffffffffe7fffffef8fff3e00000033f7ffffffffffffffffffffffffffffffee78ffffffffffffff1e3ffffffffffffffffffffffff
G2[89] <= 640'hffffffffffffffffe01000000000000000000000890c3ffffffffffffffffbff3cfeff0fb6c00000103ffefffffffffffffffffffffffffffffff0c63fffffffffffe3ffffffffffffffffffffffffff
G2[90] <= 640'hfffffffffffffffefc080000000000000000000081007effffffffffffff1fffffffff0f96c00000083fffffff3fffe3ffffffffffffffffffff7c803fffffffffffff3cffffffffffffffffffffffff
G2[91] <= 640'hfffffffffffffffefc0c0000000000000000000000007e7ffffffffffffe1fffe3ffff0f92800000071e9f7ee01fffc03fffffffffffffffffffc700ffffffff7fff3e3cff7fffffffffffffffffffff
G2[92] <= 640'hfffffffffffffeffcc0c0000000000000000000000010f7fffffffffffff99ffefffff07b3000000000efdfff01fffcc1ffffffeffffffffffffc0000fffffffffff1eff7f7fffffffffffffffffffff
G2[93] <= 640'hffffffffffffffffcc800000000000000000000000017ffffffffffffffec0ffffffff0733800000000effe7f01cffd883ffffffffffffffffff880007ffffffc7ffc3ff3ff9ffffffffffffffffffff
G2[94] <= 640'hffffffffffffffffcc40000000000000000000000000fffffffffffffffe67cf3cf8ffff32c0000000000fff0000ff0001ffffffffffffffffff9c0003ffffff87ffcf6083f1ffffffffffffffffffff
G2[95] <= 640'hfffffffffffffff0cc00000000000000000000000018ffffffffffffffffe6effff83fce12c00000000166ff1c00c00100fffffffffffffffffff80000fffffffce3fe7183f33fefffffffffffffffff
G2[96] <= 640'hfefffffffffffffc70000000000000000000000000337fffffffffffffffc0889ff38f790081600000034d389901000080fffffffffffffffffe4000013fffffefff7f0030f3e7fffeffffffffffffff
G2[97] <= 640'hfffffffffffffffff0000030080000000000000000b3ffffffffffffffff07c78f7087398181000000004101f800000001ffffffffffffffffff4600033fffffffffff0000ffe6ffffffffffffffffff
G2[98] <= 640'hfffffffffffffff3f0000078ff80000000c0000000b3feffffffffffffff07cf9f00011f83800000000000016000000001fffffffffffffffffe06f0069ffffffffffc008c7ffeffffffffffffffffff
G2[99] <= 640'hfffffffffffffff3f100007fffc000000330000000b3ffffffffffffffffc0cf1c00008f180000000001000006000000003ffffffffffffffffe0698069ffffffffffc00803f3d7fffffffffffffffff
G2[100] <= 640'hfffffffffffffff90f0000ffff700000033800000032ffffffffffffffff06f81800008e180000000000000006000000001ffffffffffffffffe00904099feffc7fffc000038397fffffffffffffffff
G2[101] <= 640'hfffffffffffffff81e0000fffe30001007fc000000163fffffffffffffffc01080000007010000000000000000000000000ffffffffffffffffe90800018defd1cc31e000038337fffffffffffffffff
G2[102] <= 640'hfffffffffffffff9180001fffff000187ffc000000073bffffffffffffffe000000000000100000000000000000000000007fffffffffffffffff8008000ffd918c000000000636fffffffffffffffff
G2[103] <= 640'hfffffffffffffef1380001ffffe0000cff78000000077bfffffffffffffd0600080000001800000000000000000000000003fffffffffffffffffc600001ff19800000000000666fffffffffffffffff
G2[104] <= 640'hffffffffffff9f70800001fffff8000ccfd8000000037ffffffffffffff8000800000001000000000000000000000c010003fffffffffffffffffc00000046e000000080000cf1cfffffffffffffffff
G2[105] <= 640'hffffffffffffff20800001ffffe0000ceffc0000000cfffffffffffffff9000000000000000000000000000000000c000003fffffffffffffffffe00000027000000000003007fefffffffffffffffff
G2[106] <= 640'hffffffffffffee60b080037fffe000017ffe0000000cfeffffffffffffff01000000000000000000000000000000388000037ffffffffffffffffe000000030c0000000003000fffffffffffffffffff
G2[107] <= 640'hffffffffffffee803000037fffe00001ffee00000001fffffffffffffff8000000000000000000000000c000000019e600017ffffffffffffffffe80008000000000000000e30fffffffffffffffffff
G2[108] <= 640'hffffffffffff7e003200037ffff00000fffe00000001773ffffffffffff800000000000000000000000fe000000019e360007ffffffffffffffffe80000000000000000000c387ffffffffffffffffff
G2[109] <= 640'hfffffffffffffe803200013ffffc0004ffffc08000002307ffffffffffe000000000000000000000001ce00010019df13c007ffffffffffffffffe0000000000000000000083c3ffffffffffffffffff
G2[110] <= 640'hffffffff7fffcc800200013ffffc000cffffc38000000077ffffffffffe00000000000000000000001fcf8001003b9990e007ffffffffffffffffe0000000000000000000001ffffffffffffffffffff
G2[111] <= 640'hffffffffcfffc8800200010f77c0811fffff0f8000008063ffffffffffe00000000000000000000001effc80023ff9dfeee0077efffffffffffff08000000000000000000103fffeffffffffffffffff
G2[112] <= 640'hffffff79fffff800100000107fc0807efffffe6000000103f7ffffdffff000000000000000000c0007efe3008170f9f7f3807bfffffffffffffff1000000000000001801001fffffffffffffffffffff
G2[113] <= 640'hfffffffefffff800000000003fc0080efffffee40000000bffffffffffc000000000000000010c0207effc00003fffffb200317ffffffffffffff000000000000000000003ffffffffffffffffffffff
G2[114] <= 640'hffffffcefbfff000040000003f81000fffffffc4000000199fffffffffc00000000180017ff88e0707fffc001c1fffffbe00000ffffffffffffff800000000000000001813ffffffffffffffffffffff
G2[115] <= 640'hffffffceffffc00006000000ff000001fffffffe010000189fffff7fffe0000007138e31fffc8f0317fffc1c1ffffffffa0080027ffffffffffffc00000000000000001cfbffffffffffffffffffffff
G2[116] <= 640'hfffffffcffffc00004000000cf000001fffffffe80c00001bfffffffffe0000000fb1f39ffffff80b6ffd9fe7ffffffff0808000fffffffffffffc000000000000000013ffffffffffffffffffffffff
G2[117] <= 640'hffffff78cfffc0000000000080800000fffffffc80400001ffff7ffffff000010c993019fffffefc1ffffc3ffffffffff0808000fffffffffffffc000000000001000023ffffffffffffffffffffffff
G2[118] <= 640'hfeffff210fffc0000000000280000000cfffffff02000001fefffffffff800000f9d0c1fffffffff1ffffc1fffffff9ff00000013ffffffffffffc000000000000000107ffffffffffffffffffffffff
G2[119] <= 640'hfffffc013fffc00000000003cc0c00000fffffffe00000006efffffffff800001f9f0c8fffffffffbffffd3ffffffff080000001fffffffffffff8c6000000000000000f7fffffffffffffffffffffff
G2[120] <= 640'hfffffe600f7fc000000000021c0600004fffffffe8000000fffeffffffe000019f7f02fcffffffffff7fff3ffffffff0c000000037ffffffffffff0fc00000000000041fffffffffffffffffffffffff
G2[121] <= 640'h7eff7e0006ff81020000001003001800efffe0fffe0000033fffffff7ff000031f01100ffffffffffffff87ffffffff80000000037fffffffffffcfff40000000000021fffffffffffffffffffffffff
G2[122] <= 640'hff7ffe0006ff98300c000010030c9c000ffc00302ec000003ffffefffefc00071f433003ffffffffffe7fc7ffffffff80400000013fffffffffffcfffc1c00800000037fffffffffffffffffffffffff
G2[123] <= 640'hff7ff30007ff8000000000123880c0000fdc0420000003c03f7ffefffffc00061fe316f7ffffffffffffff3fffffffe80000000013ffffffffffffffff3e0000000003ffffffffffffffffffffffffff
G2[124] <= 640'hc6ff078007ff80800000000339c007f0ff0f40000000037ffffffffffffe00009f703f7fffffffffffffffffffffffe80040000001bfffffffffffffffff000000000cffffffffffffffffffffffffff
G2[125] <= 640'h3efe3f2002ffc0000100000293e17ff807c6010000031e7ffffffffffffe00008378ffffffc7dfffffe3ffffffffffec000000000017fffffffffffffff9e0c000000fffffffffffffffffffffffffff
G2[126] <= 640'h7ffc782002ffe0000000000091e07c7f07f4898000000cffffffffffffff800003ffffffee011ffffff3ffffffffffff000c00000017fefffffffffffff9eec000009fffffffffffffffffffffffffff
G2[127] <= 640'hf1f0072007fc00300000000010000601823e89f0000083f7ffffffffffff8000037f3fffee001fffff7fffffffffffff0048000080103effffffffffffffffc00000bfffffffffffffffffffffffffff
G2[128] <= 640'h38660461011bc904000000000000080e231f0ee0b000337ffffffffffffe8000661ffffecc003ffffffffffffffff7ff0080000130061bff97fffffffffffbf880063fffffffffffffffffffffffffff
G2[129] <= 640'he30006e040b3d8000000000000000046469e3fe7100000e7ffffffffffff8000071ffffff0000fffffffffffffffff7ff1000003300099fffffffffffffffff8c00fffffffffffffffffffffffffffff
G2[130] <= 640'hc00060800d63580100000000000001648e0e3ffff00000e7ffffffffffff8000f81fffff70000ffffffffffffffffffff80001c7780003fffffffffffffffffe87ffffffffffffffffffffffffffffff
G2[131] <= 640'h567e90000000000000001efccc611fff000013fffffffffffff800899ffffff700007fffffffffffffffbfff88001e7ff80031bbfffffffffffffff02ffffffffffffffffffffffffffffff
G2[132] <= 640'h7ef900000000000000037ffce48150960001fcfffffffffff9800c1fffff7ecc0007fffffffffffffffbfff8c03be7ff40001933ff7fffffffffffff7fffffffffffffffffffffffffffff
G2[133] <= 640'h7e7800000000000000057ff97e8710060003f1ffffff7ffff9000cfffffd7fcc0017fffffffffffffffffff3303fffffc1000023ff7fffffffffffffffffffffffffffffffffffffffffff
G2[134] <= 640'h9d78000000000000000c4fff7f0618c0000703ffffffffff7900cffffffdffe0001ffffffffffffffffffff371fffffff0e00003ffffffffffffffffffffffffffffffffffffffffffffff
G2[135] <= 640'h8b60000000000000000d4fffff7effe2820010ffffffffff3901effffffffff1001ffffffffffebffffffff8c3ffffffffff00023e7edffffffffffffffffffffffffffff7ffffffffffff
G2[136] <= 640'h24800000000000000006dffffffeffffc00112dfffee1e8f8803fffffffffff8007ffffffff7fdfffffffff13fffffffffffe600318efffffffffffdffffffffbfffffffffffffffffffff
G2[137] <= 640'h6800000000000000007bfffffeffffec0000207ffee8fc180003ffffffffff88c7ffffffffffdfffffffff91ffffffffffffe0000c08fffffffffffffffffffffffffffffffffffffffff
G2[138] <= 640'h20000006008000000000000003fffffffffffe58000003ff04017000017ffffffffefc8cfffffffffffdbffffffffc1fffffffffffff0000000fffffffffffffffffffffffffdfffffffffffffff
G2[139] <= 640'h100000000000000000000000003fffffffffffec88000213b1100380001fffffffffffe99ffff7f1fffec3fffffff78fffffffffffff8000000073fffffffffffffffffffffffffffffffffffffff
G2[140] <= 640'h2000000000000000019fffffffffeffc9180000ff0100300009fffffffffffe9bffffffffffec7ffffffe787ffffffffffff8000000013ffffffffffffffffffffffffdffffffffffffff
G2[141] <= 640'h3ffffffffffff7d00000030008001000cffffffffffff73ff9dfffebfec7ffffffeff7fffffffffffd8200000011fffffffff7fdfffffffffffffffffffffffffff
G2[142] <= 640'h29fffffffffff7de0000000000000000cffffffffffff77ff9dffffbffc6fffffffff7ffffffffff8800000000107ffffffffffffffffffffffffffffffffffffff
G2[143] <= 640'h2110000010000000000000080049ffffffff73ff96000000060080000017ffffffff7fffffbddffffbffd67fffff3fcffffffffffe30000000000077ffffffffffffffffeffffcffeffffffffffff
G2[144] <= 640'h6800980100000000000084c0188fffffffddfefbc93000004000000010fffffffbfffffffdd6c6ffdff81fffffff0e7fffff7fffe000000000003ffffffffffffffffff9ff7ffffefeffffffffff
G2[145] <= 640'h10000000000001c00183fffffffffff7ffde0000200000000007ffffef9fffffff9f20ffffffdf1ffffffe37ffffe7fffc000000000007fffffffffffffffffff1f1ef97fffffffffffff
G2[146] <= 640'h1400000000000000000003800003fffffffffffffffe0000000000000017ffffcffffffffc1120ec13f7dc3ffffffe3fffffeffff80000000000076ffffffffffffffffffff8c983fffffffffffff
G2[147] <= 640'hc000000040000000000001000061ffffffffffffffe000000000000001ffffff7fefffffc0030080064c07fefff83ff9f6f8ffffc0000000000020fffffffffffffffffffc8c88c0dbffffffffff
G2[148] <= 640'h61ffffffffffffffc000000000000003ffffff60ce7ffbd8800000040046fef91f1fd93690ffffe00000010000017ffeffffffffffffffff708c00f9ffffffffff
G2[149] <= 640'hc000031ffffffffffffffc000000000000003fffff9201c7fff9c800000000000e7310e860122009fffe000000100000131fef7ffffffffffffff200000f17fffffffff
G2[150] <= 640'h10000000000000c000009ffffffffffffffc080000000000002fffef01f3effffdc0000000000016100008040e0001ffff00008c0000001387ffffffffffffffffc00000023ffffffffff
G2[151] <= 640'h37800831ffffffffffffdc0000000008000027ef7f7fbe7fffffc800000000001600000106420009dfff8001802000080307fffffffffffffff0c00000003ff7fffffff
G2[152] <= 640'h1822000000000010010000000030001e1fffffffffffff3000000000000006fffe78ba7ffffffe000000000000000000803300000f7fe0000100000001000ecfffffffffffffe0000000047fffffffff
G2[153] <= 640'h816000000000001000000000003e00880fffffffffffffe000000000000003997fff937fffffff00000000001000000000120000801fe00000000000000039ffffffffffffff300000000177ffffffff
G2[154] <= 640'h83008000000000100000000000700000cfffffffffffffe000000000000003107fcf97ffffffff00000000000000000000020000810e700000000000000171ffffffffffffff2000000001f7ffffffff
G2[155] <= 640'h188080000000000000000000006000008fffffffffff7e18000000000000001100fe97ffff7ffb8000000000000000000000008019007000000000000001e13fffffffffffffe000000001ffffffffff
G2[156] <= 640'h1cc080000000000000000000000600103ffffffffffd7e8800000000000000011f7fbf9fff7ff880000000000030e0000000000018002000000000000000861fffffffffffffc0000000193fffffffff
G2[157] <= 640'h198300000000000203000000000e001c3fffffffffffffc0000000000000000003f3bedf7efff880000000003e7bf80000000000800000000000000000008c3fffffffffffffc0000000193fffffffff
G2[158] <= 640'h9b27800000000003cec00000000c000c7fffffffffffffc000000000000000000083bac73efff880000000017fffff00000000004000000000000000000004ffffffffffffff0000000100ffffffffff
G2[159] <= 640'h18f0c01000000003fc180000000c000cfffffffffffffe980000000000000000010092c68c81e08000000001fffffff8000000006000000000000000000100ffffffffffffff00000000009bffffffff
G2[160] <= 640'hcf8402000000003ffe4000000872003ffffffffffffffeb200000000000000000010747f0c0e00000000003ffffffe03000000110000000000000000000006387fffffffffc00000000000fffffffff
G2[161] <= 640'h87f8000001000003fffe800000010003ffffffffffffffeaf800000000000000000000060301e00000000007ffffffe080000000000000000000000000000077e7ffffffff8e0000000008ff0fffffff
G2[162] <= 640'hc7b8000001000001ffe6800000000c07bfffffffffffffeac00000000000000000000004000080000000000ffffffff08000000080000000000300400000003effffffffffdc000000000023ffffffff
G2[163] <= 640'h6e1b4c0000000000ffc6000000000003ffffffffffffffea000000000000000000000000000000000000000fffffffb00c00000480000000000fe060000000183ffffffffffc008000000103ffffffff
G2[164] <= 640'h7e83480000000000ffc6800000000000ffffffffffffffeb7000000000000000000000200000000000000003fffffff01800000000000000001fe36c000000013fffffffff1f0000000000f11fffffff
G2[165] <= 640'h67810880010100001fff000000000000ffffffffffffffeb7000000000000000000000000400000000000001b3cffef000000000000f00000087f76c000000013fffffffff00000000000031ffffffff
G2[166] <= 640'he3900880010000003ffe0c00000000003fffffffffffffeb70020000000000000000000004000000000000009003fe600000000086fcf0080087ff6e000000011ffffffffec0000000000007f0ffffff
G2[167] <= 640'h62bfdc1c180080007ffe8000000000007effffffffff7eb9fe800000000000000000000400420000008000001000e600000001001effbec00c1fffefe20000000ffffefffe8100000000011c7fffffff
G2[168] <= 640'h9c6fe30000203003dff78000000000003fffffffffffffcff1880000000000000000100000000000000000000000000000000011ffff7ff7813bfdfe600000001dfbfffffc1800000000003e3fffffff
G2[169] <= 640'h83fdff80006000001ffef800000000003ffffffefffffecfff980000000000000080000000800000000000000000000000000011ffffffffdd3bffffe000000001fffffff800000000000001e3ffffff
G2[170] <= 640'ha3cd3fcc0c900c00fcfef800000000001efeffffffffffeffef00000000100000000020000000000000000000000000000000083ffffffffffffffffe000000003bffffbf000000000000003f3ffffff
G2[171] <= 640'h770f3cc61c988cc3f8ffc100000000003fdffffffffffffffee000000001000000000200000000000000000000000000000000fffffffffffffffefff600000001fffff900000000000000037c7fffff
G2[172] <= 640'h764fe06000bffee39fffc760000000007fdb7ffefffffbfffbf8000000000000000026000100000000000000000000000000017fffffffffffff7fffff00000001fffe9800000000000000073effffff
G2[173] <= 640'hf2fde06101bf7b39bf7ffc400000000027bd7fffe0cffffdfbe0000000000000000002000000000000000000000000000000037ffffffffffffffffffe000000001ffc88000000000000000ccfe7ffff
G2[174] <= 640'h8279e32001277b3cf97ffe400000000003bc7767c06ffffdff4000000000e000000002e0400000000000000000000000000006fffffffffffffffdfffff00000003700000000000000010000cfffffff
G2[175] <= 640'h9a61ff0c0066ffffffefffe0000000000fdc76e00777fffffee000000000000006101880000000000000000000000000800006fffffffffffffffff3dff0000000e000010000000002208303fc7fffff
G2[176] <= 640'hd831c322001feeffffffff80200000000efffe3338cdfffffdc000000000000000000606000000008000000000000080000000fffffffffffffffffe9fce000000001106011100000200000f7e7fffff
G2[177] <= 640'h1830102003ffffffffffff182000000007fffff0c04fffffff00000000000000001000e0000000000000000000000000000000ffffffffffffffffff9ffe0000000000000000000000000081f7ffffff
G2[178] <= 640'h1800004003ffffdfffffff980080000003fffff88101fff9ff0000000000000000100400000000000000000000000000000000ffffffffffffffffcf9fff000000000000000000000c000000f7ffffff
G2[179] <= 640'h8000ffffffffffffc30480000000bfffff0100e7fbf98000000010000001010c000000000000000000000000000000010ffffffffffffffff37fff00000000000000020030081000017ecfffff
G2[180] <= 640'h8000000000fffff9ffffffe76c80000100f9fffe000007fff880000000030000c40300c000000000000000000000000000000107fffffffffffffff973fb800000000000000200c000b200013fffffff
G2[181] <= 640'h81000000417ffffbfffffffffc8c000000fffffec00007fff8000000000300010460000000000000000000000000000000000007bfffffffffffffff73fbc000000000000000008001120080439fefff
G2[182] <= 640'h8000000000fffefffffffffef6f80000017ffffe800007fdf9800000000000010470b100000000000000000000000000000000009fffffffffffffffe7f380000000000000000100010200c0679fffff
G2[183] <= 640'hd000011000ffffffffffffe767e80000037ffffe800060cff3c00000000400103e66b160000000000000000004000000000000009efffffeff7bfdffe7c780003ec08ff00000013c309700997cffffff
G2[184] <= 640'hc0000000007fffff7fffffffe790000080c6fffc8000006778060000003080c0b9cc0780000000000000000000000000000001077bf7ff7fffdf7f6f601f8008fffffffc000001039866ff7338feffff
G2[185] <= 640'h3fffff7ffffffffff80300097fffff800000037d800000003b8c0791fc00800000000000000000000000000000000000f3fee3ff8fffe7e6f8004dffffffff1800010018e7c3ffb9ffffff
G2[186] <= 640'h1ffffffffffffffffe0700001fffff0000003f4fb00000063fff3381fcc1662000000000000000000000000018000000fffec1018ff7f7f600004dfffffffffc00003809c3f7cefbffffff
G2[187] <= 640'h1fffffffffffffffeec0000091fffc000000004f90000006fef9f081fb876600000000000000000000000000100000013f0c1900ff73fefe00004fffffffffff00001009f9e78ef7ffffff
G2[188] <= 640'hfffffefffffffffe6c00003f9fffc000000006190000127fff9c7f8f7ffe6c00000000000000000000000000000000003e0190000387f7c00000fffffffffffc0000011b9011f23ffffff
G2[189] <= 640'hf7effcfffffffffff98000318fffc00000006638000013fff7bcff8ffffeef80000000000000000000000000000000001c000000038df7800001dffffffffffe00001109f033f7fffffff
G2[190] <= 640'h3fc9f4fffffffffff98000018fff800000000448000001f7ffffff91ffffffc00000000000000000000000020000000000000c10010816000000dfffffffffffc000010077f7bffffffff
G2[191] <= 640'h13f9f0ffffffffffb910000c03f980800000044020004ffffff7ffb1efffff800000080000800000000000020800000000026c10091984000004dfffffffffffe8000107e3ffe67ffffff
G2[192] <= 640'hc40c07fffffffffbc08c00001ec00000000001c080007f7fff7ff8c3efffff0000800000000000000000000098000000000166800c0004000033ffffffffffe380000e0187cfffffe7ff
G2[193] <= 640'h6c547ffffffffffc48c0000000000000000000000067cfffffff801effffc00000000000000000000000031f800000000006600000000000003fffffffffff600008081fcffdfffffff
G2[194] <= 640'h4143ffffffffff8718000000000000000000000006eccffefff9003ffffc00000000003000100800000033e00000000000000000000000000273c7fffffffc000000987effffffffff
G2[195] <= 640'h37fffffffffe000000000000000000000000006c5c7fe0ffbb1bfffffc0000000027000364c00000c7fe2400000000000000000000000000101ffffffec00000081077fffffffff
G2[196] <= 640'h803ffffffe7fef000000000000000000000000003cff3ff1f7183bfffffc0000000309c0196ec00000e3f76c0000000000080000000000000001f4fffff8000000083f3fb7fffffff
G2[197] <= 640'h7fc00000000ffffffff7ff3c00000000000000000000000217c79f31800033fffff9980000012de8b9fec0010873f7e8000000000000000000000000000000dff710000000083ff7bff7fffff
G2[198] <= 640'hf00ffe000000008fffff7e7ff1c00000000000000000000000204c7cfce08019ffffff9c80000007ffffffec0000831fff80000000000000000000000000000000790000000001013f3fff7fffff
G2[199] <= 640'h201f00ffe9e000000ff9ff7fe7ef0c8000000000000000000000102c39c9cc08d99ffffffdca0000086fffffeec00009c3f9f9800000000000000000000000000000000000000001008fffbffffffff
G2[200] <= 640'h7c3fe9ffff3000000cffefff99ff3c00000000000000000000000030cc780003ff1ffffff7e00000003fffffff1000fc0fff7c60000810000000000000000000000000000000000001919fe6f7fffff
G2[201] <= 640'h3fffffffffff8000001e3ffef9190700000000000000000000000001003080000ff3ffffffffe000007ffffffffc0007c7ffff660000000000000000000000000000000000000000000f81ffffffffff
G2[202] <= 640'hffffffffffffd6910018fffb38000700000000000000000000000000003081c087ffffffffffe000007ffffffffe0007fffffffcc000000000000000000000000000000000000000000699ffffffffff
G2[203] <= 640'hfffffffffffffeff0000f0f700608000000000000000000000000000000199c007fffffffffff4061f7ffffffffe801ffffffffce00000000000000000000000000000000000000000243c0fffffffff
G2[204] <= 640'hfffffffffffffffe8006dff3c060800000000000800000000000000000809830377ffffffffffc043fffffffffff81fff97fffffc000000000000000000000000000000000000000000018cfefffffff
G2[205] <= 640'hfffffffffffffffe00070fe080000000000000000000000000000000008098003bfffffffffffe06ffffffffffffc1fff8ffffff8000000000000000000000000000000000000000000100ffecffffff
G2[206] <= 640'hfffb7fdfffffffff0000000000000000000000000000000000000000008010007fffffffffffff1ffffffffffffff3fffffffffd0000000000000000000000000000000000000000000107ffffffff7f
G2[207] <= 640'hfffc2689ffffffff80000000000000000000010c0000808080000000000000ffffffffffffffffdfffffffffffff76ffffffffff300000000000000000000000000000000000000000083eff67ffffff
G2[208] <= 640'hfff9670004ffffffc40000000000000000001827000000860000000001431f7fffffffffffffffffffffffffffffffffffffffffe00000000000000000000000800000000000000000011cbeebffffff
G2[209] <= 640'hfff97600001ff9ffe000000000000000000080008000000720000000006c1f2fffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000190fe6fbffffff
G2[210] <= 640'hffffe000000efcfff0000000000000000000022000000108f0000000007cdeffffffffffffffffffffff310380fffffffffffffffe00000000000000000000000000000000000000001807e67bffffff
G2[211] <= 640'hff7fc0000000b83ff80000000000080000000200000000fff0800000016fcffbfffffffffffffffffffe0080000ffffffffffffffc000000000000000000000000000000000000000000807eefffffff
G2[212] <= 640'hff7ee0000000001ffc0000000000811003000000000000fff000000033edffbffffffffffffffffffffe00000001ffffe3c00ffffc000000000000010000000000000000000000000001007fecffffff
G2[213] <= 640'hfffe78000000000fff0000000000c7fc03000000000083fffd00000037fc3fffffffffffffffffffffff80000000ffffe00003ffff0000000000000344000000000000000000000000000983ef7fffff
G2[214] <= 640'hfffebc0008000007ff0080000fc7effec0000000000087fffe80000077fc7fffffffffffffffffffffe100000000fffe6000001ffff8000000000003fff00000000000000000000000000383577fffff
G2[215] <= 640'hffff88003c0000007fffc0c11fff7fffff00000001001ffffe8c000177cd7fffffffffffffffffffffc000000000fffe000000007fff636000018673fff18000000000000000000000000193473fffff
G2[216] <= 640'hffffc000ff00c0017ffffff99fffffffdd0000000007ffffff33c1111fe37ffffffffffffffffffffe00000000000f00000000001fffff03000019dfffffe03000000000000000000000004c49abff5f
G2[217] <= 640'hd3ffe000fffff000ffffffffffffffffff8000000002ffffffffe011bffcfffffffffffffffffff0f80000003c000000000f70000ffffff3ff0f99fffffff7000000000000000000000000aea1ebffff
G2[218] <= 640'h807e8007fffffc000fffffffffffffffff00000000c7fffffffffc9bff7cfffffffffffffffe38c00000001cff7c0000007ffe0000ffffffffffdfffffffffc400000000000000000000008cf2ebffbf
G2[219] <= 640'h2601fffffffe0007ffffffffffffffff0000020347ffffffffffffffffffffffffffffffff30000000003fffff000003fffff8004ffffffffffffffffffff800000000000000000000025dd2eaffbf
G2[220] <= 640'h1fffffffe0001ffffffffffffffff00000207effffffffffffffff7ffffffffffffffff2000000000ffffffc023fffffffe000dfffffffffffffffffff800000000000000040000005fc26f7fef
G2[221] <= 640'h3ffffffff00003ffffffffffffffff000100fffffffffffffffffffffffffffffffffff0000000000ffffffffffffffffff00017ffffffffffffffffff3000000000000000c0000001eb6ebffeb
G2[222] <= 640'h3cfffffffff00000fffffffffffffffc0001efffffffffffffffffffffffffffffffffffe00000000003fffffffffffffffffe0017fffffffffffffffffff80000000000000040000008e8269ff7b
G2[223] <= 640'h26ffffff3fff800000ffffffffff7fff000097fffffffffffffffffffffffffffff9fffffe00000000003fffffffffffffffffe001fffffffffffffffffffc1800000000000000800000083049ffb2
G2[224] <= 640'h3bfffffc63ffe3040003fffffff3ffffc000ffffffffffffffffffffffffffcf9f0cfffffb0000000c803ffffffffffffffffff0003fffffffffffffffffffc0000000000000468290003f005f4d7c
G2[225] <= 640'h7ffffff823ffff7f8000fffffff1fffff000ffffffffffffffffffffffffffcfffc1fffffc8000003fc07ffffffffffffffffff8001fffffffffffffffffffc00000000000008097000024962b6dfc
G2[226] <= 640'h1fffffff801ffffffe0003cffff71fffff007ffffffffffffffffffffffffffcfffc13fff7c0000017fec7ffffffffffffffffffc000ffffffffffffffffffff800000000000136f600013412614f5c
G2[227] <= 640'h99fffffff0017ffffff000181cff00ffff981ffffffec3c7ffffffffffffffffcfe7c33eff3c017003ffff7ffffffffffffffffffc0007fffffffffffffffffff88000000000012b228010320000416c
G2[228] <= 640'hf87ffffff000fffffff0000000f800ffff983fffffff8103ffffffffffffffffeee7833effc0013801fffffffffffffffffffffffe0003fffffffffffffffffffcc000000000016008000138f0285369
G2[229] <= 640'h7fffffffe000fffffffb0000002000ffff89ffffffee0001ffffffffffffffffdc7f081cffc0003800ffffffffffffffffffffffff0003fffffffffffffffffffc000000000001f8214001d98b24d509
G2[230] <= 640'hfffffffd0000ffffffffc0000000003fffcfffffffe000000ef3ffffff9fb9f8fcbf00083fe0001e00ffffffffffffffffffffffff0003fffffffffffffffffffe000000000000ecaad00540034817b8
G2[231] <= 640'hffffffff00003fffffffe0000000001fffdfffffffc000000021fc00ff8319009c990001077800c703ffffffffffffffffffffffff8003ffffffffffffffffffff0000000000004943c805868240197c
G2[232] <= 640'hfffffffe80000ffffbfff00000000007ffffffffff00000000200100b8000000063801008000000fc7fffffffffffffffffffffffc0001ffffffffffffffffffffc00000000000a83e0049125061b980
G2[233] <= 640'hfffffffe00000ffff3ffff0000000007fffffffc38000000000000000000000006bc00000000003ffffffffffffffffffffffffffe0001ffffffffffffffffffff8000000000015c02c80f58401b2968
G2[234] <= 640'hfffffffe1800ffffffffff8000000001fffffffc00000000000000000000000000000000000000ffffffffffdfffffffffffffffff00007fffffffffffffffffffff0000000001baa2501f502011ab4c
G2[235] <= 640'h1ffffffc0007ffffffffffe0000000007ffffff800000000000000000000000000000000000000ffffffffffffffffffffffffffff00007ffffffffffffffffffffc00000000803690800d1d1b7aaa00
G2[236] <= 640'h7fffffe830fc17ffffffff8000000003fffff0000000000000000000000000000000000000000ffffffffff7fffffffffffffffff00007bffffffffffff073ffff000000000181a5440090108214e72
G2[237] <= 640'h8371ffdfc300831ffffffff8000000003fffff00000000000000000000000000000000000000007fffffffff7fffffffffffffffff0000fbffffffffffe0033ffff80000f8001016a1ca0c963dc0de3b
G2[238] <= 640'h373ffffffc03fffdfffffff000000001ffff800000000000000000000000000000000000000003fffffffff7fffffffffffffffff8000fffffffffffe00000ffffcf701ff0051345ec888a1d20f1ea5
G2[239] <= 640'hf7fffffff01effdffffffff00000000ffff820000000000000000000000000000000000000001fffffffffe7fffffeffffffffffd000fffffffffffe000003ffffff7effc0913460b735b594471d8c
G2[240] <= 640'hfeffffffffffffffffffffffe1f8000001dff000000000000000008000000000000000000000003ff8ffffff87fffffffffffffffff000f87ffffffffb000083afffffafaa24e0600640405b0403cce1
G2[241] <= 640'hffffffffffffffffffffffffffff0000008ef0000000000000007cf800000000000000000000001fffffffffdffffffffffffffffff0000000ffffffe0000001afffff2faa869dbb0675a814303ed6bf
G2[242] <= 640'hfffffffffffffffffffffffffffff0000000c000000000000000fffc00007bfc00000000000000003fffffffffffffffffffffffffc00000000fffff000000002ffffdbffb870f40d28b2c6b680e8d57
G2[243] <= 640'hfffffffffffffffffffffffffffffc0000008000000000000000fffc003efffe00000100000000001fffffffffffffffffffffffffc000000000fff00000000017fffdbeef64c50dac4a7526482b7290
G2[244] <= 640'hffffffffffffffffffffffffffffffc000000000000000000000ffff83ffffffc0003f0f790000001fffffffdfffffffffffffffff000000000018700000000055fffd9fee42f356287c3442086f5a97
G2[245] <= 640'hffffffffffffffffffffffffffffffe000000000000000000018ffffcfffffffc0003ffffde00000079ffffffffffffffffffffffff00000000000000000000001effcdfee4590626c89958088eb74a2
G2[246] <= 640'hffffffffffffffffffffffffffffffe00000000000000000867ffffffffffffff8007ffffff00000079cfffffffffffffffffffffff000000000000000000000016fedfffe561c282462d9920cee6c40
G2[247] <= 640'hfffffffffffffffffffffffffffffff0000000000000001ffffffffffffffffffc0063fffff80000079cf7fffffffffffffffffffff000000000000000000000052ff74f7e45b644816c8c41a04ac81e
G2[248] <= 640'hffffffffffffffffffffffffffffffc000000000000003ffffffffffffffffffff807ffffffc00000073fffffffffffffffffffffffe000000000000000000002faebc4f3d45418416aa8d42d40d6e26
G2[249] <= 640'hffffffffffffffffffffffffffffffc00000000000041fffffffffffffffffffffe3fffffffe000000017fffffffffffffffffffffff00000000000000000000156d78cebf212f1420eb6e401830825e
G2[250] <= 640'hfffffffffffffffffffffeffffffffc000000000001ffffffffffffffffffffffffffffffffff10000003fffffffffffff03ffffffffe0000000000081fc0e40b003feb3df7d66a0bb873e480c02c40c
G2[251] <= 640'hffffffffffffffffffffffffffffffc00000000000fffffffffffffffffffffffffffffffffffff07ffcffffffffffffff01fffffffff00000000007fffffff1bf828b819f9250038007d0a29c539481
G2[252] <= 640'hffffffffffffffffffffffffffffffc00000000063fffffffffffffffffffffffffffffffffffffffffffffffffffffffe01ffffffffff000000015ffffffff93ea11832bf1e8d0c1586dfd96b2988c9
G2[253] <= 640'hffffffffffffffffffffffffffffffc00000001f7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00ffffffffff0000000ffffffffff54b45295b7aa92eb485b8ebc6425d1128
G2[254] <= 640'hffffffffffffffffffffffffffffffe000000e3f7fffffe07fffffffffffffffffffffffffffffffffffffffffffffffe000007fffffffe0010ffffffffffff12709306dfb8df03910c4e2a248e8c5c3
G2[255] <= 640'hfeffffffffffffffffffffffffffffc000001e3ffbffffe03ffffffffffffffff0ffffffffffffffffffffffffffffffc000003ffffffff3c3fffffffffffff04bc3ca1e798cf49e21047bf22180a085
G2[256] <= 640'hfffffffffffffffffffffffffffffffc000083ffe3ffffe01fffffffffffffffc17ffffffffefffffffffffffffffffff800000ffffffeffc3ffffffffffffd78a52a438fd12909b0242eda9c712104a
G2[257] <= 640'hffffffffffffffffffffffffffffffffc000c7ffe1ffffe007ffffffffffffffc01ffef8ff003ffffffffffffffffef800000003ffffffffffffffffffffffae03f5e5b829120710808d94e8a20cc8b3
G2[258] <= 640'hc107fffffffffffffffffffffffffffffc00fffff8bfffc083ffffff9ffffff9001ff800000007fffffffffffff81ff80000000fffffffffffffffffffffff36c380aa8bf9cc718213bcda9ea16b91f8
G2[259] <= 640'he003ffffffefffffc7fffffffefffffffffffffffefffe0003ffffcf1fffffe0000ff000000000000003ffffffe007f80000003ffffffbffffffffffffffffa5673e430528c228e65c92c1fde64f40e8
G2[260] <= 640'hf01fffffffcfffffc01cffffffffe0fffffffffffffffe0000ffff86ffffffc00007f000000000000000fbffe00001000000003fffffffffffffffffffffff85231447b26e31100c406406726339a7c0
G2[261] <= 640'hf81fffffff9c47ffe00037fffffe001ffffffffffffffe00007fff80ffffff800003f00000000000000038000000000000000003bbffffffffffffffffffff513d0c6add52ca10e04d3364d52b421208
G2[262] <= 640'hfc3ffffffffc013ffe0001fffff80001fffffffffffffe00007fff000fffff000000800000000000000000000000000000000000007ffffffffffffffffffe05a4c3092b390b8749fc846c54631a0725
G2[263] <= 640'hffffffffffe00001ffe001fabff8000067ffffffffffff00017ff00000fff8000000000000000000000000000000000000000000003fffffffffe3fffffffc2890b94b31821d06e59380ef81324f02a1
G2[264] <= 640'hfffffffffffc0000fffff0033f00000000fffffffffffe0000fff8000007c0000000c00000000000000000000000000000000000000c7e80e000000081807113a13ba390a44d0fb628ab8cdf8904af2a
G2[265] <= 640'hffffffffffffc002fffff8c300000000000fffffffffff8000fff800000300000000c0000000000000000000000000000000000000000000000000000000b957bd3cf820aa3e827349b2c12450050df7
G2[266] <= 640'hffffffffffffffffffffffe300000000000000003fffffc000fff8000001000000000000000000000000000000000000000000000000000000000000000076ea03bb8e0ea7a44966e8e0a92f2db2004b
G2[267] <= 640'hffffffffff07ffffffffffe000000000000000003ff87f80003ff000000000000000000000000000000000000000000000000000000000000000000000006321c189ab0ddbe62e92060c01bee5860a72
G2[268] <= 640'h3ffffff4000ffffffffff0000000000000000003ff00080001f8000000000000000000000000000000000000000000800000000000000000000000000009fadfbbc932067e7d9254eae34d11f108a18
G2[269] <= 640'h7fffff0000000ffffff800000000000000000039000000001f8000000000000000000000000000000000000000001805c70000000000000000000000000e2166102b470241052d1a42da7c09b1c581
G2[270] <= 640'h1fffff00000000e7ffe000000000000000000030000000000f000000000000000000000000000000000000000000303fff00f0500000000000000000004beca470fbe50c6110cbe34150cbc0a44ec0
G2[271] <= 640'h7fffffd00000001800000000000000000000000000000000f000000000000000000000000000000000000000001607bff8f604000000000000000000005880221c4d1760ba91cb977b977389ed100
G2[272] <= 640'hfffffa800000000000000000000000000000000000000001f80000000000000000000000000000000550080070001fffff9ff000000000000000000003fdea60a66c58553574500182e84ac943104
G2[273] <= 640'hffffff800000000000000000000000000000000000000000f80000000000000000000000000000000ff1fff0f0000ffffffffff0000000000000000007a0b8c0798dda43fd27e20104c16d473ac72
G2[274] <= 640'h7fffff000000000000000000000000000000000000000000700000000000000000000000000000007fffffffe3e00ffffffffff00000000000000000037707a67a2126ffe01fa16489a87fe8db14c
G2[275] <= 640'h7ffff000000000000000000000000000000000000000000077800000000000000000000000000001fffffffff8f00ffffffffff0000000000000000000382d211060f3a6b9ec7c5ea4691508b1852
G2[276] <= 640'h3efffffe00000000000000000000000000000000000000000003f8000000000000000000000000000007ffffffffc767fffffffffff000000000000000010bd1b01cc58a282c021a473be1e1b24b922c
G2[277] <= 640'hfffffe8000000000000000000000000000000000000000000103f800000000000000000000000000000ffffffffffedfffffffffffff0000000000000001427f135fe511011c4c1427d3d0efb85fbd94
G2[278] <= 640'hfffff00000000000000000000000000000000000000000000783e000000000000000000000000000000ffffffffffeffffffffffffff0000000000000000ff1427f9835062b808892085610553a104b0
G2[279] <= 640'hffffc00000000000000000000000000000000000000000000fc3e100000000000000000000000000001fffffffffffffffffffffffff800000000000000045dfc8e31189400553b5769e8ff27c0dcc3c
G2[280] <= 640'he0000000000000000000000000000000000000000000000000e3f3380000000000000000000000000000ffffffffffff07ffffffffff0000000000000040b13b1b8cc4f03baec9a7c183bcc2a8af56db
G2[281] <= 640'he3f1100000000000000000000000000000ffffffffffff07ffffffffffc000000000000000ccffc1447aa90e8b096223b0ed8745220adf
G2[282] <= 640'h3f1f8000000000000000000000000000000fffffffffffe07ffffffffffe0000000000000020db9294c504973960c9481a285c201483b11
G2[283] <= 640'h3f1fc000000000000000000000000000000ffff7ffffff807fffffffffff000000000000043ee50cb450c136142ca239627a444f429bc82
G2[284] <= 640'hf0ff000000000000000000000000000000ffff1ff3ff7803fffffffffffffc000000000066d1ad37b1c27111a91c6ba370121a75e69231
G2[285] <= 640'h70ff0000000000000000000000000000007fff1fe3fffe00fffffffffffffc000000000044c62403f2a258d448d9d1704a3e1af200c024
G2[286] <= 640'hf10000000000000000000000000000003fffbf637cff837ffffffffffffc0000000000124bc2d1d586843392c5eab034441962a2d2f4
G2[287] <= 640'he000000000000000000000000000000007ffff6638c7033ffffffffffefc0000000000276f6a9717e883b28e7684532ca7402437fd8e
G2[288] <= 640'h848000000000000000000000000000000001ff0723f0c0c01c1ffffffcff3800000000002424c94c9a34144bad869f43244a1c9de2c52a
G2[289] <= 640'h700000000000000000000000000000002001f0000f000030807fffffcbf300000000000da9bfe3ac1a14496bef8930452d84e9726e63d
G2[290] <= 640'h3f03ff00040000071800fffffcf000000000000152439b00447b1727bacd0f2525be951fd1f6d7
G2[291] <= 640'h1860000000000000000000000000000000ff03ffc00c00000300000100f800000000000000f261daaa37840da6a8b70002d3003101880f1f
G2[292] <= 640'h800000000000000000000000000000003ff0ffff00000000000000000000000000000000055d14d110fd740795992fdc72d539a3c99f3fc
G2[293] <= 640'h3ffffffe0000000000000000000000000000000003250d247a93e816fd8b848408daaa8be883426
G2[294] <= 640'h8000000000000000000000000000000005ffffe1e180000000000000000000000000000021d071aab9c2037b092c66627677101fa02198
G2[295] <= 640'hfffff161e000000000000000000000000000005ea0d5c79032cb327a12048409dda08e915d73
G2[296] <= 640'h10000000000000000000383ffff7bc1fc00000000000000000000000000000ca8450a54994c605e02870100de427d58e750
G2[297] <= 640'h80000000000000000000000ff7f77fffec00000000000000000000000000040479d15bcb710a5f65d0d402973c11674e468
G2[298] <= 640'h1831fffff000000000000000080000000000916c2c0868cd01dbd6a69ed318f60061240b66
G2[299] <= 640'h7dfff8000000000000001e8000000000b0f329571668d5eb15b8b085980ac252515c87
G2[300] <= 640'hff000000000000000000f000000000000000f1e80000080005120fc4932ab08dbd3cf3f0131130444100497
G2[301] <= 640'h10000000000000000000000980008000000ee000e000000000000000000000000000001fd8c00000e0001eb2ee323320096646bc37d2d33c5e7079499c
G2[302] <= 640'hc00600000000e0ffe0c000000000000000000000000000ffd2e40c0bb803c49532f62e4f2f83f2538193e3f8c99579d8fa
G2[303] <= 640'h10000000000000000000000be07d30000000c1ff00c000000000000000000000000000ff6ee40cff3fffe44afea8846a664da21c16801e839ff83c4a12
G2[304] <= 640'h1af0778400000000c3e000000000000100980000000000036f3db66abe7fff508b21659f06638732413ba1bd54bc1704c08a
G2[305] <= 640'h37df0e386000400e1f81ff0000000000006010000000000007fec253800077e9683309d6a4e4168de3b7063be4230c5c8ccb0
G2[306] <= 640'h1b9f905fbc000c0080f807fc00000000008000000000000000012fa9a7007f8596efca022f11089503648583004d7c60e03305
G2[307] <= 640'h2a3af3ffc0000000017800ff000000000000000301c89000001bfdd07a013fdd8a16a22402048560c0183672f49b0fb6516607
G2[308] <= 640'h863f4efffda000000000500f8000000000200007fffe04fe0ffe6291eba863fdc0235946a4b1624a447d83961daf6499c38cad2
G2[309] <= 640'h3fbfc7ffffe6000000000000ffff0000000fff0c0003fcbf9c0f004710de863c3803c27384b0a51638a055f9917b2c446a00e822
G2[310] <= 640'h7f044ef3fff60020000000003fffff0000001ff1ff20042070c100f890b68000380bafa0965a0e5247e2cfb4881e6c361cb9687f
G2[311] <= 640'h27906fcefffbc790001fffff0018fffff80000007fff81df3e00b07c659900001c230a24992a68867a187b20e0ef4d81c8f95970
G2[312] <= 640'hf7ef91ffffb000c000f3ffff7ffc209f7fffff8009e02eb3e1add3445df8400655e854d2d2e5640f4cb396391faff1b02385e4c
G2[313] <= 640'h8000000000000f0000000000000007fa00dc00031e79f3fff8005ff10e1b0038ffff7e0cff5f3ed8fd73f87b4c00b751994a8c3008c0e9ef498da05210a641681499
G2[314] <= 640'h30000000000ffffff0000007ff001fcc00003216371930f80070000fe0020fe7ffe167fb07ef87c1e00ba4ffc9b6d9c3b0ff110e2b65e7d1ba8f8cbc0d24c424c
G2[315] <= 640'h307fffffffcf3000fffffffffe00001e0bfc100fff7c7a600008000001e006cffffe01738c13f3e7d6be9d3ddffd1d1a21ff0c104f1ed6922cce2d952342e444ceb
G2[316] <= 640'hfffff8c0000fffffffffffffffffeff800ffffff87e3e1fcd8c78080069804000300c007ffe01f80011fbfd7f88df3f5ffe7f764a5797a8543523637a62062531fff948e50
G2[317] <= 640'h7f1f000000000ffff800000007ffffffffffff00000fffff000000e3ffffff003000fffc017e39749c031001800001fff80001001fa50ba24dc2017fa6537ee0b9b224a652210b9c4bf2d9491d2ee400
G2[318] <= 640'hffffffffffffff000000000007ffffff00030000000000077ffffffff000007ffe83ff8f7f7f1337808011013f38000000fb0758e9608f117f1db27c50389516039a8bad0ee1e21a542becce8b
G2[319] <= 640'he3ffffe0000000fff800000000000000000000000000000000000033fffffffe04601fff83fff0ff90efe6400001002000001e41fb78e66ded38df7f9e8d8e526a7858d30886defb62cad4bf1fa85236
G2[320] <= 640'h3ffffffffe17ff83ffe7fffff97f3fffecf100000000011ef6449a63e572f8a837d25780e6a3388e4b814ef2e280092aaa8802bf81
G2[321] <= 640'h1fffffffff7ff80f83ffffff9dffc014f1f00000100303f55b4a910d8c95b2613a146ac1a8cb4900141844e2d61873826d4501161
G2[322] <= 640'h1fffffffff37f000839fffff801ffffffffa000000003996d2f604556d59a5403a966f71aec11b002879a0ca1e01060932f407267
G2[323] <= 640'h3fffffffff37f000001fffffc1d7f386dffe50000000299ca0530edb5005176542b83c17f81801038009b459fcb61458462f66e4c
G2[324] <= 640'h7fffffffffffff0000007ffff9070004cc7f9800000f09f3a7c865851278cdc1b007aa583086e04583429122149e212d281646e13
G2[325] <= 640'h1ffffffffffff10000003fffe80b80000ffff7e00030f0e2de6706d1fb01e4112d991f1988f51421440bd47208a1b9fd165126270
G2[326] <= 640'hffffffffffff7f8000004effdf9d01cffeffe0fc0000004f4fadc7a01a73bffa09df0b2edc7dbe34140746d7189aee620e362283
G2[327] <= 640'hc00000000000000000000000000000000000000000000000000000003fffffffffffffffcff0001ffc0000000001fbc000001dc89bb7a7a49475a7a5880f0f1bd46136c4b970176c0015fe2a5205c0b
G2[328] <= 640'h3fffef000f080f8000000000038000000000000000040c100c000000000fffffffc800000007fffde3c84000007c033f980010425d871b8404510596e1e34733c05883a45c92d298493605df21e094f
G2[329] <= 640'hfffffffefffffffff0e0fef0ffffffffffffffffffffffffffffffff0ffc0000000f3fffffff8000703ffffffbfffc63003ffcb0abaebfc65be5eb5bb7e0905a0181341417487784c05c799210347f17
G2[330] <= 640'h80001e00ffffff000000ffffffffffffffffffffffffffffffff007fff009fffffffffff03000000000ffe0000c0fc30807ffc2363d839695b2fb30b6aed005d4802d21c8f40861c4014d60a1dd66452
G2[331] <= 640'h1effefffffffffffffff800000000000000000f01fd000000006ffffffffffffffffffff007ffff6fffffffff83ffffce001fc612f1e15f35362614860fa6a649187cda0632a12a9c05b14f229084308
G2[332] <= 640'h1c03fffffffffff3fffffff87ffffffffffffffffffffffffffffffffffc000000000000000007ffffefffe8ff84000e000fdd4f73f20885836af22526697637e120f20c5a3714800c861db7464528e
G2[333] <= 640'hfe1e000000000000000000000000000000000001ffff037eff8f000000000000000000000000000003800108010000000000a3e806e9085b30f742c37fda963d38c1188a5147810a00bbc84eec6e44ee
G2[334] <= 640'he101c00000008000000000000000000000000000000000000000000000000000000000000000000004000000000000000000b7d28e8369b3cb4d9dc98332e31915ca4c840c4885f0016dd1760c642683
G2[335] <= 640'h7c03be000000000000000000000000000000000000000000000000000000000000000000000000001c0000000000000000015033f60705fc46bd653e0926181b84cb2b80e83951fd8425d99813181ae2
G2[336] <= 640'hbb807effc00083c0000000000000000000000000000000000000000000000000000000ff000000001cff019000000000004967c86918f10f0f13925a4d2efb7984adcc84618ca4d6c447da528d08538e
G2[337] <= 640'hbbff001fff8007c0000000000000000000000000000000000000000000000000000000ff0000000000fe00086100080001003449e68246b4923f708e6eb7bed068a4028a4182a54c840478170f987693
G2[338] <= 640'hff007fcfffc31c0300000000000000000000000000000000000000000000000000004cfffccc00000000000000074ff103b6ac3fffdc3df01914132eae4e366b17c38585711b28bf0807ac6b457218b1
G2[339] <= 640'hb3c07f07f7c03c03e000000000000000000000000000000000000000000001000000fcfffff83800cfc000000003effffcbf595b85fe56187775b9e8e9786f3f45677ce11a8c7a28406828de79a22435
G2[340] <= 640'hfeffec0fff300000f0000000000000000000000000000000000000000000070f7fffffffff700ee0c7ff8f1000004f7fff785e8916522a604a27958323125e88e52092491a4006c11400bceed1005701
G2[341] <= 640'h33ffe97ffe7c8100f800000000000000000000000000000000000000000007ffffffffffffe006fffefffffe84307ffe03782c2281b98f442002b38d73359775c55404e0930945c38071193045414464
G2[342] <= 640'ha6fe607ffcfe0000fe00000000000000000000000000000000000000010ffffffffffffffff76fff7c7fffe0463fc06007017a6cea0690e77c98aa272d98371060e8110111732c4c8464e77f21e64027
G2[343] <= 640'hdff600ffff0001e3d0000000000000000000000000000000000000107ffffffffffffffffff2ffcfcfff01cff8fd10c0c0505bfffe757505e861f0f28932e502079021304d440a286031e9a1ad2052d
G2[344] <= 640'h3ffe007ffff771fff0000000000000000000000000000000000010383ffffff6dffffffff7fe7eedcfbf3f819e7e038c76d281f2a20a1c91a9372f56a340ec19282a899c5482f941b1a9ea65611284e
G2[345] <= 640'h1fff007ffffffffff0000000000000000000000000000000000000fff010cffff375bffffd1fffffc3b0200ff01ffc0006e5fc0da89c05b1b8f176ee92e8517b2c45a0190a582048d2b9b24fce87b10
G2[346] <= 640'h3fff007ffffffffff0000000000000000000000000000000000000000ff6f07a35bffffffbdfff63c3405ffff81ffffffcc4639ddfc86f6d9078061f776aec259f8608050c1983c0232915088e00946
G2[347] <= 640'h1e36006ffffffffff00000000000000000000000000000000000083c798457eb49f0fe4fffa58462c32fcffffe3dfffffff9fc25a7737a239ad18f6d8a0ba0555d4441c80602160001a4613ab441e52
G2[348] <= 640'h3c3000000017fffff80000000000000000000000000000000000104e67c6f7ff282b7100ff6567fc57b00c1fff93fffeff9e05d23be987c04827e4fec88b2c2e23a0160c86c28cb2482b36240402747
G2[349] <= 640'h3fe3f98000007fffffc000000000000000000000000000000000003ff739efc1bba232378e8dfff6d55fffffffcfe264002d0b9b3451899bb688958aff2e81c5d0dbb5842449e80199442406e843d51
G2[350] <= 640'h9fffffcc08007ffffffc0000000000000000000000000000000000201fffff819c19560878c4bf0f25321cfffffb00fba012fd437191627db8bbc881eecb6c199e3c048074c69dc2584a0109682335c
G2[351] <= 640'h3ffffdc03800fffffffc00000000000000000000000000000000003063fffffa961f3fe0614b41febdbfe3fffff9c03cf905062b1c0979a997b2c378c407392ddbe66004502604046421856dc520949
G2[352] <= 640'hafffffcc0001fffffff8c6600000000000000000000000000000000ffe1ffbc7ad38a9d56249940bc91edfff7ff821f8efa526862609c167f9674d0c37a55a0310798b0c18a1c98074208482c443512
G2[353] <= 640'h3ffffffc000003ffffffff0810000000100000000000000000000007fff067b67ac01e240745abfbb9a407ffff9c20e0002ad74b15623ce114a49e12210affc6fb907f0001a31761002822304c2468e
G2[354] <= 640'h3ffffefff0000003ffef3ffe1018000000000000000000000000000ffffe0ca88321e8dac884fa059f6a980036006060025f3524b1ce59ecfe121d6bb29321ec95f424c4f0202b33605c2206c902b0b
G2[355] <= 640'h3ffffffffff3803401ffffff8f80fffc100000000000003e0000ffcfffff6647cc50984eeed59504f29c0f80008f0003c2d6eee5d9a43ccd6f7b94ff0846db48c052e60230283640b20390088d03a81
G2[356] <= 640'h3ffffffffffcc000410f00fff7fe07fc90000000000000ffffffffffffffe30a960288d7034b30c00699bfe07470ff97cbc99ee7814132769ead2bc80ad18af442af0200081c1306b00218a70581e02
G2[357] <= 640'h3ffffffffffce000039f1ffffe0387f3d80c3c7000000013ffffffffffffef3ca9dd0eaf40e07c00da8723fffde3ffffc9740a0108aaa2d43d50d123f130178a226004d0200ec5c03011080abda0320
G2[358] <= 640'h3ffffffffffcffc008001ffff0300006e3f9ffe70000000163fff1ffffc7ffb39e64571f12489007505320000e13ffffe9ee28ca0ed9583b2111687de8969998f118ccb0000200290300010228a75b1
G2[359] <= 640'h3fffffffffffffefbffe6410199afffe0f801ffcf200000bffffe00fe6601fb5d2595e09210fd2c47cf38007f013ffffe9c9c705f4b727d01481541af5b43eea0041c2000012008c04826018bd40100
G2[360] <= 640'h3fadfffffffffffffe3ffff1f7fff5fbfffffff3f0b063fefff7c0002c07c6aa616e1e2d125551c49c68801fe1a2ffffede3f7c827b4939492f43d4402033731012606300c6c03040e0330008407800
G2[361] <= 640'hadabbb7ffffffffffffffe2fffffff03ffffff8ffc0f70ffffcc4000018f0738373a820ef1de9e289939203fc1c47ffff566748325b39b35828c43e814b541c0207200e80001810c800206446442409
G2[362] <= 640'h1f2011ef1fffffffffffffffffffffff5ffffff0107e9ffffff08000007e70235810ac4743964a7c955883fffc400fffffc30c908d8b9c88847c4edfb062006eca081301c3410811201002480aa63f00
G2[363] <= 640'h1c0001bffffffffffffffffffffff405dffffc7fff00efffff0002462070c2a62c8860c86e650046615e11ffc760f7fff1be1ed0311a7087a3c0c9755e8e061739911800131ce08e23000c019c60108
G2[364] <= 640'he80003d7fffffffffffffffffffffe073ffffffe000c3ff7fe00004e007001d187596d22a799f1133c0621ff8f5947fff6943e95954a2550d1df847f518a0b0e182104c40804b08020410440042080c
G2[365] <= 640'h13000309ffffffffffffffffffffffe057fffffffc00000061e40041f09f3046448baa2f1c84020046a0049ffcfd387fffe8ccb83e0a40fb254417cc19f79cd3c2c0000780100000320000c09020020c
G2[366] <= 640'h1c004001b3fffffffffffffffffffff07ffffffffeffffc00007b14867c0df78ab228388461e0572b4ea90fffc565c7fbf2462935e31361da80863d7fd35cb1201b0003680003c01f230004080061022
G2[367] <= 640'h80000109e67fffffffffffffffffff057ffffffffffffffc181ff565fff106d1a1d65bb36c9fb44dcbe487ffcf67eff3f915c8200628c738f3ccc4335988a9b20c81b0830d028005000000043840060
G2[368] <= 640'h806e597ffffffffffffffffd07efffffffffffffffcc06ecda3dda53e5e477b249d4e463dc3bbc17ff27522575ee576cea3f0fb63c0fb046c0d571a1c0000390050c05c0182000000002a30a8
G2[369] <= 640'h800a0bfff9bfffffffffff003fffffffffffffffffc03d50a13c34bd290dd268770723c8be76b97ff04166962e4b880ba034d148b1ec64773d8e0e502480022850444e00b88c000001a0208c
G2[370] <= 640'h700103df1cdfffffffffff700effffffffffffffffc03f2ea0271825a26014307c9a4db4714a5c7ff7e06e8602111622c2433714e9d238bc09a5314bd4823ae2080043100d800000113300a0
G2[371] <= 640'h100001267dffffffffffff63b0bf7cffffffffffffe3ffebd06419accf9167e898f084f0a1d2c97ffce1fe67935a43faa4a78631811bc1f298e5833b4b4287e9080000100c020300806400ec
G2[372] <= 640'hf00001276e7f9fffffff99403180ffffffffffffff1f99823f1216624ba41f5bc897d487027e83fff7031612e4e0a82578facadd80b763660250f28634802d2000020003300020080100008
G2[373] <= 640'h21000001dd0ffffffffefc0023fc0f387ffffffe3c3e4ea0322334e0a9d113a11cbddefd076dd7feda6471c127c66b9a20279097a810e7ea20d3a044000c3a0800012000a1c000000620002
G2[374] <= 640'hc1c00000c339ffffffe800007fff4007f8ffffc007b8543e2ad051dd13908533905e11558135fcc18296fc4265b141461d5cc0e2862c71f9d4001950096611cc001318101a06000020000c
G2[375] <= 640'h1803800000d6bfffffe000007fffffe0007f800fc0cdbb651750869bc53361220a824c91eb2080184429fb0f3b0224073724a309c68c5702a44e31a0c0336b80001008201a0000001b0000
G2[376] <= 640'h2780e000020dffffde000007ffffff9f1815ee000e041bc3a60d80a0086454781c72895947233e04487f94387f246023e88229383cf5453a83c860008c0a9000000000038080000010005
G2[377] <= 640'h7ff01f000005ab67e000017ffffffffc003e019e70ad36ee4672193b158844476c5696b85de3cc993fe0df4e404a600804e0ab85de8c0088120db000d0c4c0030044000c180000000008
G2[378] <= 640'h7fffe0380001cfbf100000ffffffffe0103e019f5b4442b577d2044002e65ba4410ed30bfbc78412b5d091017412908baae31238f216b2118f1e1084409008030004008c180000000000
G2[379] <= 640'h231fffe0380002d1f80003fffffffe03fffffffcc1215740e20028a4d63c64a4af30f80af10fd1a176803100280580010d6ae82036401125532141a69e0c580000000080000000000000
G2[380] <= 640'h1cc47fcee0f80024240003fffffffc07fffffffe05709f10bc4da1624a54e486023dfc16b8c7cf8b920c76e33000000000932aa83c94904c630f26426c0c000000000000000000000000
G2[381] <= 640'h3ffe030ffe1c0021c0003ffffff001efffffffd7a110021781cbc46bf0fea43184db23767c7f4ea8053025f0000002000158114a75c23e5f00384603801000000000000000000000000
G2[382] <= 640'he6ffc1ff5f1f80000001783fff3f3ffffffffdb739ba3a337e20808dd5a1e11fe9b8e981bfb87aa21ea0f4000000084000b004b44e9923018346006200200000000000000000000000
G2[383] <= 640'h137fffb3bffe84000003b7df7f7fffffef7ffca7a6916e1b4a2c82088d663f6fa4ea1de2e3d4f59048f06000000000000223c33a1d704e188064200000000000000000000000000000
G2[384] <= 640'h1f0fffffc79fffc0000168b7ffffffffefff76863c71c81d62cc76e20fb0b6a181c80042eb962d09a00a0000000000000001fd6cd4a362848ce4300000000000000000000000000000
G2[385] <= 640'hcf907ffffff9ff018003805bffffffffffece3f590a0c0a610d07f896e1c1ee768051db44251fb795000000000000000000f42ad5f306058346000000000000000000000000000000
G2[386] <= 640'h30ff007ffffff0fff400003fdffffffffffee5e4898c0c4046b8082625ab4da74404a1bcd25f48c22000000000000000008060247276f008680000000000000000000000000000000
G2[387] <= 640'hc7ff000f7ffffc7e767f80ddffffffffff50aaa0191a0d28f0066b107ad211e1ec4df2de26f81408000000000000000000000000020085c3e0000000000000000000000000000000
G2[388] <= 640'h303fffe30000ffe70763b47dffffffffe38037a0d9aa47488360557f10604003004398054748226c800000000000000000306202000001c000000000000000000000000000000000
G2[389] <= 640'h1903fffffffc07f0ffffff1bffffffff0f80031888543b1602630eb52422e90080042a1241bc58640000000000000000008402108048000000000000000000000000000000000000
G2[390] <= 640'h38000000000000cf000ffffff783ffd9f2b8efffffffe10240000004075144a524c03a08200003440635234449f0000000000000000000048020000c0080000000000000000000000000000000000
G2[391] <= 640'h6c00000000000023ff001307fffe07fff6ff23ffffcf406894220240093aece6a0552140000017a08b8100bbc2000000000000000000000b2022444000a0008000000000000000000000000000000
G2[392] <= 640'h68000000000000083ff0301c0c0fff81ffffc78bffc003f99c0004720032ec940140f40000000031c2900000000000000000000000000000000646280000000000000000000000000000000000000
G2[393] <= 640'h3c0000000000000307ffeffffff07fffb7ffe08322303ff9960000000000431d15c67e000000000000000000000000000000000000000000000646380000000000000000000000000000000000000
G2[394] <= 640'he07fffffffffc07fffc7f4217fe00000000000000000094bb50840000000000000000000000000000000000000000000800246280000000000000000000000000000000000000
G2[395] <= 640'h3f0037ffffffff803fff0f8118000000000000c030f8004f2740000000000000000000000000000000000000000000000002c4080000000000000000000000000000000000000
G2[396] <= 640'h1ffc00187f000fff8e7ff2e0080007fc08000081f8fc00000400000000000000000000000000000000000000000000001000c4000000000000000000000000000000000000000
G2[397] <= 640'hc3f8c004037007ffe03f26863e037f00cc00003b83805210020000000000000000000000000000000000000000000001000c4000000000000000000000000000000000000000
G2[398] <= 640'h303ffeffffffe007ffec6d40ef03ffe2640020f80f974c1820000000000000000000000000000000000000000000000fa6004000000000000000000000000000000000000000
G2[399] <= 640'h207fffffffffee020ff9be43382dce660006038085e2c1840200000000000000000000000000000000000000000000fe4054000000000000000000000000000000000000000
G2[400] <= 640'h100041ffefc8fff7c1fffff01820070600060300c9ffe88200000000000000000000000000000000000000000000002921c0000000000000000000000000000000000000000
G2[401] <= 640'h4c0000ffe0017ffff87fffe102000000001f13c49ffc8020000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000
G2[402] <= 640'h4ff00000000001ffffe0fff003800000001f13e38fcf8020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[403] <= 640'h10fffc0007ffe0001ffffffc03018000000d12e3c06e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[404] <= 640'h40ffffffffffff0001ffffc00008000000003f8c0060000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[405] <= 640'h7fffffffffff007fff80000000000003f800060000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000000
G2[406] <= 640'h600000f800003ffffd07ff600000000000017000060800000000000000000000000000000000000000000000000000000003e00000000000000000000000000000000000
G2[407] <= 640'h3c00000000800006ffffcfd80000000000000000040800000000000000000000000000000000000000000000000000100003700000000000000000000000000000000000
G2[408] <= 640'hff800000030f00020fffffa00000000000010000e0000000000000000000000000000000000000000000000000000100002200000000000000000000000000000000000
G2[409] <= 640'h33ffe0fff7ffff800001fff8000000000300000000000000000000000000000000000000000000000000000000000000001c00000000000000000000000000000000000
G2[410] <= 640'hc7ffffff7fdfffffff07be20000000001e000880000000000000000000000000000000000000000000000000000000000082c000000000000000000000000000000000
G2[411] <= 640'h2001780780000f8fffff8f983000000007400000000000000000000000000000000000000000000000000000000000000006c000000000000000000000000000000000
G2[412] <= 640'h80000010000000000fffff22400000001b400800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[413] <= 640'h218000000008000000077f30c000000003d00900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[414] <= 640'h1dfc4001cfffff97fe0010cc0000000000620340000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[415] <= 640'h43fffffffffffffffffb3f90000000000380040000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000
G2[416] <= 640'h10100611800000031f73ffe4501000000056000000000000000000000000000000000000000000000000000000000000470000000000000000000000000000000000
G2[417] <= 640'h40000000800000000010091bc2000000014400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[418] <= 640'h18000000000007c80000638800000000004500e00000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000
G2[419] <= 640'h7ff000003ffeffff8cfffff000000000002a02c00000000000000000000000000000000000000000000002c0000000000000000000000000000000000000000000
G2[420] <= 640'h3fffffe7ff0c00018c00998400000000002a8090000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000
G2[421] <= 640'h80cfe0fe000000000000096000000000003c00a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[422] <= 640'h600000000c0000000006610000000000002fc01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[423] <= 640'h8000000000107ee1c78b152000000000007e00c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[424] <= 640'h210039c003ff01000100078800000000001fa0300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[425] <= 640'hef07f037c80000000000003000000000005ec000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000
G2[426] <= 640'h3f88e000c00000000000020c00000000000b5000000000000000000000000000000000000000000000003b00000000000000000000000000000000000000000
G2[427] <= 640'h18000000000000787000000cf0ffc00000026000000000000000000000000000000000000000000000003800000000000004000000000000000000000000000
G2[428] <= 640'h40000000001fc00000000007ffff8606000a000000000000000000000000000000000000000000000000028000000000004000000000000000000000000000
G2[429] <= 640'h100003f080ffc0000000000f00e1e0f80000000000000000000000000000000000000000000000000000060000000000000000000000000000000000000000
G2[430] <= 640'h2ffe3ffff0000000001218083e7f8388000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[431] <= 640'h1fff80000000003ffe780001e3c0d810000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[432] <= 640'h400000000000ffff8000000dff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[433] <= 640'h30000000003ffef880000084fe00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[434] <= 640'hc00003c83ff0c00000007d80000000000000000000000000000000000000000000000000000000000878000000000000000000000000000000000000000
G2[435] <= 640'hc81ffffff000001887fe000000000000000008000000000000000000000000000000000000000000030000000000000000000000000000000000000000
G2[436] <= 640'h7fffe138c000037ff800000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000
G2[437] <= 640'hfff00000030fffc00000000000000000000000000000000800000000000000000000004c0000000000000000000000000000000000000000000000000
G2[438] <= 640'h63c0000007ffe000000000000000000a20000000000000000000000000000000000000380000000000000000000000000000000000000000000000000
G2[439] <= 640'h100011cfffdc0000000000000000000fdc009000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[440] <= 640'h41cffffe0000000000000000000000fe00a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[441] <= 640'h30ffff2000000000000000000000007d7f20000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[442] <= 640'hcff800000000000000000000000007c3fe0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[443] <= 640'h3d8000000000000000000000000007c7f80000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G2[444] <= 640'h3ec000000000000000000000000000000000000000000000000000006000000000000000000000000000000000
G2[445] <= 640'h12000000000000000000000000000000000000000000000000000000a000000000000000000000000000000000
G2[446] <= 640'h12000000000000000000000000000000000
G2[447] <= 640'h1f00fb100000000000000000000000000000000
G2[448] <= 640'h40000000000000000000000000000000000000000000000000003800000000000af6d20f00000000000000000000000000000000
G2[449] <= 640'hc000000000019fd900000000000000000000000000000000000
G2[450] <= 640'h240000000000000000000000000000000140000000000000000000100000000200284200000000000000000000000000000000000
G2[451] <= 640'h6400000000000000000000000000000000600000000000000000001400000000f0183e00000000000000000000000000000000000
G2[452] <= 640'h80060000000000000000000000000000000000201c000340000000000000000000000000000000000000000000000000000000000000
G2[453] <= 640'h7800000000000000000000000000000000000003033000040000000000000000000008000000000000000000000000000000000000000
G2[454] <= 640'h7e800000000000000000000000000000000000006086601818000000001fd3000000000000000000000000000000000000000000000000
G2[455] <= 640'h608000000000000000000000000000000000000140030c001cf44f31000010000000000000000000000000000000000000000000000000
G2[456] <= 640'h6e0000000000000000000000000000001180380000602bff00c70dbff4cf8f0000000000000000000000003806c0080000000000000000
G2[457] <= 640'h60000000000000070007a280000ff1c001801e80000430001f7eb4a006034a000000000000006440000000c000010c0000000000000000
G2[458] <= 640'h9118cf738f81ff1800000038000087ffffe80075b83014a00000000cc007bcc7c000100c00000000000020000000000
G2[459] <= 640'h1000000000000000000000000000000000041080003fc000000000000000001c000006c00d900c038388000000cc002004280000002400e0000000000000000000
G2[460] <= 640'h8000000000000000000000000000000000000fe00874500fb8308000000cc00602c688000183c0000000002000000000000
G2[461] <= 640'h80000000000000e0000000000000000000000000000000000000000000000001103000f9419f10003608001000c40024746c020000400000000000000300000000
G2[462] <= 640'h80000000000000e0000000000000000000000000016000000000000000000018e1001f0c406500002c94800000c00000000c000000c00000000000000100000300
G2[463] <= 640'h16000000000000000400000000001f2f80000000000000000183000f25200331000181f308000400004046c0000c3000000000000000000000000
G2[464] <= 640'h7200000000000000042001043c080000000000000000000000920e3d2c0008e80001a14024000000020047c0000000c0080000000000000000000
G2[465] <= 640'h100000000000000000000000000000000002610984000000000000000000000000001f97fe00000877bff0b0960900c0200143c640000c08c000c000010000c01c00000
G2[466] <= 640'h700300000000000000000000000000000000000000100840000000000000000000000000000000000000000300da5cdded1c00003e3847001fe7ff003c000018000000000000
G2[467] <= 640'h3ffe4fe00100000000000000000000000000000000000000c4f780000000000000000000000000000000000000000020123fb000000000000000000000000000000000000000000
G2[468] <= 640'h1e381ffff6bc0fac00000000000000000000000000000000000184418a00000000000000000000000fffffc000000000083c010c18200000000000000000000000000000c00000000000
G2[469] <= 640'h3e387ffff29bcb90000000000000000000000000000000000000c600e8800000000000000000000007fe87400000800000e9c715fef4000018000000c3ffff0010061001400000000000
G2[470] <= 640'h3fffff901fcd80000000000000000000000000000000000000c004732000000000000000000000047f00000000800000045632001bc1000818c700c100fc0000180400000000000000
G2[471] <= 640'h1f3ffffff901c0100000000000000000000000000000000000000420c7ec30000000000000000000007f8008000701c00000000c01880c1000130460000c040000fc088e8480007d00e00
G2[472] <= 640'h7f00000004ffffffffffc360c00000000000000000000000000000000000001040007e7b00000000000000000000073ff9802201040000000003c0018800042067209cdec3a31900492c800353680800
G2[473] <= 640'hff800000c7c7ffffffff8700e00000000000000000000000000000000000001000007ef00000000000000000000001807d00308100000000000007014a00001880011800080cc98770717c0362000000
G2[474] <= 640'hff0000ef41ffffffffff8700000000000000000000000000000000000000001000003f780000000000000000000003ffc0063801c00000000000001e63c0000000000027f10f83fec800f60010000000
G2[475] <= 640'hfffffeffc3ffffff3ffe8930000000000000000000000000000000000000000000003f400000000000000000000006c004021900000000000000000060200000000101e00008080010250e0000000000
G2[476] <= 640'hffc7ffffc5fffffcfd7f2390000000000000000000000000000000000000000020003f943c000170000000000000038000031de000000000000000000000000181780c000ee9443c003b910000000000
G2[477] <= 640'hfff00efe5f3fffce076c800000000000000000000000000000000000000000040001f80220006080000000000000000000098000000000000000000000000011270702df7058c074c038a003800000c
G2[478] <= 640'h7f73fffc1f1ff7c7fff800000000000000000000000000000000000000008004000008000000278000000000000000000006000000000000000000000000000025a071fe00e01c3c0000000b20a000b
G2[479] <= 640'h1ffffffbc1f8fffcfff8028c00000000000000000000000000000000000000002000000000000078000000000000000000000000000000000000000000000000002d3fd1cc00c6e000f8000026c40a00
end
always @(posedge vga_clk) begin
G3[0] <= 640'hf08cc0e087c0ee008100000080000000000000000008000001000020000000000000000000006000000000000003000000801f037fff
G3[1] <= 640'h200ff8c30f0c186e600000000000000000000000000000100000000000000000000000000000000000000000000000000000000f8f0feff
G3[2] <= 640'h3001fcc3cfce00363000000000000000000000000000000000000000000000000000000000000010000000000000000000000300f78fcff
G3[3] <= 640'h13c000fc03cff00716200000000010000000100000000000000000000000000000000000000000000810000000000000000000101241e78ff
G3[4] <= 640'h13c0000e003ff00306400000000010000008100000000000000000000000000000000000000000000810000000000000000000180e003041f
G3[5] <= 640'h3000070800300006c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000c66c1071f
G3[6] <= 640'h20000710003010c200000000000000000000000000000000000000000800000000000000000000000000000000000000000000807e087df
G3[7] <= 640'h8000000000000000000000000000713000c0c82100000000000000000000000000008000000000000000000000000000000000008080000000000000000003601ef0fc
G3[8] <= 640'h70018c0fff00003000000000000000000000000000000000000010001000000000000000006000000000000000080000100110300893c3f
G3[9] <= 640'h1001800ff8c000000010000000000000000000000000000000001000000000000000000000000000000000000000000000001000181383f
G3[10] <= 640'h31000031008c80e000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000081007f
G3[11] <= 640'h300000310084c0c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010163
G3[12] <= 640'h83f0000000000000000000000000000000000000000000000000000000000080000000000000000000000000000080000101e3
G3[13] <= 640'he1e000000000000000000000000000000000000000000000000000000000000000000000000000000080000000000000000023
G3[14] <= 640'h800000807fc00000008000000000000000000000000000004000000000000000000000000000000000000000000000000000000001000023
G3[15] <= 640'h300000000980000000000000000000000800000807f8c0100000000000000000000800000000000000000000000000000000000000000000000000000000080000000010001040833
G3[16] <= 640'h100000000000000000000000000080000000000800004060001000800600300000000000000000000002000000100000000000000000000000000000000000000000000000001000000000000070880
G3[17] <= 640'h100000000000000000000000018800000000000000000000001808001000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c00800
G3[18] <= 640'h10018800000000000000000000030018001002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000700
G3[19] <= 640'h66000000000000000000000100c001000000000008000000003000803c00400000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000001070e
G3[20] <= 640'h66000020000000000000800000c000800000000000010000000118881c00c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000070030e
G3[21] <= 640'h600000000000000001080000038000000000000000000000001080883802000000000000080000000000000000000000000000000000000000000000000000000000000000000000001000000300100
G3[22] <= 640'h8801008000000000000000000018800000000000401000000000000001000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000038000
G3[23] <= 640'h980300830000040000011cc0008380090021000000c00000000080001800020000020000900001380600000001000000800000000000000000000000000000000000000000000000000080000080c0c0
G3[24] <= 640'hc1f80000001032104c100820001000000000001012000000000008000000000000000000000008100000100800000048000000000000000000000000000000000000000000000000006000000000003
G3[25] <= 640'hf8e0800000010060040700120618000080000020030000000000008000000000000000000000001880000000800000040080000000000000000000000000000000000000000000000000000000000001
G3[26] <= 640'hfcc11800000100e0000300120038c00000000000000400000000000004800000000000000001010080000000000000060100000000000000000000000000000000000000000000000080000000000020
G3[27] <= 640'hcf8730000001000000c00012f03c03000000000e000000000000000000000000000000018001018102000400000000060100000000000000000000000000000000000000000000000000000000000000
G3[28] <= 640'h871c41008001010001e03c3207ff00000000010e000100000000000020000000000000008000000012000c00000000022100000000000000000000000000000000000000000000000000000000000001
G3[29] <= 640'hc0f8c100c0018007033fffb21fffc0000001018c1c1100000000000000000000000000010000183cb000c00100000000200000000000000000000400000000000000000000000000c000000000000001
G3[30] <= 640'hfcf08e000001000633ffc3b7f8fec000000080000e9000000000000000000000000001000100037e3000e001000080000000000000000000000000000000000000000000000000000000000000000001
G3[31] <= 640'h1ec38cff0010078e3fffc3b71efc03000000fc0000808400000000000000000000001100030383e71030e130113ec6000001000000010000000020000000000000000000000000000022000000000081
G3[32] <= 640'h3ef0191e86198efb03ffffdf3bfc789c000016013001980000008000000000000000000100870e98c1463000000e0166f109000080001800040000800000000000000001000001000000000001000000
G3[33] <= 640'h3c3399388311ce3f07ff7fffff7fe199000032010003980000000000000000000000000001c01e98e006b001038e31671949000084000000000000800000000000000000000000000000000000000000
G3[34] <= 640'hc30fd9e0816038079fff7fffffffe31300009220070161000000000000000000000000c0031ef8f8f8060200c1c4fb061849000004c08100000060800000000000000000000000000000000000000000
G3[35] <= 640'hccc1e101663cc3defffeffffff3e11803c17300f3c63800000000000000000010001801f1ffbfcf8068280e0c4ffe0f869000000c081009000f0000000000000000000000010000000000000000000
G3[36] <= 640'h3cecc7c731669ee3defffeffffff7e98c03f0300181826800000000000000000802101041cf0ffffe306f0803fcf1ff0f169000000000000110000000000000000000000000000000000000000000000
G3[37] <= 640'h3cfe670f3c66ceffffffffffffffe79ccc3fb2c018088c0000000000000000000000000cc3f37fffc70633047e3f0f99e74d008000010000010000000000000000000000080800000000000000000000
G3[38] <= 640'hff7f7efffe8ce7fffffffffffffee7fccc83b0c0181f990100000000000000000800001fc33f87ff1ee4330ef03f0ef9674c800000000081000000000000000000000000000000000000010000000000
G3[39] <= 640'hff73fefccf9973fff3ff7efffffffef9dc03b2c0c73f9b300000000000000000000ce07fff7f86ff3ce4708c073ecef8744cc000e30000c3041800000400000000000000088000000000000000000000
G3[40] <= 640'hff7f7f78fffc7c6edffeffffffff3fcffcfffe0f1fe3fe00010000000000000001e0e1ff7f67fffec77f00717ffc19ffce4020e01806e798000010800000000000000000000030000000000000000100
G3[41] <= 640'hff7fef3fff7ffffffffffffffffffccff3fffffe3e1fff8000000000000000000100793fff7fffffc0efe77ffb7cb9ffffc071e1c0060018000081000000000000000000000120000000000000000000
G3[42] <= 640'hff7fe67fffffffffffffffffffffffff733efffefcfcfbc0000000000000000000003d3fe3fffffffee7e71ff07cff3f71f8f9e3c0067e188f0081000000000000000000000100000000000000000000
G3[43] <= 640'hffffe7fffeffffffffffbffefeffdffeff9efffffcfc73c00000000000000000000273f3e3ffffffffe3ff8ef0ffff7f73fff9f73806ff09cf0019006600000000000007000000000000000000000000
G3[44] <= 640'hffffe7fbfffffffffffffffefffffefefecf0ec33f8e33000000000000000000000777f3ffff7ffffe387fccf0c3ffffc7ff80371802ff01010018006600000000000007000000000000000000000000
G3[45] <= 640'hffff677ffffffeffffffffffe7fffffffee71fe03f8f1700000000000000000000c77eff7ffe7fffef383cf0f1c36effcfff803f83023c812000c1006200000000000000000000000000000000008000
G3[46] <= 640'hffff7fffffffffffffff7ffffffffffffef3fffcffff0f800000000000000000067ffffefffefffffffc7efbffff6efff3fecc31c1020091780081000000000008000000000004000000000000000000
G3[47] <= 640'hffff7ffffffffffffff7ffff7ffffffffffbff3ff8ff8fe008000000000000000e7effdffffffffffffffffffffcee8ff1c0de307806e7d908ff18381800000003000000000000000000000000010000
G3[48] <= 640'hfe99f3f93ffffffffff3fffffffffffe99de7fd387707fe0000000000000300133cffddfffff7ffffe67f9df787e1c7ffbfcfe71cffc30e07e7098e000301c7000810100181860800000000000000000
G3[49] <= 640'hffff737fffffffffffbfffffffffffff99dfffff0f7b7fc00000000000002018fffefffffffffffffffff9dfc7ffe7fcff1ffeff80e37183000101000000808100180100810020000000000000000001
G3[50] <= 640'hffff777ffefffeffffbffffffffffffffffffffc1f7f1f000000000000000018f8ffffffff7ffffffffffbffffffffffff0ffece8033ff83810381000000830100180100818000000000000000000000
G3[51] <= 640'hffff7ffffeffffffffffffffff7fffffffffffffff3fde0000000000000000c3f0fffffffffffffffffffffffefffe7fffc0e7fecf3d8f83c300800000000000008100003881040c0000000000000080
G3[52] <= 640'hfffffffefffffffffff7ffffff7fffffefffffffff79dc8000000000000000c3fffffffffffffffffffffffffcfffefcffe0f37fcf3f8f0000c0100080001c1000030000380004000000000000000080
G3[53] <= 640'hfffffffcffffffffffbffffffffffffffffffffefffefce00000000000000006ff7fffffffdfffffffffffffe7fff7ffffffff7b84c7df7800001800e01c010080060000630000000000000000000000
G3[54] <= 640'hfffffbfeffffffffffbedffffeffff7ffffffffcfffeff00000000000000010e713fffffffffffffffffffffe7fffffffffeff7e84c7ffffff111910c00c41038c260000630020800000000000000000
G3[55] <= 640'hfffffbdfffff7fffffe6dfeffefedf7fffffffe7fffc7f000000000000003146ffe7fe7ffffff9ffff7ffee6ffff7ffffffcfffedf9c7cff1838c1fcc08630000ee20400740160000000000000000000
G3[56] <= 640'hffff77ffffffffff7ffbff3ceefe7fcffffffffefefff8060000000000000c0cffffffff738f7feffffffffffcffffff9fe71fff77ffff78f30e66c3e13000801c2070003880e3001801000000000000
G3[57] <= 640'hffffffffffffffff7ff8ffff7fe7fefffffffffffee7ffe08000000000000406ff7effffffff7fffffffffffffffffffdfffe37f77fffeff7f046618f101000083013100000062000000000000000000
G3[58] <= 640'hfffffffffffffffffeffffefffe7defbffffffffffe77fe000000000000301877ffeffe7feff7ffffffffffffffc3efff3ffc33f668f3c871c000618fc011f1c0103070080013e000000000000000004
G3[59] <= 640'hfffff9fffffffffffe9fefdff3ffc47bffffffffff7fffe000000000000001cf7ff7fffe7cfffffffffffffffffeff7ff3ffe3ff8c073e8e8c7003001c017f1c3c018f00e70024000000000000000004
G3[60] <= 640'hfffffdfffffffffffefcffffe7ff711f07ffffffff7efff0000000000000003fffe7fffedffffd9fffffffffffffef3ff37f7eff8ec7ff8eccf13b0008387fc31c20fe00ff0060c00000000000000001
G3[61] <= 640'hfffffffefffffffffffdffff7fff739ffffffffffffffef8000000000000013fffffffe7dffffd9fffffffffffffe7fffb7f3eff9cffdf1ee7ff39c38c387fe30070f0003000c0c06000000000000001
G3[62] <= 640'hfffffefeffffffffff1fffe7fcfff3fcff99fffffffffed8000000000000077fffffffffffffcddfffffffffffffe7fffffffeff9dfffcfd7ffff9ffce317f73833131004010c6000000008000000000
G3[63] <= 640'hffffeefcffffffff39f9ff3fff7ce0ff67997b77feffde990080000000008773fffffffffcfccd81ffffffffffff7ffffffff8c3bffefce13fdff97ecfe31779ff03317ce03f0e00000200c000000000
G3[64] <= 640'hfffffefefffffffffff10737fff321f99cff9fffffdfdfe40000000000003f7fff7ff7ff4dffff8fffffffffff1ffff7fff8e740ffbec73ffef33c8e6639f1e7e0d9663071c138808080000000000000
G3[65] <= 640'hfffffffffffffffffff13f70fff3615999ffbfeeffdfdfe40000000000003fffffffffffecfcfffeffffffffffffffbffefffff1ffb7cffffef1ff9e633f99fff0dde030fb7f38800080000000000000
G3[66] <= 640'hffffffffffffffffff7bf870ff73f04939f07fe6fffbff9800000000000027ffffffffffed3ffefffffffffffffcffbefeff7ef1ffb3c7f9fe78ff9eb97f8f7ff0dd7ff1ff3f0e000080000000000000
G3[67] <= 640'hfffeff7fffffffffe03fc326c7e0ccc139fb7ffffff3ff980000000000083ffffffffbffef3fcf1fffffffffffffdfbeffffffffffb7cffffef8c33f99fe8f3ffcff1ff3ff3f0c000000000000000000
G3[68] <= 640'hffffff7fffffffffff0f0f0ec71f8ec10c7f67ffffffef9800000000001c3ffffffffbfff8f8cff9ffffffffffffdff7fffcffff7fffff06ffc3007f99f8f13fff9ffff3fecf8c000000800080000020
G3[69] <= 640'hffffffffffff7fffff8e3c6ecf0f8e0c0437277ffffee7d800000000000c7ffffffffbfff9f0cfd1fffffeffffffdff7fffffffd3fffffc8ffc7ff7ff9cef1ffff9ffffffee7e0210100000000000000
G3[70] <= 640'hfffffcffffffffffffcc3cc60f1e804c04010f7fffee67e40000000000057ffffefeffff6f3fcf9bfffffffffffdf9feffffffffffbffeceffffff7ff2cf99ffff9f9ffffffff1610300000000000000
G3[71] <= 640'h7e73fcfefffff3ffffccc3860ffcc0c720f019ffffc66766000000008007ffff7ffef2ff69fe8719ffbffefffffff9fefeffff00f0b7fe9ffffee77fe6df8fffffdff9fffffe73e3e001000000000084
G3[72] <= 640'hfffffd9f8fffffff7f3e993107ffe4c3638c0efffb9cf73c000000000301ffffff7fffdfe0ef2107ffffffffffdf9ff3fffe9fd8ffbfe0fffff9fffffffef3ffcfffffb7ff9cdeff8e00000200000000
G3[73] <= 640'hfffffc8ffffffffff0f88100803e0eff780006ff7fdc7c7c00000000000fffffffffcfffffcf87f1fffffffffffffffffe7ff999cffffffffff3fffffffff3ffffffffbfffcf7800f800000000000000
G3[74] <= 640'hfeffbe837ffffffff3f88100801efcff7e008b737fce3c7c00000000001ffffffeefef7ffffece3ffffffffffffdfbfe3c5bf9198efffffffffffffffffff3fffffffffff3ff79007000002000000000
G3[75] <= 640'hfeffbf897bffffff3f9f0000001ef43fcf011b63ffefc3fc00000000019fffffffffff7ffefece3ffffffffffffffbfeff73f831cfffe7ffff7ffffffffffffffffffffff7fffffc3fc0612000000000
G3[76] <= 640'hffffff9e71fffffff89c2000000f0707c400198fffffc3fc00000000010ffffffffffffeffffcef9fffffefffffffffffff7fff1fbfffffffffffffffffcffff7ffffffefffdfeff8fe0712000000000
G3[77] <= 640'hffffffbef1ffffffe398c000000002cfbc00008fffff7efc00000000100ffffffffff9ffffffc03bffff7ffffffffff7ffe7fff07b7f7fffffeffffffffcffffffffffffff78defccef0302000000000
G3[78] <= 640'hffdfffbfffffffffc39800000000603e1e00303f7fff7ef8000000001837fffffffff03fffffc01fffffffff7fffffff7ffefffe7f7ffeffffffffffffffffffffffffffff71feffcff81c0000000000
G3[79] <= 640'hffdfffdffffffffffd813e0000086038c0007e7ff3fffff8000000000036defffffef0f8fef3e0303fff6fffffff7bff7ffef6ee1fffe3ffff7fffffffffffffdffffffff9f37fff77f81c0200000000
G3[80] <= 640'hfffff0f77ffffffffc980000a0010600180107efefbf7fde000000000123ffffffefcf7ffefff040fffffefffffffef7dffffce6ffff7ffffffff7fffeffffeffffffffffffffc73ff99f08000000000
G3[81] <= 640'h3fffffffffffffffc79d0000000080000000017e66fffffc000000000007ffffffeff07fffffe000fffffffffffffe7fffffff6f7fff7fffffffff7ffffffffffffffffffffffefffff9f00000000000
G3[82] <= 640'hffffff7f9fcfff7ee78f00000000c0808008003f70ffffff00000000080fffffff7fffffffffc0001fffffffffff7fffffffff9f7fffffff7ffffffffffffffffffffffffffffffcc7f9f00000000000
G3[83] <= 640'hff7ffc7f9bcffffffc0f0000a00001808003000371ffffffc0000000008fffffff7f7fbffffcc00000ffffffffffffffffffffd9ffffffff7ffff7fffffffffffffffffffffffffefff9ff3000000000
G3[84] <= 640'hffff7f7fb9ffffef3e3c0000200001800003000163fffff8e0000001018ffffffffff8bffffc80001f7ffffffffffffffffffff9deffffffffffe7ffffffffffffffffffffffffffff9f7f3000000000
G3[85] <= 640'hffffffff7b7fffffc230c0004000000000000018637ffff8e0000000830fff7ffffdfdffffc300000f7ffffffffffffffffffffffeffffffffff3f8fffffffffffffff7fffffffff7fffff0000000000
G3[86] <= 640'hfffffcffffffffffe020c000000000000038000c00671ffec0000000013f9ffffffdffffffc00000007fffffffffffffffffffffffffdfffffff3cfcffffffffffffff7ffffffffffff9ff0000000000
G3[87] <= 640'hff7f3f7feeffffff7e0300001c0000800000008704661b3cc00000003c37cffefefdff7ffffc010000baf7fffffffffffffffffffbfedffffffee3ffffffffffffffeffffffffffffff8ff0c00000000
G3[88] <= 640'h9cfffe7cefffffff001100fce0001000010c0000818efc7cc0000000998fe7fffffef8fff3e000e0033f7fffffffffffffffffffdffffffffffee78ffffffffffffff1e3fffffefffff7676010000000
G3[89] <= 640'h9fe77fe3ffffffffe010000000000000001c0000890c3ff9c00000009dfffbff3cfeff0fb6c00000103ffefffffffffffffffffffffffffffffff0c63fffffffffffe3ffffffffffffff662100000000
G3[90] <= 640'hffcfffe3fffffffefc0800000c0000000078000081007efb78000000bf7f1fffffffff0f96c0001ec83fffffff3fffe3ffffffffffffffffffff7c803fffffffffffff3cfffffffefffeee2300000000
G3[91] <= 640'hfffffe3fcffffffefc0c01f83c1800000030000000007e7f7e008000ff7e1fffe3ffff0f9280001e671e9f7ee01fffc03fffffffffffffffffffc700ffffffff7fff3e3cff7ffffffffcceff00000000
G3[92] <= 640'hfbff7f3eeffffeffcc0c01fffc1800000321000000010f7eff0000007fff99ffefffff07b30000cf000efdfff01fffcc1ffffffeffffffffffffc0000fffffffffff1eff7f7fffffffffdefe00000000
G3[93] <= 640'h77ff7fdf7fffffffcc8003fffe00000007c3000000017ffeff0000007ffec0ffffffff07338000cf000effe7f01cffd883fffffffffeffffffff880007ffffffc7ffc3ff3ff9fffffffffffc00000000
G3[94] <= 640'he77bfeff7dffffffcc4003ffff66000066ff80000000ffffff0000007f7e67cf3cf8ffff32c0001fc0000fff0000ff0001ffffffffffffffffff9c0003ffffff87ffcf6083f1fffffffcfdec00000000
G3[95] <= 640'hf67ffefffbfffff0cc0017ffff660c007effc9800018ff7ff800000067ffe6effff83fce12c0003f808166ff1c00c00100ffff7ffffffbffffff780000fffffffce3fe7183f33fedfffff9ce00000000
G3[96] <= 640'hdecffef39ffffffc70003ffffff1003fe7ffe20000337fff7c010001ffffc0889ff38f79008160ffe0034d389901000080ffffffffffff7ffffe4000013fffffefff7f0030f3e7fffefffc8600000000
G3[97] <= 640'hffc7fffffffffffff0003fcff7ff001ffffff70100b3fffffc0180211fff07c78f7087398181013fe0004101f800000001ffffffffffffffffff4600033fffffffffff0000ffe6fffffffffc00000000
G3[98] <= 640'hffffff3ffffffff3f0007f87007f31ffff3fff8700b3feffff00c07b3fff07cf9f00011f8380017ee08000016000000001fffffffffffffffffe06f0069ffffffffffc008c7ffefffffff3fc00000000
G3[99] <= 640'he7ffff9ffffffff3f1007f80003f7ffffccfff8400b3fffeff000eff7fffc0cf1c00008f1800017ef001100006001e03003fffffffff1ffffffe0698069ffffffffffc00803f3d7ffffff3fc00000000
G3[100] <= 640'he7efffdffffffff90f007f00008f7ffffcc7ffcc0032fffeff008effffff06f81800008e1800000ff00010000603ff87c81fffdffffefffffffe00904099feffc7fffc000038397fffffffff80000000
G3[101] <= 640'h7eeffffffffffff81e017f0001cf7feff803fdfc00163ffffff1c0ffffffc01080000007010004eff88310180007ffcfd00ffffffffefeff7ffe90800018defd1cc31e000038337ffffffeff80000000
G3[102] <= 640'hfffffffffffffff91801fe00000f7fe78003f97800073bffffffc07fffffe00000000400010000fff8c71238003fffef9007fffffffffeff3ffff8008000ffd918c000000000636ffffffefe80000000
G3[103] <= 640'hff79ef7ffffffef13800fe00001f7ff30087f92100077bffffff007ffffd0600090680001818603f98f81f00663fffeffb03ffffffe7ffdf3f9ffc600001ff19800000000000666fffffcffc00000000
G3[104] <= 640'hffcffbffffff9f708001ee000007fbf33027ffc600037ff8ffff71fcfff8000800039f010004183f98ccfe3f937ff3ba7f03ffffffff7fc74dfffc00800046e000000084010cf1cffffff20f00000000
G3[105] <= 640'hfffffddfffffff2080093e00001ffff31003ffc6000cfffffffff3fffff900020000fc0000009800f87dfeffbefff3fff603fffffeff7fe0fdfffe00008027000000000003007fefffffb20f00000000
G3[106] <= 640'hfffffeffffffee60b08d3c80001efffe8001ffe6000cfefffffff3ffefff010080003f8000309863f9fcffffbeffc77ff7c37fff7eff7f73fffffe030c00030c01e0000003000fffffff960f00000000
G3[107] <= 640'hffff9fffffffee803044dc80001efffe0011ffff0001fffffffffffeeff80000811f1fc000308037fbef3fffbfffe619ffc17fff7efffd3f4ffffe801c80000001c0000000e30fffffffbed800000000
G3[108] <= 640'hfff7ff7fffff7e003244cc80080fdfff0001ffff9801773fffff7f7feff80003191ffff8800cce3bfff01fffbfffe61c9fc07ffffffffdf94ffffe801c0000008680200000c387ffffffbff003100000
G3[109] <= 640'hff7ffb7ffffffe8032413ec00003bffb01c03f7f99002307ffff7fffffe021021fffffff820e7e3fffe31fffeffe620ec3e07fffffffffff7dfffe01108300008eff60000083c3ffffffb6f803800000
G3[110] <= 640'hffffffff7fffcc8002013ec02003fff309803c7f99000077ffffffffffe000029fffffffbefffefffe0307ffeffc4666f1f07fffffffffcf7cfffe01000700000fff40000001ffffffffb3fc01800000
G3[111] <= 640'hffffffffcfffc880020936f0a83f7ee00d80f07f99008063fffffffffde00036fffffffffefbfefffe10037fbdc006a01110077efff7ffc00cff7098011c22017fff40010103fffefffef31f00180000
G3[112] <= 640'hffffff79fffff80010033fef803f7f811880019fe7d80103f7fcfe57ff700003dffffffffffff3fff8101cff7e8f06080c787bfff3ffff79df7ff1001f41180077f7d805001fffffffffff7f1c980000
G3[113] <= 640'hfffffffefffff80000037fffc03ff7f10198011bf6e9000bffffffffffc00097fffffffffffef3fdf81003ffffc000a04df8317fffffbf7ddffff00008c983807fe7000003fffffffffffffff8800000
G3[114] <= 640'hffffffcefbfff00204007fffc07efff0011c003bffc100199fffffffffc0009ffffe7ffe800771f8fa0003ffe3e0190041f8000ffffffbfdffcff8003fcc8bc1ffff001813fffffbfffffecee0810000
G3[115] <= 640'hffffffceffffc0020600ffff00fffffe117e1081bec100189fffff7fffe00037f8ec71ce001370fce80003e3e000790005f880027efff9fdfffffc003fccfc03ffffc01cfbffffffffffeeece3000000
G3[116] <= 640'hfefffffcffffc0000400bfff30fffffe007610817f3d0001bffffffb7fe00033ff04e0c60018007f49002601800040802f788000ffffbffdfefffc000f79f807fffec0137ffffeffffffeef8c7000000
G3[117] <= 640'hffffff78cfffc00000001fff7f7ffeff017612037fbc6001ffff7fff7ff000b2f366cfe604180103e08003c0000145000f7c8000fffffefffffffc004f7dc2077efe0023ffffffdfffffff7b07000000
G3[118] <= 640'hfeffff210fffc00000001ffd7fffffff307f9310fdecf001fefffffffff801fff062f3e004f80000e3c803e000027fe00ff800013fcffeffeffffc1007ed4207ffff8107ffffffdfffffffff00400000
G3[119] <= 640'hfffffc013fffc000001c1bfc33f3ff7ff03f93f91fefff006efffffefff801dfe060f37007fc000043f982c000047f8f7e388301ffcfe7f96f9ef8c600c87c8cffdf800f5d7fffff7fffffcf00c00000
G3[120] <= 640'hfffffe600f7fc60000033ffde3f9ffffb01981b817fffe00fffeffffffe0007e6080fd03363f8800017f20c00027ffcf3ef8090037cffffffeff7f0fc01000c3fffe841ffff9fff9fffffef8c7c88000
G3[121] <= 640'h7eff7e0006ff810200087feffcffe7ff10001f0021ffc7e33fffffff7ff00cfce0feeff0277f80001fff078000673fc7fef8fc0037fffffffffffcfff400000efffe021ffbfbff9bffffffffc38c0000
G3[122] <= 640'hff7ffe0006ff98300c0ce7effcf363fff003ffcfd13fc0003ffffefffefc0fe8e0bccffc07ffc0013fe78380122ffe07fb7ffc0013ffffffffbffcfffc1c008ffffc037fffff7ebfffffff9f000c0200
G3[123] <= 640'h7f7ff30007ff800000007fedc77f3ffff023fbde2fff03c03f7ffefffffc0ff9e01ce9080ffff1817fffc0c61e07f917fffffc0013ffffffffffffffff3e0003ff8003fffd66fcffffffff9900004000
G3[124] <= 640'hc6ff078007ff80800001fffcc63ff80f00f0bffea000037ffffffffffffe00ff608fc083ffffffb9ffffc0079a260717ffbfe88041bfffffffffffffffff0001ff800cffff66ffffdfffffff00204000
G3[125] <= 640'h3efe3f2002ffc0000100e3fd6c1e8007f839feff60031e7fff1ffffffffe01ff7c870003ffc7de3fffe3c00692fe3c53ffffe5014017fffffffffffffef9e0c0e0000fffffefe7cffffffff980300000
G3[126] <= 640'h7ffc782002ffe0000008c3ff6e1f8380f80b767f2a000cffff19ffffffff83fffc0010c6ee011efffff3c006927ff8c0fff3ef0ffc17feffffffffffff79eec000009ffff7ffff0fffffff98c0000000
G3[127] <= 640'hf1f0072007fc003000007ffeedfff9fe7dc17409ea0083f7fff1bffe7ffb81cffc80c3cfee001ff97f7fc006831c81e0ffb7fd7f7d103efffffffff1f7ffffc08000bfc777dffeceffffff9fe10c1800
G3[128] <= 640'h38660461011ac9040000008f7fe2f571dce0f11f4a01337fff4ecffffefe80fd99e0127ecc003fdf7effe080367e2900ff7fff7ecf861aff97ff7fffdffffbf880063fffdeffe6fc3fffffe779c02000
G3[129] <= 640'he30006e040b3d8000000803ffc60ffb9b961c018ef8080e7ffefffffffff800df8e0833ff0000fff7effc20e326600900efffffccf8099fffffffffffffffff8c00fff9f0fde7ffffffffffffbc02000
G3[130] <= 640'hc00060800d635a010007c07b9f707e9b71f1c0000f8c00e7ffc7ffffffff800f07e0023f70000fffffffc08c0226003007fffe3887c403fffffff7ffff7ffffe87fffffde7cffbfffefffeffffc02080
G3[131] <= 640'h600567e9000003807b9f707e103339ee000e06813fffe7ffff7fff8077660800ff700007f3ff7f80f0037f84b2077ffe18007e031bbfffffffffffffff02fffffcfbfff9ffff7efffeffc02080
G3[132] <= 640'h1000002007ef90000001c3fc0717c80031b7eaf69c001fcffffeffffff980f3e0dc3f7ecc0007e1ffff0430137605f7073fc41800bf3f9933ff7fffffffffffff7ffffff9fffffffffefffe3c800000
G3[133] <= 640'h71c00000007e78010030011f60017a80068178eff9c003f1ffffef7ffff909f3009ffd77cc0017e07eff7c301200113e8ccfc000003effc023ff7fffffffffffffffffff3cffffffffffffff3c801008
G3[134] <= 640'h7f600010309d78010300019f330173b00080f9e73f800703ffffffffff791f30389ffdf3e0001ee0180020c010003ffe8c8e1800008f1fe403fffffffffffffffffffffefffffeffffffffff8c801800
G3[135] <= 640'h37fc0d1028b6009e00020ff600812b0008081001d42c010ffff7fffff391e103ffffffbf1001ee000040081404067f2073d3c00038000fec23e7adfffff7fffffffff7ffffffefffff7ffffc7801900
G3[136] <= 640'h8786c18c1ca4808ec6e63c83d8e269200031010000016112dfffea1e8f886c003ffff7e378007fc00406280200183ef90ec0fe0019876019e0318efffffffffffdfffbffffbfffffe7fffff7b9e00400
G3[137] <= 640'h9ef9f14ff886800e3ee7f81cffe6f84080e01000013dc00207ffee8fc1807fc03fffff78788c76c0060020020000fef006e3fe0001fff4c1f000c08fffffffffffffffffff7ffffffffffffef9e08000
G3[138] <= 640'h1effdaffe00600a33ec7f33c7ffffc00808e003001a7cf4803ff040170007e8033fffe197c8cf700000000024001fee003e7fe6107ffde60f700000fffffffffffffffffffffffffdffffffef901c000
G3[139] <= 640'h87befee3e00004637fe77fff6ffffc00060e001001377c7c213b110038003e0033fcf8003e99ff0080e00013c001ff008707ffe106ffdb07f7f880073fffffffbf7fffffffeffffffffffffe3f0fc000
G3[140] <= 640'h83fdeeeffce204e79fff7ff37fffe60000c000050036e47d00ff01003000d60033fe80003e9bfe00000000138000ff018783ff8020fff107fffc00013ffffffffffcf3fffffffffffdffffff3f070e00
G3[141] <= 640'h37fffe7ffcc007fc3efdfe7ffffffc00003000000082ffffe03000800101f30332f800003f72906200014013800718010083ff8031fff027dff038011fffffffff7f5ffffffdfffffffffff7f6390f00
G3[142] <= 640'hb77fff7ffe0407393df9feffffff3d600019800000821ffff00000000003f307b21000003b77906200004003900700000083fd8019ff677fffe0300107fffffffffffffffffdfffffffffffff6f8ce00
G3[143] <= 640'h8375eaefff8103b9f19bcfdeff7ffb6000389808c0069ffff0006108008f6e803738000833d9f422000040029840f10c0307fde019ffdcfffff0c100077fffffefffeefffffeffffcffefffe77f8d400
G3[144] <= 640'h1df97ff67c102fbdf271f7f7b3fe770000e30a2010536cfc00040018100af008360040101fc822939002007e0007e80f1a73864a67f9ffedf9901003ffffffffbfffffffff9ff7ffffefef7ff98030c
G3[145] <= 640'hf3ffffffffb100df1806d9ffe3ffe7c0030ff0810081021ffc0200010022bf80fee106000160060df00000020e0606001c80b2c187f83ffedf9900007fffffffffffffffffff1f1ef97fffffffc1380c
G3[146] <= 640'h80febfffff10038c1802f8ffc7ffffc0004792c00019001ffc0000180000be803a93000000003eedf13ec0823c0400001c00e00103e07efc8f80000076ffffffffffffffffffff8c983ffffffec338c0
G3[147] <= 640'h7f3fff7f004188810221c7feffff9e0063876000e1401ffc800280c000be000310801000603ffcff7ff9b3f8010007c006090703873f0003c0000020fffffffffffffffffffc8c88c0dbfff7fcc0f1
G3[148] <= 640'h801efffefea000810100310fffffff9e0063b2678107c03fff001283cf10bc0017109f318004277ffffffbffb90106e0e026c96f01c01fc800010000017ffeffffffffffffffff708c00f9ffff7cc3f1
G3[149] <= 640'h801e7ffcff30012100006108f3ffffce000132768007c03fff0012073c103c001006dfe380006373f1ffffffff18cef179feddff607c1ff0000100000131fef7ffff7fffffffff200000f17f7efe3e71
G3[150] <= 640'h7ffef901030000006000f3fffff6000413700074c03f7c801207fc017d60010fe0c1000023fff00e9ffffe9effff7fbf16ffe03e0fe008c0000001387ffffffffffffffffc00000023ffffe73c30
G3[151] <= 640'h7dfe990240000100c401fc87ff7ce18c310702e6ca3fff80077f771f3d81080804180000037819061feffe9ffeffef9bdfff620007ff1802000080307ffffffffffeffff0c00000003ff63fec008
G3[152] <= 640'h18a21ff9c7cc9810010031847fcfffe1e0121ec4dcdc30cfffe666effb1f390101874580008001ffc48083997fffff7f7fccfefff0801fe30100000001000ecfffffffffffffe0600020047fffffde03
G3[153] <= 640'h81601f39fcc818100000101877c1ff77f093fff8dec1001fffe066c7fcc7746680006c80000000fe840018bb6fffffffffedffff7fe01fff80000000000039ffffffffffffff300000000177fffec7f0
G3[154] <= 640'h83008f19fec02410000101197f8fffff3192ffff1fc1001ffff006e7fce1f4ef80306800012400ff8400083ffffff3fffffdffff7ef18e3fe0000000000171ffffffffffffff2000000001f7fffec7f0
G3[155] <= 640'h1880808383406600000001997f9fffff713fff1f3f0081e7cf7f06ffdf389feeff0168000086e47fce928067fffffbff7fffff7ee6ff8f01fef000000001e13fffffffffffffe001000001fffffecf0f
G3[156] <= 640'h1cc080c7010066000000809c6ff9ffefc3bffffc200a8177ff7be7ffdf389efee08040600086c77ffff287f7ffcf1fffffb7fcffe5ffdfc01cffe0000000861fffffffffffffc0010000193ffffffe1f
G3[157] <= 640'h1983000410006602030000bcc7f1ffe3c2933ffec000003ffff9e7f99c6383c3fc0c41208103077fffb23ef7c18407ffffb39cff7f7ffff81e9ff00000008c3fffffffffffffc0000000193fffff7efe
G3[158] <= 640'h9b27800000000783cec0017ec7f3fff380b3f33fcc8000bffff9c0733ce183cfff7c4538c100877ffcb2379e802020fdffb319ffbffefff81f9ff000000004ffffffffffffff0000000100fffffffef8
G3[159] <= 640'h18f0c010c0000f8bfc1801661c73fff3003ee1ffce000167ffffbe4391f8338cfeff6d39737e9f7ff8f0239e00307007cf82193f9e8ffec003dfff80000100ffffffffffffff00200000009bfffedfff
G3[160] <= 640'hcf8502100001983ffe4003003b8dffc0203393ffbc00014dfbf7f0e67b800667ffef8b80f3f1ffc62e79cfc0200f01fc9803ffeeeecff0031fff7690000006387fffffffffc000c0000000fffff1f73
G3[161] <= 640'h87f8000001000183fffe833083fefffc0018e3f7dfc0001507fffc666e9218067ffffff9fcfe1f1f77f18ff93f00f01f7b817cffbf0f3f7003fffffd40000077e7fffeffff8e0000000008ff0ffff971
G3[162] <= 640'hc7b8000001000099ffe6800081eff3f8403cc3e3dfe000153ffffd737f9f1c007ffffffbffff7f0f193901f016c0f00f7fd11fff77f7beff0ffcffbfe6c0003efffffeffffdc000000000023fffff830
G3[163] <= 640'h6e1b4c0000000080ffc60080004ffffc0001c3e0dff00015ffbfd9f37f3fc49d3effffffffffffc0991101700080784ff3f33ffb7efbfec31e701f9ffff000183ffffffffffc008000000103fffffb10
G3[164] <= 640'h7e83480100000000ffc6800000ffffff102307087ff000148ffff8ffff3ee3991cffffdfff7ffc069880017c0000200f67f73ffffe7fffff3fe01c93ffff00013fffff7fff1f0000000000f11fffff18
G3[165] <= 640'h67810880010100001fff000000efffef00380c0027e000148ffff99ffff6fb999ffffefffb7ffc04fcc001fe4c30010fffffffffff70fffeff780893ffff00013fff7fffff00000000000031ffffffc8
G3[166] <= 640'he3900880010000803ffe0c00026fffefc0100000070000948ffde71ffff7fe71df7f7efffbffffc06c66007f6ffc019fffffffff79030ff7ff780091ffffc0011ffffffffec0000000000007f0fff6cc
G3[167] <= 640'h62bfdc5c980082807ffe8000027dbcef81010000060081c6017ee63bfffffe739f7ffffbffbdf80004a6001fefff19ff7f7ffeffe100413ff3e000101dfce0000ffffefffe8180000000051c7ffff6ce
G3[168] <= 640'h9c6fe30000203003dff78000019f7effc1010000000000300e770499fffff9fcefffaf7ecfffee0160000083fefbff7fff3fffee000080087ec49a019fff80001dfbfffffc1800000000003e3ffffff8
G3[169] <= 640'h83fdff80006000001ffef800009bfe8fc0000001000001300067e08bbffffffcff7fbf7fcf7ef00901000003dfc3fef3efffffee0000000022c400001fffc00001fffffff800000000000001e3feffff
G3[170] <= 640'ha3cd3fcc0c900c00fcfef8000083ef83e101000000000010010fc78bfffeffffffdffde7ffd7f148400009010781b2c34fffff7c01101fe7000080001ffff00003bffffbf000000000000003f3ffffc3
G3[171] <= 640'h770f3cc61c988cc3f8ffc1000183efc1c420000000000000011f1fbffffefc3fffbffde7ff976340c000091003c0920e6fffff000038ffff8000010009fff88001fffff900000000000000037c7ffff0
G3[172] <= 640'h764fe06000bffee39fffc7600003eff882248001000004000406fcffbfff7c1f7fffd9ff6efff0c00000099871f0820e00fffe80381ffffff000800000fffcc001fffe9800000000000000073efffffc
G3[173] <= 640'hf2fde06101bf7b39bf7ffc400007ffffd84280001f300002041ec1fffffff071fbfffdffeffaf8400006019c7f708000401ffc80380f7ffff400000001fffe00001ffc88000000000000000ccfe7ff7f
G3[174] <= 640'h8279e32001277b3cf97ffe400007f3fffc4388983f90010200be87e7ffff177bfffffd1ebcbf7b404006401fff710000053ff9007e3f3ffff600c200000fff30003700000000000000010000cfffffff
G3[175] <= 640'h9a61ff0c0066ffffffefffe1000671fbf0a3891ff888080001171c7efefffe3f89efe77f7cbff90801066011ffef0000817c6900c73e3fffee38800c200ffff800e000010000000002248303fc7fffff
G3[176] <= 640'hd831c322001feeffffffff80a0010ffff10001ccc732000802389ffffefffe3ffffff9f9b7ef77008011190fe77c0080008fff00e206fffefc1840016031fff880001106011100000200000f7e7ffff9
G3[177] <= 640'h1830102003ffffffffffff182000063ff800000f3fb0000000fc9f9fffffffbfffefff1fb787ff000001800fffff0000009bff007207ffffe08160006001ffff800000000000000000000081f7ffffff
G3[178] <= 640'h1800004003ffffdfffffff98008000fffc0000077efe000600fc81ff9fffffffffeffbfff383e00000009003fffc000007f3ff003007ffc7008121306000ff7f18000000000000000c000000f7ffffff
G3[179] <= 640'h8000ffffffffffffc3048000dfff400000feff1804067f83ffffefffdffefef3fff2e0000000000133fffc000000fbfef03007fe1e0000000c8000ffff1800214400020030081000017ecffff6
G3[180] <= 640'h8000000000fffff9ffffffe76c80000eff061181f9fff801077fc73ffefcfedf3bfcff3ff2e066000000003fffff400004cffef80000f81e000000068c047fffee0371e6c08200c000b200013fffff7f
G3[181] <= 640'h81000000417ffffbfffffffffc8c0007ff00031139fff80007fee7ff07fcfffefb9fffffb70106000000003fffff40030fcf1ff84000f881000000008c043fffff7ffffee000008001120080439feeff
G3[182] <= 640'h8000000000fffefffffffffef6f80007fe8003317ffff802067eeffc07fffffefb8f4effbf0004000000803fffff6003dfff9fff6000000000000000180c7ffffffffffff8000100010200c0679ffff8
G3[183] <= 640'hd001011000fffb7fffff9fe767e80007fc8009f15eff9f300c3fef3ffffbffefc1994e9ffee00c000000001c7b3f603cfff7ffff6101000100a4020018387fffc13f700fff60013c309700997cffffbf
G3[184] <= 640'hc0000000007fffff7ff3ffffe79000037f3907737f6fff9887f9df6fe7cf7f3f4633f85fff8000000002817f7fff6067fffffef884080080002080909fe07ff700000003ffc101039866ff7338feff7f
G3[185] <= 640'h3fffff7ff7bffffff80303f68002e07a2ffffc827ffdffefc473f86e03ff7ffe840800000280ff7ffff03fffffffffff0c011c007000181907ffb200002700e6c0010018e7c3ffb9ffffff
G3[186] <= 640'h1000000001ffffffffffffffffe0713ffe002e0f826ffc0b04ffffff9c000cc7e033e99de000c00000000ffffffee7fffe7ffdfff00013efe70080809ffffb200003ff003fcc03809c3f7cefbfff7ff
G3[187] <= 640'h1000000001fffffffbfffffffeec011ff6e0233f000ff7fb06ff7fff901060f7e047899ff004000000007fefeffc6feffefffcffec0f3e6ff008c0101ffffb000003ff900fec01009f9e78ef7ffffff
G3[188] <= 640'h80301000000fffffefffffffffe6c001fc060212f003c1ff9e6ff1fed8000638070800193ff04000000060ff7fffc6fffffffff7fffc1fe6ffffc78083fffff000006ff8003fd80011b9011f23fffeff
G3[189] <= 640'h1e300000060f7effcfffffffffff9800fce70003b081c3f99c7bfffec00084300700001107f04000000243ff7ffffffffffffff3fffe3fffffffc72087ffffe2000007fc001f9801109f033f7ffffeff
G3[190] <= 640'h9f3098837783fc9f4ff7feffffff9800ffe7000720f0ff0fbb7f7fffe080000006e0000003f0400004121ffffffffffeffdfffffcfffffff3effef7e9ffffff2000007ff7803c80010077f7bffffffff
G3[191] <= 640'hf030d98c7f813f9f0ff37ffffffa91009f3fc06428183c7fbbfdfffb0000008004e1000007fe00008417f47fffff7f3edf5f7ffc873ffed93eff6e67bf3fffb200000f66f8014100907e3ffe67ffffff
G3[192] <= 640'hf00e4e03ff70c40c07fedffffffbc08c3fffe13e000026e7fe3f7fff80800080073c100000f703800027ffcff7fdffff7fff67f90183fffe997ff3fffaffffcc000001f8fc1c60200e0187cfffffe7f9
G3[193] <= 640'hf07fefffffc006c547ffffffffffc48c3ffffffe0000067efffffff98300000007fe100033ff830000e2ffffffffffffffce07ffc1b81fff99fffffffffffffc000001209c09f7008081fcffdffffff9
G3[194] <= 640'hf37fe7ffffc0004143ffffffffff87189ffffffc0000c67e7ffffff91330010006ffc0003bff82c01877cfffeff7ffffffcc1ffee03006fffffffffffffffffd8c3801000003f80010987efffffffff9
G3[195] <= 640'hf237effffffc0080037fff7fffffe0009ffffffc0000c7c7fffffff93a3801f0044e4000003fbc00197d8fffc9b3fffff3801dbee002047ffffffffffffffbfffefe00000013f8800081077ffffefffb
G3[196] <= 640'hf2fffffffffc000a83ffffffe7fef0009fff3e9f00011fe7efbffbfc300c00e08e7c4000803ff60003cf63fe6913ff7ff1c0893fe002107fff5f7cff7fffd9feffe0b000007ffc000083f3fb7ffffff9
G3[197] <= 640'hf2fffff803ffd812c0ffffffff7ff3c00f3e3cc100013b7e3fff7fde83860ce7fffcc0000066633007ed21746013ffef78c0817ff0320007fffffffff3ff993efffff2008efffc000083ff7bff7ffff9
G3[198] <= 640'hffff0ff001fff8bf608fffff7e7ff1c0277c10c00001f97e7e7f3fdfb383031f7fe60000006373d8e7f800000013ffff7ce0007ffc100001fffffff3c97f9937ffffff86fffff00001013f3fff7ffffc
G3[199] <= 640'hfdfe0ff00161df9f70ff9ff7fe7ef0c823e0000101001fe7ee6732fd3c63633f7266000080235a8d7f7900000113ffff63c06067fc808001fffbf3e39c0399a2ffffffffffffc0601008fffbfffffefc
G3[200] <= 640'hf83d2160000cfffff0cffefff99ff3c01ffe81c00001ffcf909c67fcf3387fffc00e00000081f9fbfffc0080000ef7f03f000839f800c100cf8c9966f39ff087fefffffffffc3200001919fe6f7ffffe
G3[201] <= 640'hc000600000007ffff81e3ffef91907008f0001000007fe1f921e67feffcf7ffff00c000000001ffbff8000000003fff838000099fc0000008fc0d9623c8100077fe33fffff3f1280000f81ffffffffb7
G3[202] <= 640'h3d7e01f800296efc18fffb380007008fc00000808edfffb30203ffffcf7e3f7800080000001f7fff817c080001fff8000000033e00000001001b191c810000f0037f738ff89280000699fffffffff3
G3[203] <= 640'hffff83f8000100fe80f0f7006080001fe0000000fcffffb08003fffffe663ff800000000000a79e0817efc80017fe0000000031fc0000030030119c0180030e003f87b0ff0020000243c0ffffffffe
G3[204] <= 640'hffffe3f9c010017f06dff3c06080001fc08000803fffeff00001ffff7f67cfc8800000000002fbc0037fe782007e00068000003fc0000030000019c13880300000077ff0030200000018cf6fffffbe
G3[205] <= 640'hc0fffffffff03341ff670fe080000000cfc38200007f7fffba1200ffff7f67ffc4000804010c01f90007ffe383c03e00070000007fd84000780001198ee300000000033331000000000100ff2cfffff7
G3[206] <= 640'hfffb7fdffff8bfe0ffc0000001000001e7ef820000fbfffffe02809fff7fefff80001c0f233b80e000fffffff3800c0000000082fff84400fc0103769ee300000000f07b07e01000000107ff9fffff72
G3[207] <= 640'hfffc2689fffcbfe47f800000016606017fe0a10c008f7f7f7e20809f7fffff0000c1c78773f3982003fefeffff80890000000000cef8e6c08e607066cc60f000001b1fff6300100400083eff07ffffff
G3[208] <= 640'hfff9670004ff7ffc3b3000003107660e7ff87827073fff79fff08107febce08000008f8e1806c2000effffffffc00003008000001ff880607c3c39ff7c7f0000810161e3f0200c0001011cbe8bffffff
G3[209] <= 640'hfff97600001ff9fe1ff0000033ff7efe1ffe8000813ffff8df0f8003ff93e0d0000067ce9dfefc0287fffffffffc0003eeff000000ffcc70741ff0c77e38180000002027f020000000190fe69bffffff
G3[210] <= 640'hffffe000000efcff8ff0018033fffffffffc022001fffef70fcc9000ff832100003877fcc7fffcc0c7ff310380fc8003fffffec001ff8039c2f9dce3ff3878000000202698004080001807e64bffffff
G3[211] <= 640'hff7fc0000000b83f87fcfdc07ffff7ffffff020001ffff000f78e10ffe903004003c7ff867ffffc7effe0080000fc603ffffffe003fffc99c6ffffffffffff18000000008c002000000080789fffffff
G3[212] <= 640'hff7ee003f400001f83ffffffffff7eeffcff000009ffff000fffe10fcc12004100fffff867ffffc7fffe00000c01ff77e3c00fe483ffff8f9e1f7ffeffffff7c000000408cc104000001007d1cffffff
G3[213] <= 640'hfffe7803fff8000fc0ffffffffff3803fcff40000fff7c0002fffcffc803c000c043fffc67ffffffffff8010de80ffffe00003ffc0ffff8effbffffcbbffffe70004000389c1860000000983977fffff
G3[214] <= 640'hfffebc33f7ff6007f0ff7ffff03810013fff4000ffff7800017fffff88038060f83ffffefbffffffffe100ffffe0fffe6000001ff807ffc6fffffffc000fffff1f4546609180000000000383a97fffff
G3[215] <= 640'hffff883fc3fffe0078003f3ee000800000ff40037effe00c0173fffe88328042fc7ffffed9ffffffffc00e7ffffcfffe003ffc007c009c9ffffe798c000e7ffefcf746703100004100000192993fffff
G3[216] <= 640'hfffec03f00ff3f61780000066000030022ffc1267ff8012080cc3eeee01c8000cffffffff9fffffffe001ffffffe0f0003ffff801f8000fcffffe62000001fcfe73ff801c081800000000047c0a3ff0f
G3[217] <= 640'hd3ffe1ff00000fe0ff80000000018f70007f0136fffd007000001fee40030070fffffffffffffff0f8001fffc3ff0000fff08ffc0ff0000c00f06600000008fffeffef3800000000000000a98eebffef
G3[218] <= 640'h807e83f8000003e00fc080001033fff000fe0c77ff381efe00000364008301f1fffffffffffe38c000003fe30083e033ff8001fe00fec000000020000000003bffffdff1000000800000008b2debff25
G3[219] <= 640'h263e001f0001e007ffd000663ffff000ffccf5fcb81fff008000000000003fffffffffffff300000073fc00000fffffc000007e04ff8000000000000000007ffffffe304000118000002750aeaffb7
G3[220] <= 640'h7e00fff801f001fff800661ffff000ffedfdf8103ffff80000000008003fffffffffff7f2000007fff0000003fdc00000001fc0dfc000000000000000007ffffffe38400001500000077de6f7fa7
G3[221] <= 640'h187fc00fffc00ff003ffc1867ffffe0000f6feff00077fff8000000000000ffffffffffffff000f00ffff000000000000033000fc017cc0000000000000000cfffffffcc000008d210000123d6bff87
G3[222] <= 640'h1ec3004ffff80fff80fff9ffffffffc003fefe100007ffffc1c0006710003fffffffffffffe003f0fffffc0004000000007ff9c1f817ff800000000000000007ffffffecc1804850400008425a9ff5d
G3[223] <= 640'h19590c17ff3ff87fff00ffffffffff7c60ffff6800067fffc79c034671001ffffffff9fffffe03ffffffffc001e2c08e0107ffbe1fb1ffff8000000000008003e7ffffefccc10c1884020023a2c17f84
G3[224] <= 640'h7fc403fffc63f81cfbe003fffffff3ff003fff000007ffffff7ffffff7d067ffcf9e0cfffffb01fffff37fc00703f004ff1ffffe0ffc3ff18c000000000300003fffffff1006335e919180a3d9f50d69
G3[225] <= 640'hff8007fff823f800807800fffffff1ff000fff0000ffffffffffffffffc37fffcfffc1fffffc81ffffc03f8003e7ff8ffffffffe07fe1fff9c000000010300003ffffffff8063029ece100ae745ce9ee
G3[226] <= 640'hfe007ffff801f000001f003cffff71ff000ff803007ffffffffffffffffbffffcfffc13fff7c0ffffe80138000ffffdfffffffff03ff0ffffc0000000101c80007ffffffff603784910000ea57260f57
G3[227] <= 640'h6601fffff0017f10000fe0181cff00ff8067e00f037ec3c7ffffffffffffffffcfe7c33eff3c028ffc000080007fffdfffffffff03ff07fffc0000000001cc00077fffffffe0a7fcc59811eeb4a38662
G3[228] <= 640'h79cfffff000fffc1c0ff00000f800fff067c01fcfff8103ffffffffffffffffeee7833effc002c7fe000000001fffdfffffffff01ff83ffff0000000037ce00033ffffffff6ef306c18626860f6c446
G3[229] <= 640'h801cffffe000ffffff84fc80002000fff876003fffee0001ffffffffffffffffdc7f081cffc00fc7ff000000000ffffffffffffe00ff83fbfff00081007fff0003fffffffff6e77ba9080a986a1c8426
G3[230] <= 640'h1ffffd0000ffffffc03f800000003ff830007fffe000000ef3ffffff9fb9f8fcbf00083fe01fe1ff0000000003fffffffffffe00ff83fffffc03fe00ffffe001ffffffffff36adda980f0c7e6d94d5
G3[231] <= 640'h76cfffff00003fffffe01f0e0000001f1c2003ffffc000000021fc00ff8319009c99000107784f38fc0000000001fffffffffffe007f03fffffc0ffe83fffff800ffffffffff36359dc40bc62dc9ba9f
G3[232] <= 640'hff7ffffe80000ffffbc00fc080000007fb00077fff00000000200100b80000000638010080000ff0380000000007ffffffffffff03ff01fffffe1dff07fffffc003fffffffdf76d974f889406112c82c
G3[233] <= 640'hfffffffe00000ffff3e000fe81800007ff801ffc3800c000000000000000000006bc000000001fc0000000000006ffffffffffff81ff01fffffe1fffffffffff007ffffffffec68896a6a838ab109a11
G3[234] <= 640'hfffffffe1800fffffffcc07fffc00001ffc43ffc0003f00000000000000000000000000000019f00000000002004ffffffffffff80ff007ffffeffffffffffff4000fffffffecea8926dbf14003ad70f
G3[235] <= 640'h1ffffffc0007fffffffee01ffff000007ffc7ff80003ff700000000000000000000000000001ff000000000000007fffffffffffc0ff807ffffeffffffffffffd803ffffffff48af08466a3c21345e92
G3[236] <= 640'h7fffffe830fc17fffede007ffff01803ff3ff000003fffc0000000800000000000003000003ff000000000080003fffffffffffc0ff807bfffee7ffffff073ff80fffffffffd4a3c6b87c9904760385
G3[237] <= 640'h8371ffdfc300831fffe0e007ffffe1c03ff3ff000001ffff000100ff00000000040037c13c07ff800000000080001fffffffffff80ff80fbffffffffffe0033ff807ffff07feccbc47d3ab36188ae687
G3[238] <= 640'h373ffffffc03fffdfc04000fffffbf01ffff80000007fff0033ffffc0007f009e707fffffffffc00000000080000ffffffffffe007f80fffffffffffe00000ffc0308fe00feadaaabe61f360c4e2e16
G3[239] <= 640'hf7fe3ffff01effdff000000ffffff80ffff82000007fff007fffffc00f7fffffffffffffffffe000000000180007feffff3ffc002f80fffffffffffe000003fc000081003eed7508ace614aa2f2e1f
G3[240] <= 640'hfeffc007fffffffffff800001e07fffc01dff00000001fff99ffff7ff03fffffffffffffffffffc007000000780003fffffcff00000f80f87ffffffffb0000838a00007055c5bdbc6a9fc79c252d2619
G3[241] <= 640'hffff8087feffffffff3800000000fffe008ef00000003fff99ff8307fcffffffffffffffffffffe000000000200001ffffffff80000fc00000ffffffe0000001ab0000d0556e8711a44a0bcbb533886c
G3[242] <= 640'hffff038ffef83fffc000000000000fff0000c00000007fff9fff0003ffff8403ffffffffffffffffc0000000000000ffffffffcc003fe000000fffff0000000029804340047b52931688db4adab9a129
G3[243] <= 640'hfff8018fffffff7fc0000000000003ffc000800000007fff9fff0003ffc10001fffffeffffffffffe0000000000000ffffffffdc003ff0000800fff000000000119243c1109a4c7ecca385492b136227
G3[244] <= 640'hfffc01ffffffff3ff00000000000003fe080000000000fffffff00007c0000003fffc0f086ffffffe00000002000000fffffffcc00fff0003ec018700000000057b3582011b54c2710ce81a595458263
G3[245] <= 640'hffffe1ffffffffe7fc0300000000001ff180000000004fffffe70000300000003fffc000021ffffff860000000000003ffffff80000ff8007fe00000077fc00001a35f40103ab5b22262e8c9dc2e09ed
G3[246] <= 640'hfffffffffffffff7f80300000000001ff1fc00000000ffff798000040000000007ff8000000ffffff863002000000001ffffff80000ffffffff000017ffffc00052346f4016811092c21870b884d4bca
G3[247] <= 640'hfffffffffffffffcf00080000000000ff1fe80310000ffe0000000460000000003ff9c000007fffff863083104000001ffffff00000ffffffff83003ffffffc30163dd4da3611caccd2168e8469c5204
G3[248] <= 640'h790fffffffffe7fe8000000001c0003ffffff3c3c0fffc00000000fb00000000007f80800003ffffff8c0004f8000000ffffffc00001ffff1f7fff3fffffffe833a20489a23f9d2b8ca142817c0c981c
G3[249] <= 640'h11c7ffffffff87ffc80000000104003ffffff3ff07fbe003c00000ff00000000001c00d64001fffffffe801ff8000000ffffff8c0000ffff1f01fffffffffff9304be6406105f827a206b605e80262cb
G3[250] <= 640'hc0f13ffffffffffc0001000039003fffffffffdfe000fffc0003ffc0001007f0000fffe0000effffffc03ffc000001ff03fffe00001fff1fc3ffff7e03f1b8d09e0735000fed880a93f3c390ea8c53
G3[251] <= 640'h11ffffffffffe3000000070003fffffffffff0007fffff023ffc0003dffff001fffe000000f8003003ffe000001ff01fffc00000ffffffffff80000000d25cd9c45c0fab4d91a707ec282c5a468
G3[252] <= 640'h1800077ffffffffffe70000070003fffffffff9c0ffffffffc37ffe4007fffffe13ffff000f800000000fffe000003fe01fffec00000fffffffea0000000071d90e81629d040a330ec61f00e2984e6
G3[253] <= 640'hc03ffffffffffef0000011003fffffffe0803ffffffffc7ffffc007ffffffffffffffffc00001e00fffc000003fc00fffff88000fffffff0000000000ba224743b240472a0d6367dc8327c0828
G3[254] <= 640'h17ffffffffcc000001fc01ffffff1c0817fffe07fffffffff607ffffffffffffffffe60003f00ffff000c1fe000007ffffc001ffef00000000001afaf87bc1c659b7c591295a10000723c66
G3[255] <= 640'h10000000007fffffffc800003fef03fffffe1c0047fffe03fffffffff60fffff0fffffffffffff10079001fffe0ffffc000003ffffe000c3c00000000000326a20a11e0ee906d66a3c125439c2a81b7
G3[256] <= 640'h17f7ffff8c4c01ffff803ffff7c001c3fffe01ffefffffee0ffffc17ffffffffeffff8000003ffffffffff800000ff7ff81003c000800c03098be1417ce146a0a0aac9f0a0cf54489a2f3
G3[257] <= 640'hc00000033ffffcc0007ffffc003fff38001e0fffe007feffffffffffffc01ffef8ff003fffff3c837ffffffef800000003ffffc0000001fffffcc00076d6dd0a32b00f4a71819d4596272f1cb3
G3[258] <= 640'h3ef8000000000007fffffe07ffffffc003ff0000074fffc083ffffff9ffffff9001ff800000007ffffff8ffffff81ff80000000ffffe6000003fffffffc000c2446fb78b4f1720c267129e27014238c5
G3[259] <= 640'h1ffc0000001000c3c7ffff3ffeffffff800000000100fe0003ffffcf1fffffe0000ff000000000000003ffffffe007f8005c603ffffe2400007fffffffe0005ca1646ebfcfd19d2284004a840319a89b
G3[260] <= 640'hfe000e0f0300003c01cffffffffe0ffcc00001fc001fe0000ffff86ffffffc00007f000000000000000fbffe000310003ffe03ffffe0000007ffffffff80073cfe6b29a6f1f60258c03434e99110000
G3[261] <= 640'h7e000c7fc63b801e00037fffffe001fffc13ffff8017e00007fff80ffffff800003f0000000000007ff380000003f2107fff003bbff800000ffffffffff008a9be732d9aa22267e46808e668824954d
G3[262] <= 640'h3c0000ffe03fec07e0001fffff80001ffffffffff007e00007fff000fffff000000800000000000ffff80000001ffffe3fffc80007fcc00f3ffffffffffc171001472c1667a410341120246121fc09f
G3[263] <= 640'h1cff1ffffe1fe001fabff8780067ffffffffc03f00017ff00000fff800000000000018e001ffff7000001ffffff0fffff8003fffffffffe3ffffffe21395de6a8e99a7c036c1c6c55617292204
G3[264] <= 640'h200000ffffc3ffff07fff0033f01fff800fffffffff80e0000fff8000007c0000000c000001ff0f0ffffc00001ffffffc33ffffefc0c7e80e000000081806ae316e9411f762c17a22976a74c8326c31e
G3[265] <= 640'h33c000fffffc3ffd03fff8c300007ffe000fffffffffcf8000fff800000300000000c000007fffffffffc100380ffffff83fffffffc00000000000000000a383e1e9c335ef16a5064a6cce6a28086113
G3[266] <= 640'h3ffc0ffffff800000ffffe30000ffffc00000003fffffc000fff800000100000000000001ffffffffffe3e018003fff0c7ffffffffc003c0000c7c0000071e63c503d391c6c6231609042a00581a1ea
G3[267] <= 640'h7fffffff07fd71017fffe00ec0ffffff8000003ff87f80803ff000000000180000000001fffffffffffff8017f7ffe07ffffffffffc3fee0f103c0000066430eb6950a417034f2a6f072ace4389200
G3[268] <= 640'hfc1fffff4000fffffffcff001e01ffffffc000003ff00080801f80000000001e8000000003ffffffffffffff83fffff40ffffffffffffffc00e01c000800d71c9f8c6311416e7289856041d279b021b5
G3[269] <= 640'h3f83ffff0000000ffffff8001c1fffffffe0000039000000801f80000000003fe000000003ffffffffffffffff7fffe67a38fffffffffffe07803f18e10000caa73081096b9168270f36b9c8eaaf44f4
G3[270] <= 640'h3fe01fff00000000e7ffe0007fffffffffff000030000000800f0000000000fffc00000007ffffffffffffffff3fffcf4000ff0fafffffff1ff0ffffe100d401303c5b9bcb47cdac545c0c9f72b92708
G3[271] <= 640'h3ff80ffffd000000018000001fffffffffffc100000100c0000f0000000000fffd00000007ffffffffffffffff3ffe9f8400709fbfffffffffffc7ff3e789bf98b8fdad3e5f3617fa3059589a0413246
G3[272] <= 640'hfff07fffa8000000000000010fffffffffffd57100000370801f80000000001fe00000001fffffffffffaaff7ff8e3fe00000600ffffffffffffffffffffad101d2e3c43ad97036cd7ab001814404398
G3[273] <= 640'hf7f01ffff8000000000000073ffffffffffffff900000070000f80000000003ff70000001fffffffffff00e000f0ffff0000000000ffffffffffffffffffac36170f2851467dba244f2124c1498d89ad
G3[274] <= 640'hfff81ffff00000000000000fffffffffffffffffc000000000070000000000ffff8000001ffffffffff800000001c1ff0000000000ffffffffffffffffff486edb1364813a6c4588b40e187a7e9822c2
G3[275] <= 640'hfff87fff0000001c80030f3fffffffffffffffffe000000000077800000000f8cfe000001fffffffffe00000000070ff0000000000ffffffffffffffffff3df626348fc3441f60e76596155479885338
G3[276] <= 640'hc101fffe0000003ff8d7fffffffffffffffffffff80000000003f800000000005fff00003ffffffffff800000000389800000000000ffffffffffffffffefce252dd09809888422edc9b0069e887b426
G3[277] <= 640'h3ffe800000017ffcfffffffffffffffffffffffc0000000103f8000000000003ff001ffffffffffff0000000000120000000000000fffffffffffffffe35baf5dbf188b221f13a4431d8068ed73606
G3[278] <= 640'hfffff00000001ffffffffffffffffffffffffffffe0400000783e00000000000000740fffffffffffff0000000000100000000000000ffffffffffffffffe6a675b91a5a9df8a15d9d8a1731846e9371
G3[279] <= 640'hffffc000000018fffffffffffffffffffffffffffe8e00000fc3e100000000000000e0ffffffffffffe00000000000000000000000007ffffffffffffffe8d99b6c9ee442fa40dc3a54ffde23704d054
G3[280] <= 640'he0000000000107fffffffffffffffffffffffffffe1fc00000e3f338000000000061ffffffffffffffff000000000000f80000000000ffffffffffffffb4e68e1df6a635b19e9d61c7f8daa048012213
G3[281] <= 640'h107fffffffffffffffffffffffffffe3fe00000e3f110000000000021ffffffffffffffff000000000000f800000000003ffffffffffffffd2ec48e7ffc3ae425ef6da638c586848074a9
G3[282] <= 640'h3ffffffffffffffffffffffffffffe7ff00003f1f800000000000001ffffffffffffffff000000000001f800000000001fffffffffffffcaf864e962155d5a12822b01acc205a8247cc1
G3[283] <= 640'h3ffffffffffffffffffffffffffffffff80003f1fc0000000000000cffffffffffffffff000080000007f800000000000fffffffffffff8c55ab9f541c283be085c811ece0ccc8a5162c
G3[284] <= 640'h187ffffffffffffffffffffffffffffffffe0000f0ff0000000000001fffffffffffffffff0000e00c0087fc00000000000003ffffffffffa822123ab9056159b99713e32019426546ba71
G3[285] <= 640'h800000000000fffffffffffffffffffffffffffffffff0000070ff0000000000000effffffffffffffff8000e01c0001ff00000000000003ffffffffff8beba984a3badcf970badc960b848b025383dc
G3[286] <= 640'he00000000001fffffffffffffffffffffffffffffbff00000000f10000000000008effffffffffffffffc000409c83007c80000000000003fffffffffff787c92b8393ac182fea042b4b424f91520106
G3[287] <= 640'hf00000000003fffffffffffffffffffffffffff773ff00000000e0000000000001c6fffffffffffffffff8000099c738fcc0000000000103ffffffffffd188248d69c699fb598c41743eba81eeb1a31e
G3[288] <= 640'h310000000000ffffffffffffffffffffffffffffffff0000008480000000000000c7fffffffffffffffffe00f8dc0f3f3fe3e000000300c7fffffffffecad757405d24d89698bdab064590591ed0a350
G3[289] <= 640'h8000c0000000ffffffffffffffffffffffffffffffff000000070000000000000086fffffffffffffffdffe0ffff0ffffcf7f800000340cfffffffffffa5c2c0ef02d9d03b7ff73136a73696d6c010f7
G3[290] <= 640'hf000f80000f0ffffffffffffffffffffffffffff07ff0c0000000000000000000004ffffffffffffffc0fc00fffbfffff8e7ff0000030ffffffffffffeadd309ad8fbea14b120a543e9096176f69ebc3
G3[291] <= 640'hf081ff0003f87fffffffffffffffffffffffffff03f08e00186000000000000003cfffffffffffffff00fc003ff3fffffcfffffeff07ffffffffffffff6e33811091a048656ff11803aa8272869bf684
G3[292] <= 640'hf8c3ff0007fc7fffffffffffffffffffffffffff83008000080000000000000003e7fffffffffffffc00f0000fffffffffffffffffffffffffffffffffcdd3b68c9250680ad1139ac1d0496aa67196b6
G3[293] <= 640'hfcc3ffff0fffffffffffffffffffffffffffffffc0000000000000000000000001c3fffffffffffffc0000001ffffffffffffffffffffffffffffffffefc62d6c20051cdba8b37da87128dfc04b805c0
G3[294] <= 640'hffffffff1ffffffffffffffffffffffffffffffff80000000080000000000000007ffffffffffffffffa00001e1e7fffffffffffffffffff1fffffffc070809d960aecc481e72dbe87d04123f368204e
G3[295] <= 640'hffffffff1ffffffffffffffffffffffffffffffff80000000000000000000000007fffffffffffffffff00000e9e1fffffffffffffffff7c07ffffffc1f35e0571e0e81ebd9ae771801876ffc658f017
G3[296] <= 640'hfffffffffffffffffffffffffffffffffffffffff8000000000000000000070077fffffffffffffffc7c0000843e03ffffffffffffffff821e96ffc0000eb20cabb4914963e8a02a474ee5777b91c7de
G3[297] <= 640'hfffffffffffffffffffffffffffffffffffffffffc0000000000000000000807ffffffffffffffffffff00808800013fffffff7fffffc4108012c080008a3f4db68d1a10b3cb14c4d5f5f83e76c944c4
G3[298] <= 640'hffffffffffffffffffffffffffffffffffffffffff000000000000000000317fffffffffffffffffffffffe7ce00000fffffff3ff00f80080000000000d686841a2b8d7801323ad33f0d993d31f09709
G3[299] <= 640'hffffffffffffffffffffffffffffffffffffffffffc00000000000000000183ebfffffffffffffffffffffffff820007ffffff1f800000168200000000a27d9d93956432fdd3464a23a2c995de102f4f
G3[300] <= 640'hfffffffffffffffffffffffffffffffffffffffffff8000000000000000090e1f97ffffff00ffffffffffffffffff0fffffff03f00000f01800000800043d3be3666540e50a1d8e4f2446854ec0c265a
G3[301] <= 640'hfff3ffffffffffffffffffffffffffffffffffeffffc00000000000000002a71e77ffffff11fff1fffffffffffffffffffffc00700001fc6c00000e000626e99123f53a406d16212632fb718b031be08
G3[302] <= 640'h7ef3fffffffffffffffffffffffffffffffffffffffc000000010000000036d979ffffffff1f001f3fffffffffffffffffff80000000ff0ae40c0bb803d7e91c4208e24e152b20c8648cf74892011922
G3[303] <= 640'h18c1ffffffffffffffffffffffffffffffffffeffffc00000001008107ff774f8357ffffff3e00ff3ffffffffffffffffffd00000000ffb8a404ff3fffbff4d3b8b2eaa1b7adc2c38056340542e93139
G3[304] <= 640'hff811fffffffffffffffffffffffffffffffffffffff80000000fee09ffedd23c7b9ffffffff3c1ffffffffffffeff67fff97fb200036fba2e6ebe7ffe515a62f4805d005fcc417920799218b4cc4566
G3[305] <= 640'h701ffffffffffffffffffffffffffffffffffff800000e0fff09fc422275dbafffbff1e07e00fffff3ffffff9fefff87ff000007f63143a00077c52eb9a9c305302182844b503ff403d8ca4d142
G3[306] <= 640'hff81ffffffffffffffffffffffffffffffffffffffffe0000001fff07fe569a6209dfff3ff7f07f803fffff9ffff7fffffffffb2c000010ec9b86f807bf37305301fb1e35a0fb32240401ad006d944af
G3[307] <= 640'hff81ffffffffffffffffffffffffffffffffffffffffff000007ff007ed1c66c98617efffffe87ff00ff8099fffffffffcfe376ffcfc1a2074d67ec05de5e46aa463102f5b99108341b35149e708383f
G3[308] <= 640'hffe7fffffffffffffffffffffffffffffffffffffffffffc000fff01c84d4f0193ca3cbffffffaff07ffff01fffdff0180e01c4fe0f8189f2779063fdcb105c64140594384ced0b621ab059e29f82526
G3[309] <= 640'hffe7fffffffffffffffffffffffffffffffffffffffffffe0007c17f213e0ee6b3ee07fbffffffff0000f8fffff000cc0003fa5b9c0f0235efd4063c3adf2ec32a640211e0e589012367746afed8c8d6
G3[310] <= 640'hffe7fffffffffffffffffffffffffffffffffffffffffffe0001000040f4541210f20028ffffffffc00000c001041ceeff20feff8f3effdfd7378001380c7cb0df888807087e988e0046b9869ab811a0
G3[311] <= 640'hffe7ffffffffffffffffffffffffffffffffffffffffffff00000000a46f6ec9002cc7707fe00000fc188300f80000778380787c41ff4f8823d6eec7dce1e0a454683e67b84c43ce419a8522df8d3ccd
G3[312] <= 640'h83007f3fffffffffffffffffffffffffffffffffffffffff000000000c85f97001796d9463ef3f0ff503be7608000007ff601f75c1e523c669b37bffd10c03ad658b7d21e85de30b6373d824b7901b23
G3[313] <= 640'h3c1f00ffffffffffffffffffffff7ffffffffffff0ffffff8000000006fb0733fffdc19af31cf80fa00ecfe4ffc7000081fa0089c127423061b9c3ff4bf40c652fc1bc033a323ffac27be82db694b1b6
G3[314] <= 640'h7f01fffffffffffffffffffffffcffffffffff000000ff00c07f0f0c04bffffc3ea57174f07ff8fff901ffd101800115b8118105c3dfeedd980356de503bcf82b8c2c26ae0cf44863a147416c4b6
G3[315] <= 640'hc10000077f007ffffffffffffffffcf8000000030cf00f03ffffc01f107de73fc11ff9f8082ae63984c0fde1ff9d00001f07575ec0c2836433a0220028afc5829a4997b04c5ca652fb959eae1ef3782a
G3[316] <= 640'h507fffffffffffffff0000073ff00fffffff007fffffffeff800fffe7e47e3e113283801807698fbdc1cff31f8001fdf83fee043288aece08a007619e1b5f3e44cf6025cde4a0b0b84b1576c44c2
G3[317] <= 640'h80e0fffff0000ffff800000007fff07ff0ffff001ff00000ff3000e3ff71c090300080047d7e59659d7ae07e7ffffe0007f7e6cfe05bf517f31bae8071baba9e8b17240080ea90f34b362d893cb82008
G3[318] <= 640'hff3fff00000000003fff00000003fff8000000fffcfffffff000077fffff000c8fc66002bbc19671a1fad1bf7feefec0c79efeff04f0127b96d1f080f2d9679eb1d936c18f8de25cf20e448538b60809
G3[319] <= 640'h9c00ffe0000fff0007ffffffffffffffffffffffffffffffffc00033fffffe01fb9e10018300c68829481a1ffffeffdfffffe1be048af8a8b653b4806940cf25925b065847ccbd6f6938aa30b5a25116
G3[320] <= 640'hfffffff0000007ff00fffc7fffffffffffffffffffffffffffc0003fe7ffff01e80043ffe60022069f2000639efffffffffee1234b63937747b097c8398ea71d95284b0381243cc5c03ee10a05aa2699
G3[321] <= 640'h1fff001fc03fff1fffffffffffffffffffffffe00001fffffe0008007cf83fc0030620e3feb027fffffeffcfc0a39175562eaf0d05ec7fedec4159c2e232064a53fd889204f4dbe848ce
G3[322] <= 640'h3fff000f00c0ff3fffffffffffffffffffffff000001fcfffc000c80ff08b9e00007fe0000013feefffffffc66d39eaf048192151bfc251417a4c3baa000951013a4c5b71354fbfe9a90
G3[323] <= 640'h1f00000707e0ffffdf5fff7ffffffffffffffe000003fe1ffc000c80ffc001fe0003e280c792002e1c7efffd666be815f509faf9af707f534142c33892c904485a845800e1a55090aac5
G3[324] <= 640'h3c00080001f003ffc7ffffffffd30000007ff3fff0000000fe31006c0f06f8fffb33803b93fff0f60cb8f69a4bc6f7681e53dd05af6fcd62e38f9802353d5415f2ee6da44b7
G3[325] <= 640'h8001ff93fff3fd5d000000001ffffffc00000effc6083dff17f47ffff0019be07fcf0f1c9ef3508eb762a544cc7fe2a6f5400d81c7e891824c2044de968f6a8b6
G3[326] <= 640'h100000000000000000000000000000001f81f5414ffd000000000fffffff80000807efff84efc2062fe300101603c00ff7e7546a8f69b20650415ae46aa9ea019fa1ca508083ac20c166cf736155a
G3[327] <= 640'hf3ffffff0000000000000000000000000000f91f5cc0ffe0f800000003fffffffc0000000300f9f9f83f03000619e0fcffc06514d46e9bee3ff88f21de580012b051324222252c9fdc84f95473802b04
G3[328] <= 640'hfdfffef000f080f8011f7cffffc7ffffffffffffffffbf3eff3ffffff000fffff8037fffffe07ff821c37be700f9c0d3f9806ea841712030558b4db667a95d1cd2cf332c665825de0035f00e7346108f
G3[329] <= 640'he0fffffeffff00000f1f010f00000000ffffffffffffff3fff000000f003ffe7fff0c00000007ff8703f830004003c6507c00fa15844c6360b19dc6e543cdf0568284e1e25117df84813322fca7e7dae
G3[330] <= 640'h9fffe1ff000000fff800ffe0000000ff0000ff0f0300ffffffff007fff009fffffffffe0fcffff3f870ffe0000ccfc339f800354fdc1499cbbf834378120f2cc7e8621000a7221820803af293d3ac070
G3[331] <= 640'h26f01000000100ffffff8000007fffffffffff0fe02fffe10006ffffc01c3fffffe00000ff8000f6ffffe30007cf000361fe2357227c803524a4c4e659b5721971722418b189db70c89c245300f83aaa
G3[332] <= 640'h6c03fffffffc000c000000078005500ffffff000040ffe0000fffff81ffc000000000c3d000007ffffefffe88f84000e1ff03593649d6d1686ef302fcada7c33e54ed310d36079488c024bb80485757
G3[333] <= 640'hfe2600c7fffffffffffffffcffc3fffffffffffe0000fc810070ffffffffffffff000100000000000380010831001effdfff5ac868f8d3cab077f9e7a217c829bd2707bf83d142d12061b7be86d87446
G3[334] <= 640'he106c00000008000000000000001ffffffffff1ffffffffffff0fff078ff00fffff8c0e0f0007000040000017f1ffcfeffff40086639ca0e2b26a06a86898e603840ed540e6592ad0505369aa6784a4d
G3[335] <= 640'h7c25be00000000000000000000001fffffffffffffffffffffffff3fffffffffffffffffff7ffff81c000819fffeffff9bfec5aea498ee5724894538a16af8160e824b8c066fdf3a0c6070c838ba1cd0
G3[336] <= 640'hbb8f997fc00083c000000000000005fffffffffffffffffffffffc07ffffffffffffff00fffffeff9c9f01967fffefffffb65b00d5a6388a926b362123144718aa48590662dee00512400d9f8d1c0889
G3[337] <= 640'hbbff002fff8007c000000000000003fffffffffffffffffffffffeffffffffffffffff00ffffffff80fe0c089efff7fffefe0ead02afd2ef1c078b072c48b250213f1c0b70920c18a90d9be1e92e290b
G3[338] <= 640'h7f007fd3ffc31c0300000000000001ffffffffffffffffffffffffffffffffffffffb3000333fbfffe807ff03ff8b00efc48e6d208d8aee05d6a911b3d639308a805010a44674908912423aad00711a3
G3[339] <= 640'hb3c07f08f7c03c03e0000000000000fffffffffffffffffffffffffffffffeffffff03000007c7ff303ffffffffc100003406f007bb5e3a81f64d37730f9d881dd6400c2ab5919f608330073dcea3170
G3[340] <= 640'h72feedf1ff300000f0000000000000fffffffffffffffffffffffffffffff8f080000000008ff11f380070ef87ffb08400857a18623ee762a24c71d06d6fcea8c5514ea499a4564b72752e89f7d207c7
G3[341] <= 640'hb3ffea9ffe7c8100f80000000000007ffffffffffffffffffffffffffffff80000000000001f890001000001cfcf8001fc85d047fd5df2024499c90434cd21b514a00db8a14e2045ac7febaf3a86491f
G3[342] <= 640'h14fe619ffcfe0000fe0000000000003ffffffffffffffffffffffffffef0000000000000000870008380001f7a40319f877d39183aa2d2ba7ee386275252a7b8a41b2e631edc09846250c50e18c44b49
G3[343] <= 640'h34ff6017fff0001e3d0000000000001ffffffffffffffffffffffffef8000000000000000000000303000ff4ffb00e6cea7a362ff7cd1ff01d7a13eb08fa7dae6069dc415c1009a69e4c3b6a7d710d02
G3[344] <= 640'h1ffe0e8ffff771fff00000000000000fffffffffffffffffffffefc7c000000d2a0054919d04a1123240b06661a904776ebf4cfc767be1650f135e5919b330bf82304600137003781272bb276690f3f
G3[345] <= 640'h1fff038ffffffffff00000000000001fffffffffffffffffffffff000fef30024bee61c0faa853152c4f920ff61ff40306df196d494bb0432a688ca18bac6e7764563b980101b4ec8279b0f024036f7
G3[346] <= 640'h82fff0787fffffffff00000000000cffffffffffffffffffffffffffff0090f85c78da0945594a8fa3ec17f00181bffff74af8f0d282384336d82de0a2297cb1468c60bd5c5824f3b81808e4af4c2854
G3[347] <= 640'h31e363f9010377ffff000000000008ffffffffffffffffffffffff7c38672a8146aed15559e216367799f2f80364a1fffee647e340335716cd92ec6dd2321e4f5bd8f610401408d2031567332122a402
G3[348] <= 640'h43c30006e7fe827fff80000000000000fffffffffffffffffffffefb1903d18027bd197970044a408dd740c1e07aa3fbefe8a81ae88e201dcf41fa31b8f1483c52dac3c0446c08530980906241b61a16
G3[349] <= 640'h41fe3f980000781ffffc000000000000ff3ffffffffffffffffffffbfc53de0518977f5b2ee782c089ec01df807c39d6400001e0216c90738025fa77d67b95bdd3780924c454059a2c8820602e729d41
G3[350] <= 640'h3fffffcc080181fffffc000000000000003fffffffffffffffffff90587ff3b489741eca0730e0f808ede30007fd7e845c43092362310ebc97bebe6e4b9d553baf4cc44052a45c01e8c00116fe03c0e
G3[351] <= 640'h1bffffdc0380f00fffffc0000000000000005ffffffffffffffffcd3f9301e79053d9f62878946e0044401c0003f99f3c86d8c4d0923a0d6e90dacf7e040d1c58868132805931a6072012027a01a0b95
G3[352] <= 640'hefffffcc0016005e7ff8c660001000003c1f0f11ffffffffffff018c1d1ffd84bbccc7e1782c180d5141200086f801989f30700b9bea12dd11be0a78347fdd51d7b0c9046931c0020c3d149a9466895
G3[353] <= 640'h7ffffffc000ffc07ffffff0810000001df87ffffffbfffffdff80007de0867e4655075030b748fef859dc710799c40e2066af83e26bc1e071af060426fe68e1759e0f6c2481a4c5730ec126d502149d
G3[354] <= 640'h7ffffefff00003cc0fef3ffe1018fff860578863fff0ec47fff8000ffffdf2c45c348b6a0e1871cd322e96003631a367fc872d2fa72b2c9742d4444f515962652740cdc2d8b14c45fc24ab439a2022a
G3[355] <= 640'h7ffffffffff380343e1f800f8f88ff7c9007cdc1ffe008260000ffcfe81c99d50037b11289d9dd98c8a40c7cc74f1f843d8fe97527755364be958c77405ba315064661a26a5290e1000010533d4632c
G3[356] <= 640'h1ffffffffffcc0385ef89f07f6fd07f5af00787fffe000c08c3feff8e0101c86cb1e2626b0f3e1e0ab75bf9f8bef006824f1370d6c708c142a8e69b144d6141aaa70830a200081e48416105c7110c48
G3[357] <= 640'h5ffffffffffce03ffc60a1fffde387f3f88bc390e04000129c01c030600013b7eeae09ae4fd0b524c33223f80a7cc01e2f5ee477c8ddb6b8108c9d8a629a2e431b468cb046004c2640104120c843942
G3[358] <= 640'h1dffffffffffcffc3f81fe1998e300006ec65fe690000000163000e000038016d6a8e31f02bc08a53bedfa00c0f65ffffdf333f05102501dcb6bbf325927a839a6b88c1b460a025cc4305003640e3da1
G3[359] <= 640'h5f97ffffffffffefbffe65a9d99afffe0f801fdd7200000bdf801ff01993ed95f0b87be3aa6104a9179a10f80ac5f7ffdc8d6fff88be0ebd077389262fc551f04155000000e042c0154323183a21997
G3[360] <= 640'h3ff37b7fffeffffffe3ffff1f7fff1d3fffffff7f0b063fef8c83ecfd2e7db8f294c60279174c984f89f1de45bb3bfffd3b57b76bbbea2dddb19e0b238a169040491a090a71c8101808d700f6e4010e
G3[361] <= 640'h631c5651effffffffffffe2ffffffefbffffffb7f37350fdf033bfcf018f0043ab0d8e3b30dcdc20800ebfc7eb3bffffe79d45680ae435e7978ce14d4864836c732a4000c0010901c00928030440144
G3[362] <= 640'h855001a71b7bfffffffffffffffffff76efffff1107eadfffc0f7f010e7e7007af744ef60506ddbf114b6600faecfd7fffd87c02d52cd33565928d19cc6bc20e023aec865030d8950e32a4c601405e29
G3[363] <= 640'h1c8207723f7fffffffffffffffffff502dffffc70ff0f2c1fc0fee256d070c23b6ef8a01f8da77f54b3c20e1dae93cafff546291611bf66848f202c3c151a340b9c8da13ab90e6180c3c461533ed1204
G3[364] <= 640'h960422317ffffffffffffffeffffff5014ffffffe0183dc0811ff884e3870015172a24b41ebe2dd7df8015e6dcafcf8f1f816f0941b797e22c622e8ceae8b30a210224de04217649912c485b00227308
G3[365] <= 640'h6138084ff87ffffffe7ffffffc13fd0630f03fffc0041ff961bfbf1935f4f71f8e652c18c0aa3ed1397776ef8aba78f0f57f16978585a968ff079b590d362a109b0122410312040ca4e0d4424460123
G3[366] <= 640'h401208084af3ffe09f01fff7fe0007900a0f00e37eff7fc0e0f84e2828215fa20088ec113b4c21bc02136d0ffa518b8e4b9adf838c9106c8d88be417539012d62dc823048811b960480580e281a01675
G3[367] <= 640'h8805a129a1913cfc00000f83071000d031de003fffff7fffc1be002ecc6110cd27260abdb057d4bcbda305bfc338dd4ec1347f77ba5ef183e7e1351a5c586c157101180100cc164978965ac802820061
G3[368] <= 640'h14073ffa40a425668dfc0316700f3000333ffffffffcc1b4662609af319b6caac28513cdade1feff8faca80d1ca59fe550341dd167f4a310a1e994dc2ba04c0809208030c3ff11000142d0108d
G3[369] <= 640'hf4003b23237cd91f8ff030240618000071fffffffffc048d37e60421b8f513f3187f8fed9f1bd2e8fed6ce34a0951b4b2755f272ac7c9706481eeaf1660647a68820053110594001070131048
G3[370] <= 640'h188000c8ca9113c20f0007fd01ef20007e1dffffeffcfcaef01182efb008a3dd3d745f4a8c68530bdf91119bb17f6ef2653ccf965b226da97f463744700113ca0080804b001b41a302b4421c4
G3[371] <= 640'h2208003b83c4e603000008572b5f7300fffffffec3ec42447bf454a24f5048103ccc1f251b035e8892dbc058cd19a41816f9d0e810debddae190ba800b281e73108824a047205a2419020080
G3[372] <= 640'h78040040b20172000009a32c7e6777f7ee03ffff0f655d00af03960f07c9246f20b247c28e1e4414ac81ede9d98c512a487cd33d954563503e397cb6208a72300061448313d112048b21087
G3[373] <= 640'h3c882805b158c000000bf0001b83f0c87ffffe063cc1e5f245f34fc319fab74a54eb5b6511de68859dee29e558319b10584f23fc3cebd70e2e140280022a0c0080701e82410240004770191
G3[374] <= 640'h4d380040652100000024004147c0b3f8f8fff1df78694bc05910c1039f29e172825d8332146603380ed862e282ad1f4e95fe7562df153840210445b0d01a3160070a20961a200064270688
G3[375] <= 640'h28f20000036e390000f01200dac07e1fff9f81f0337fc15aad25105883846d1af36c18851f6c80f803d5f5fac666494647484b784643eb81f3569818400121c4081f3c14325c000e22424c
G3[376] <= 640'h1c780d80002838600a580000730000f9ce812ee006ca8390b91bbb78ecfb57008f0b97a85d994dfd8a9ebca192820f242ca695ba2e0ccd0388dd9c8c01517080031c2818141500873e03c3
G3[377] <= 640'h17e321880100736fb280002000000009dffbe7997f0277b22ce085dd8956960474339a551201d7a2a46f0568f1a5664a2e6591959204600512008760aa945e0050c1e18d20c00071f01fd
G3[378] <= 640'h63c0e0b40007713b78001180801c7fe7103e01964dbc20f11ff994e53535b7614e9fccd6363bf524e2c8e6cc8204118b941e406cecd3001fcb4331a2840130048fce18c20400000c0028
G3[379] <= 640'h6631f01e4b4400121e000111080003e03ff7fffbd7b39523111cbaa64b5cd94c703a8e901aef3e0ca8ddf01c0380510519277f9c32e801b138b00b4810e1a69818c84006c180000000022
G3[380] <= 640'h2cc470326cc6002cd80000300303fc07ffffff9abd14b83ea790c0131940c92fa260465bda5ba3f0af5cec89b040201243c2d00050696b6ab09a23633841080008010030000000000422
G3[381] <= 640'h81f0e02f01e1e000340019b73fff001e6ffffffd66b1a0161c3d014117112028de68418738594e847f9a0b3400100c00586081150e668a0c1c0124420418040000200000000000010022
G3[382] <= 640'he63cc141ab18080400437a3fff3f37fffffffd216ea1ba904abd2058c3692edc8d06bbb410c34a8851d53800a513411101d15fb8e2ab4d0a006c4006409c00000000c0000000000008
G3[383] <= 640'h337f7fb3b01e8600001a32bf7f7ffefeef7ffcc54610860f9681c2130e89600a6e9961678d2f1a234005600b48040006a01852fc7162629105c11e0013090300100000820000000000
G3[384] <= 640'h6f0fc07fc7987fbf00021c7fffe3181feffe32d0bdba7089480b70f5bce80942d96d5479042936ecd2858000000003000300319a845029d84ee3480000800000000009800000000000
G3[385] <= 640'h14f907fc07ff9f9014004028ac3c1fc0f3028312ace5645411cf27d09d5a2587702cc7bd2f6eef11020c000000000000033930dc7ddb6da3e501200000000000000009800000000000
G3[386] <= 640'h50ef007e30c3f0cffac0006b4783fe6bfff4e0d2cb4eba4acf186b6a1a9a7b112e40dcc71407a8d1a200000000000000034884b1c65aef90122000000000000000009800000000000
G3[387] <= 640'h800000000000147cf000f7ffefc7e567c531ff17ffff08720763c5682d2503477437b1050d0926033d95f2d86bd07c438800000000001bc01222000aa4a0480000000000000000000000000000000
G3[388] <= 640'h503cffe30000e1e7076336a4e3fffef32cc83ead390a9d20b7021bac8453a9455304387dc70b6c180118000000000003ad9f90518630024708000000000000000000000000000000
G3[389] <= 640'h38000000000002903ffdffffc0630766383a00fc3f83ffd0541780727dd85805252443f400f0013503281d318c3100080000000000003ec2b25e57685338964000000000000000000000000000000
G3[390] <= 640'h440000000000004f000ffffc09838e593b847ce806371a019b44804bd100053d8a60110e42001a0028a47ecdf6d0000008000000000002cd33a4a670e272463000000000000000000000000000000
G3[391] <= 640'h12000000000000627f001307fe7e07fff3be2afc0650dc976bd97c3a62c5ac70a50d90a48000181746c6a22606000420000000000000004251cc9a34a258380000000000000000000000000000000
G3[392] <= 640'h960000000000000b3ff0301c0c0eef81e19f268a0040340663f3fb8dfc5bf15204409d6600003010abc8000000000000000000000000000ed9f1a850f8f0000000000000000200000000000000000
G3[393] <= 640'h420000000000000507ffeffffff07fc7b7001ad32a18400669df0fc32c35a2303c5d440000000000040000000c100000000000000000010fcbe1b844f1e0000000000000000380000000000000000
G3[394] <= 640'h3c00000000000001607ffce9ecf7c077fdc7e88d77583e60008007c80068086194eda0000000088000200000000000000000000000000b6f4be5b8545fe0300000000000000380000000000000000
G3[395] <= 640'h470037ffffffff803fcf0f40ac0003fc0000053fcf0550508080018e000001f011600000000000000008000000000beff97532741ff0700000000000000080000000000000000
G3[396] <= 640'h2ffc00187f080fff8e71f57800382803f7c00f7e1703cef1b00200043000000001400000000000000008000000001f6fe8673a781c30000000000000000000000000000000000
G3[397] <= 640'h70000000000000052f8c004037007ffe03cb859778480ff3218fdc47c76ad79143c0001000080404100000000000000000000000001b07ef672a61c000000000000000000080000000000000000
G3[398] <= 640'h700000000000000113ffeffffc0e187ffec4e6c3984001d9b1c5f17f07aa547508c70c00000000000020000000000000000000000003010533fa61e002000000000000000080000000000000000
G3[399] <= 640'h8006c7fffe1f3f82e020e19b636c052319dff81fd7f7e82fe33f081c00000040402a00000000000000000000000000301e107aaec7814000000000000000000000000000000000
G3[400] <= 640'h206041ffefc8e077c1f0bcefe05ff8f9ff81f9bf37ffa2351c0000000000000000000000000000000000000000060056522e690800000000000000001180000000000000000
G3[401] <= 640'hcc0000ffe0017f07f87f8e9681ffffffe0602c3b6cc5ab510000000000000000000000000000000000000000006037f1bf6690030000000000000000000000000000000000
G3[402] <= 640'hcf00000000001ffffe0ffeb807fffff802c2c1c70376b58000000000000000000000000000000000000000000603fb33f6680320000000000000000000000000000000000
G3[403] <= 640'h24dffc0007ffe0001fffff7200fe7ffe00122d1c3f946a78000000000000000000000000000000000000000000203ff33f4680028000000000000080000000000000000000
G3[404] <= 640'hd8fffffffff0ff0001fc71a07e77fde00193c073bf848700000000000000000000000000000000000000000001c3fb13f078086c000000000000080000000000000000000
G3[405] <= 640'h338007fffffffffff007f844143f78e00190407f1e058610000000000000000000000000000000000000000001f1e111b070746c000000000000080000000000000000000
G3[406] <= 640'ha11000f800003fc03d07ef4177cf880018068f61be5101000000000000000000000000000000000000000000118e813b870412e000000000000080000000000000000000
G3[407] <= 640'h4c00000000800006ff3fcfdc31cc80000007ffe49d5100000000000000000000000000000000000000000000818fe12f83043bf000000000000080000000000000000000
G3[408] <= 640'h137800180030f00020fffffb0960c10000c3eff8c704210000000000000000000000000000000000000000000407e1ab87906a0800000000000000000000000000000000
G3[409] <= 640'hc37fe0fff7ffff800001fef434c0c0000788ff306000100000000000000000000000000000000000000000000067919c79eb90108000000000000000000000000000000
G3[410] <= 640'h77ffffff7fdfffffff07be33c138000c8c019444000000000000000000000000000000000000000000000000067c39c79f05200c000000000000000000000000000000
G3[411] <= 640'h7c01780780000f8fffff8f96c9c4e00e0be0881800000000000000000000000000000000000000000000000007f83e07879320c3000000000000000000000000000000
G3[412] <= 640'h1f0700010000000000ffff70008ff000228011c000000000000000000000000000000000000000000000000007c00607874c4881000000000000000000000000000000
G3[413] <= 640'h618000200008000000077f2d0fe7000006e04810000000000000000000000000000000000000000000000000640000302400800000000000000000000000000000000
G3[414] <= 640'hdfc4001cfffff97fe0010ce1d80000010683560000000000000000000000000000000000000000000000000660000180127800000000000000000000000000000000
G3[415] <= 640'hc3fffffeffffffffff7b3f990000000000180a00000000000000000000000000000000000000000000000006e08800804cf900000000000000000000000000000000
G3[416] <= 640'h3e100611800000031f73ffe65450000000330000800000000000000000000000000000000000000000060006e0000003b9fc00000000000000000000000000000100
G3[417] <= 640'h97f98000807e03c0001009440100000000c030818200000000000000000000000000000000000000002000200000000ff1e00000000000000000000000000000100
G3[418] <= 640'h3a11feec000007c800006389d00000380017847220000000000000000000000000000000000000000000005c0000000200c00000000000000000000000000000000
G3[419] <= 640'hbbf000003ffeffff8cfffff40000030000600101010000000000000000000000000000000000000000000620000000000000000000000000000000000000000000
G3[420] <= 640'h4dffffe7ff0c00018c00998820003138041a48388000000000000000000000000000000000000000010084c0000000000000000000000000000000000000000000
G3[421] <= 640'h110cfe0fe000000000000097040070c08009f120000000000000000000000000000000000000001801000000000000000000000000000000000000000000000000
G3[422] <= 640'h231808000c0c0000000671285c27883708330090000000000000000000000000000000000000000010c000c000000000000000000000000000000000000000000
G3[423] <= 640'h1b3d901e000107ee1c78b1581c21e0f8c104d802000000000000000000000000000000000000000010c820fc00000000000000000000000000000000000000000
G3[424] <= 640'h417839c003ff0100010007a0033f38600017c0080000060000000000000000000000000000000004188007620000000000000000000000000000000000000800
G3[425] <= 640'h36707f037c800003000000030000c3f000807a1900000600000000000000000000000000000007e0390083cf4000000000000000000000000000000000000000
G3[426] <= 640'h5c88e000c0007000000002620000063e021f6000000000000000000000000000000000000000741390004480000000000006000000000000000000000000000
G3[427] <= 640'h2800003f80000078700000030ccfa0000206c00000000000000000000000000000000000000001911831470000c00000000a000000000000000000000000000
G3[428] <= 640'hdd9ec01e601fc000000371f80c3f65f902020000000000000000000000000000000000000000f811c382c5600c00000001a000000000000000000000000000
G3[429] <= 640'h210003f080ffc00380010c0fff1eecc60360000000000000000000000000000000000000000ec819c38701e0830000c01c6000000000000000000000000000
G3[430] <= 640'hcffe3ffff000000000121808c190427438e0000000000000000000000000000000000000007400803870641830001f8380000000000000000000000000000
G3[431] <= 640'h2fff80000030003ffe780001ec38a428c00000000000000000000000000000000000000000060000300107808000700208000000000000000000000000800
G3[432] <= 640'hd80000180000ffff800c01ca3e4780004c000000000000000000200800000000000000000200000380003800800300000000000000000000000000000000
G3[433] <= 640'h53800080183ffef880f1008005c680004c0000011000000000000700000000000000000006e0000181c7f800000100000000000000000000000000000000
G3[434] <= 640'h14c6003c83ff0c0000000724fe0027014c00001c180000000000070000000000000000000ee0000003797e00000000000000000000000000000000000000
G3[435] <= 640'h3481ffffff000001887e180000076c37c000036000000000000000018000000000000000700000000fc1e00000000000000000000000000000100000000
G3[436] <= 640'hbfffe138c000037f074000000076ff7c0200030000000000800000180000000000000005c4000030000c00000000000000000000000000000100000000
G3[437] <= 640'h3fff00000030ff13800000000077ff4c0000000000000007400000000000000000000000a0000000000000000000000000000000000000000000000000
G3[438] <= 640'ha3c0000007f81b800000000003fff4c544018000000000fc0000000000000000000000740000000000000000000000000000000000000000000000000
G3[439] <= 640'h3c0011cfff2200000000000003fff4cf52fd6000000000400000000000000000000000000000000000000000000000000000000000000000000000000
G3[440] <= 640'hf1cffffdfc000000000000017fe7cc317f8700000000000000000000000000000000000c000000000000018200000000000000000000000400000000
G3[441] <= 640'h14fffcde000000000000000033ffecc2801800000000000000000000000000000000000e0000000000000c310000000000000000000000000000e000
G3[442] <= 640'h4fc7e00000000000000000013fffee140d8000000000000000000000000000000000000000000000000080000000000000000000000000000000000
G3[443] <= 640'h426800000000000000000007ffffcff8040000000000000000000000000000000000000000000000000000000000000000000000000000000000000
G3[444] <= 640'h1ffff7cff348000000000000000000000000000000000000f0000000000800c0000000000000000000000000000000000
G3[445] <= 640'h203fff0eac000000000000000000000000000000000000000e00000000000000a000000000000000000000000000000000
G3[446] <= 640'h80800000000000002000006001c30e80000000000000000000000000000000000000000000000000000002b0b0000000000000000000000000000000
G3[447] <= 640'h2000006001c1060100000000000000000000000000000000000060000000000003ccd75af0000000000000000000000000000000
G3[448] <= 640'ha0001061468026000000000018000000300000001020000000000000000000801506690c80000000000000000000000000000000
G3[449] <= 640'h760001061640026000000000000000000a40000010080000000009200000000002f87980c00000000000000000000000000000000
G3[450] <= 640'h5b0001070000126000000000000000000860000389900000000000ec0000e005186c480000000e000000000000000000000000000
G3[451] <= 640'h800001b0000070000336000000000000000000cee0000040000000000022f8000e000602c411000000f800000000000000000000000000
G3[452] <= 640'h34009000000301803fec00000000000000000715fea0001000000000000010000006080808c0000000000000000000000000000000000
G3[453] <= 640'h38400600000020180136800000000000000000004fd2000180000000000058000000040000000000000000008000010000000000000000
G3[454] <= 640'h1400000000020000000000000000000000000071c4a4380e00000001d60c300000011000880000000000000c0000000c0c00000000400
G3[455] <= 640'h1f40000000082000000000000000000070000002bcfd0a30380bce511dfe230000000006080000003000000187fffc00fcfce3f0000e00
G3[456] <= 640'h100000011c000000000608000000200000000012b00d400fc9c520081470c678d30ab0002000001d80123cfb0ffffc6693ff6807efe6730000200
G3[457] <= 640'h1c0000000060600b0103554000150ab01000eec000edb1ef9c9e4ac80f0c42800200c9ff09ff9bbfbfffff3f6ffef3f07ef767be000000
G3[458] <= 640'h1800000000000000000078080000004060712e748a37c4cf0840000005c000107dcf0168f93b77c26642f11fdd330d843283bffeff3fe7fffff81e35679e303300
G3[459] <= 640'h2800000000000000000000000100000f780a2d660058bc088000000000000022f80f79215249fdfd835701ffd93289dffa579fffffdbe11feff80f3f3e9e303380
G3[460] <= 640'h70000000000000fe00000100000000153800000000000000000004000010003c83ff01711aa29e1393100079dd32c99fd2177fffe7c3e1fffffc0d970f9f803000
G3[461] <= 640'h4000000000000f1f80000000000000080800000000000001000000000000003eefcfff76224b901f92f84128df2ac9db8a13fdffffbff9fffffe07838c87881700
G3[462] <= 640'h14000000000000f178000003000000000000000000290380000000000000000271efee1f361997fc1914cd0187f2ec1fefe73b7ffff3ff9fffffe0083c687881460
G3[463] <= 640'h110000000000000e9f80004001000000a400800000022c14000000000000000027cffe0e61904ed67e56736c007ea6c1fafa93f7ff3cfff9ffffff80107f879823e0
G3[464] <= 640'h30000000001000100e8010136c1c00000000000008de0000000008000012115a8c2f400100000000000000000036df1d5d200055a303c86f37e1feb6c0dffa02f7fffff3f07ffbfff020fff3803160
G3[465] <= 640'h303000000000307000010333ef8200000000000000ff000000000000000040845080180000000000000000000003e0683f36000488000e1dc9548f2b5c06b429bffff3f73fcf3fbfee80233fa383100
G3[466] <= 640'h7808000008000003f9cfc3110200000000000000e000000000001000006680c39000000000000000000000000000000c00000c1e4ff299ac36862b3804146b8ffe01800fcc3f1fee4001e99c01000
G3[467] <= 640'h60400000000003c07e8610cae000000000000000c000000000001000080110021b100000000000000000000000f3b00000000000000094a1c0a0312000038cd3000000c0820104000000000000000
G3[468] <= 640'hc00008821c7e373d4afc44a0000000000000040000000400001800000104e8f40040000000000000000000010300060e800080013c1ebde1b311b00000000000000000001000c07a0039dc40200
G3[469] <= 640'h80e010008618c1c78601fa180bec00000000000000400000000000018000001184cd504000000000000000000000180178a00801418007f1601a01c2db20677cef3f3c0000fb6fc9fb060073fc040000
G3[470] <= 640'hffc000841bf0c01fff9a1c02400000000000000040000000000000800002100609b2b0000000000000000000000b80ff0000194c000008ee878f261a6637e428ff3eff039f7fef59f0017000200400
G3[471] <= 640'hfffc0c0003e0d3fffffa30348c0000000000000000800000000000080000210a1018e5a000000000000000000000807ff000189284000001f95e74e8ae31ecca9ffff3fbf0c33cc8800380028481780
G3[472] <= 640'hcfc80080b3fffffffffda112700000000000000000c000000000000800000a0a2070e4a80000000000000000000084e86c15dfaea3c0000000dc1f880e61b35905d63313d94d6e0408b08343dd41700
G3[473] <= 640'hf84bc0010fc7ffffffff84245f0000000000000000000000000000000000002842000ee1800600000000000000000684429f4f7af48000000000791ea6071c25d60e6703100495877988481429610080
G3[474] <= 640'hc0c3cf1149ffffffffff8f38600000000000000000000000000000000000002840004f70000600000000000000000df03f19c7fe30000000000001ee47a7000000003859711913c6dc017e0109200080
G3[475] <= 640'hc011feffc23fffff3ffe8998000000000000000000000000000000000000001020004cd4000000000000000000004abcfb05f6fff00000000000000182020000040002dffb07081f981eab0000000400
G3[476] <= 640'hfcc7f80025fffffcfd7f222a000000000000000000000000000000000000000040004c045e0006480000000000000c7c6604a21c000000000000000000e000021b29cc508ee902330629c06060001800
G3[477] <= 640'h7000ff1041f3fffce076e4900c000000000000000000000000000000800018001000204048000b840000000000008000000367e0000000000000000000000013c24c70cd9703220b4e0c23204e780002
G3[478] <= 640'h3808c1efc5f1ff7c7ff94991000000000000000000000000000000008000140010001fc606000d70000000000000000001009c00000000000000000000801081f01ae44b8fcc0bc3b201e1101458061b
G3[479] <= 640'h1800e17b45f8fffcfff090c20000000000000000000000000100000080000c0001000100800240f70000000000000000000060000000000000000000000487900c52df1e2b07841803242090418d0208
end
always @(posedge vga_clk) begin
R0[0] <= 640'h0
R0[1] <= 640'h0
R0[2] <= 640'h0
R0[3] <= 640'h0
R0[4] <= 640'h0
R0[5] <= 640'h0
R0[6] <= 640'h0
R0[7] <= 640'h0
R0[8] <= 640'h0
R0[9] <= 640'h0
R0[10] <= 640'h0
R0[11] <= 640'h0
R0[12] <= 640'h0
R0[13] <= 640'h0
R0[14] <= 640'h0
R0[15] <= 640'h0
R0[16] <= 640'h0
R0[17] <= 640'h0
R0[18] <= 640'h0
R0[19] <= 640'h0
R0[20] <= 640'h0
R0[21] <= 640'h0
R0[22] <= 640'h0
R0[23] <= 640'h0
R0[24] <= 640'h0
R0[25] <= 640'h0
R0[26] <= 640'h0
R0[27] <= 640'h0
R0[28] <= 640'h0
R0[29] <= 640'h0
R0[30] <= 640'h0
R0[31] <= 640'h0
R0[32] <= 640'h0
R0[33] <= 640'h0
R0[34] <= 640'h0
R0[35] <= 640'h0
R0[36] <= 640'h0
R0[37] <= 640'h0
R0[38] <= 640'h0
R0[39] <= 640'h0
R0[40] <= 640'h0
R0[41] <= 640'h0
R0[42] <= 640'h0
R0[43] <= 640'h0
R0[44] <= 640'h0
R0[45] <= 640'h0
R0[46] <= 640'h0
R0[47] <= 640'h0
R0[48] <= 640'h0
R0[49] <= 640'h0
R0[50] <= 640'h0
R0[51] <= 640'h0
R0[52] <= 640'h0
R0[53] <= 640'h0
R0[54] <= 640'h0
R0[55] <= 640'h0
R0[56] <= 640'h0
R0[57] <= 640'h0
R0[58] <= 640'h0
R0[59] <= 640'h0
R0[60] <= 640'h0
R0[61] <= 640'h0
R0[62] <= 640'h0
R0[63] <= 640'h0
R0[64] <= 640'h0
R0[65] <= 640'h0
R0[66] <= 640'h0
R0[67] <= 640'h0
R0[68] <= 640'h0
R0[69] <= 640'h0
R0[70] <= 640'h0
R0[71] <= 640'h0
R0[72] <= 640'h0
R0[73] <= 640'h0
R0[74] <= 640'h0
R0[75] <= 640'h0
R0[76] <= 640'h0
R0[77] <= 640'h0
R0[78] <= 640'h1ee000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[79] <= 640'h1fc700000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[80] <= 640'h3fff00000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[81] <= 640'h7fff00000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[82] <= 640'hfffff0000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[83] <= 640'h1fffff0000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[84] <= 640'h2000000000010000000000000000000000000000000000000000ffffc0000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[85] <= 640'hfffff0000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[86] <= 640'h100000000000000000000000000000000000000000fffffe000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[87] <= 640'h9c00000000000000000000000000000000000000000000000001fffff8000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[88] <= 640'h9cf000000000000000000000000000000000000000000000000000fffff8000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[89] <= 640'h1800000000080000000000000000000000000000000000000000ffffe7000000000000000000000000000000000001000000000000000000000000000000000000000000
R0[90] <= 640'h1003f98000000300000000000000000000000000000000000000001ffffe3800000000000000000000000000000000001000000000000000000000000000000000000000000
R0[91] <= 640'h1fffc98000000300000000000000000000000000000000000000001fffff0800000000000000000000000000000000000000000000000000000000000000000000000000000
R0[92] <= 640'h1fffe98000000000000000000000000000000000000000000f00001fffff800000000000000c000000000000000000000e10000000000000000000000000000000000000000
R0[93] <= 640'h103ffff7f000003010000000000000000000000000000000000000001fffffb60000000000000700000000000000000000067c000000000000000000000000000000000000000
R0[94] <= 640'h3ffff6f000006ff8000000000000000000000000000000000000001ffffffc00000000000007800000000000000000000f7f000000000000000000000000000000000000000
R0[95] <= 640'h3fffff6700006efe8180000000000000000000000800000380004100ffffffc000000000001ce000000000000000000000f3f800000000000000000000000000000000000000
R0[96] <= 640'h7ffffff3003fc73ee000000000000000000000000000000c300600009ffff2000001000c1fff7000000000000000000001bdf000000000000000000000000000000000000000
R0[97] <= 640'hffffffff61fffffff701000000000000000000000000708f78c000009ffff6c00000038effff70000000000000000000001f6000000000000000000000000000000000000000
R0[98] <= 640'hffffffffffffffffff8780000000000000000000000060fffce00000fffffffe003803dffffff000000000000000000000071000000000000000000000000000000000000000
R0[99] <= 640'hfffffffffffffffeffc4800000000000000000000000e3fffe200000fffffffc900399fffffffc00000000000000000000071800000000000000000000000000000000000000
R0[100] <= 640'h1fffffffffffffffffffc00000000000000000000100167ffff000000fffffffe900fd8ffffffff00000000000000000000069900000000000000000000000000000000000000
R0[101] <= 640'h1fffffffffffffffffffc0000000000000000000000033ffffff0001ffeffffff9a3efffffffffc80000000000000000001061000000000000000000000000000000000000000
R0[102] <= 640'h1ffffffffffffffffffff7000000000000000000001037fffffd0003fffffffff9f7efffffffffd00000000000000000000037000000000000000000000000000000000000000
R0[103] <= 640'h1ffffffffffffffffffffe30000000000000000001001e7ffff99c03fffffffff9fffffffffffff00000000000000000000037ee0000000000000000000000000000000000000
R0[104] <= 640'h9ffffffffffffffffffefff0000000000000000000003bfffffe0b6dfffffffffffffffffffffff000000000000000000007efe00000400004004000000000000000000000000
R0[105] <= 640'h9ffffffffffffffffffffff00000000000000000000b7fffffff816ffffffffffffffffffffffffe000000000000000000067fff0000003800000000000000000000000000000
R0[106] <= 640'hffffffffffffffffffffffe8000000000000000008037fbfffff097ffffffffffffffffffffffffe000000000000000000007ffff806173e00000000000000000000000000000
R0[107] <= 640'h46fffffffffffffffffffffc0000000000000000000033fffffff8f6ffffffffffffffffffffffffe00000000000000000001fff3fcce1fff00000000000000000000000000000
R0[108] <= 640'h65ffffffffffffffffffffff78000000000000000021b7fffffff8ffffff3fffffffffffffffffffe00000000000000000001ffffefecfffff6000000000000000000000000000
R0[109] <= 640'h457fffffffffffffffffffffe380000000000000003193fffffffffffffffffffffffffffffffffff00000000000000000001ffffffedfffffe000000000000000000000000000
R0[110] <= 640'h97ffffffffffffffffffffff718000000000000007133fffffffffffffffffffffffffffffffffff80000000000000000001fffffffffffff8000000000000000000000000000
R0[111] <= 640'h9fffffffffffffffffffffffc3f00000000000000383ffffffffffffffffffffffffffffffffffff80000000000000000001ffffefff7ffff0000000000000000000000000000
R0[112] <= 640'h37ffffffffffffffffffffffdfe600000000000002083fffffffffffffffffffffffffffffffffffc0000000000000000003fffffffff7fffc000000000000000000000000000
R0[113] <= 640'h37ffffffffffffffffffffffffee0000000000000009ffffffffffffffffffffffffffffffffffffc0000000000000000002effffffffffff0000000000000000000000000000
R0[114] <= 640'hffffffffffffffffffffffffffc000000000000018bffffffffffffffffffffffffffffffffffff80000000000000000007fffffffffffff3000000000000000000000000000
R0[115] <= 640'h20000ffffffffffffffffffffffffff00000000000000013ffffffffffffffffffffffffffffffffffff80000000000000000007fffffffffffffe000000000000000000000000000
R0[116] <= 640'h7fffffffffffffffffffffffffe0000000000000003b7fffffffffffffffffffffffffffffffffffc0000000000000000000bfffffe9fffffc000000000000000000000000000
R0[117] <= 640'h3fffffffffffffffffffffffffe00000000000000c3f7ffffffffffffffffffffffffffffffffffff0000000000000000001fffffff9fffff8000000000000000000000000000
R0[118] <= 640'hffffffffffffffffffffffffff0000000000000003ffffffffffffffffffffffffffffffffffffff00e00000000000000019ffffe7ffffffc000000000000000000000000000
R0[119] <= 640'h1e3fffffffffffffffffffffffff000000000000001fffffffffffffffffffffffffffffffffffffffffe0000000000000000003edfeffffff8000000000000000000000000000
R0[120] <= 640'h37fffffffffffffffffffffffff0000000000000038fffffffffffffffffffffffffffffffffffffddd800000000000000000003039c7fffec000000000000000000000000000
R0[121] <= 640'h1cffffffffffffffffffffffffffe00000000000001ffffffffffffffffffffffffffffffffffffffdff0000000000000000000000101ffffe0000000000000000000000000000
R0[122] <= 640'hcfffffffffffffffffffffffffc000000000000001fffffffffffffffffffffffffffffffffffffffff0000000000000000000000000fffc00000000000000000000000000000
R0[123] <= 640'hfffffffffffffffffffffffff8000000000000008ffffffffffffffffffffffffffffffffffffffffdc04000000000000000000000073e800000000000000000000000000000
R0[124] <= 640'h1ffffffffffffffffffffeb3ce0000000000000008fffffffffffffffffffffffffffffffffffffffffc0600000000000000000000001ff000000000000000000000000000000
R0[125] <= 640'hf7fffffffffffffffffffffc80000000000000000fffffffffffffffffffffffffffffffffffffffffc7e8000000000000000000000000000000000000000000000000000000
R0[126] <= 640'h8e7ffffffffffffffffffffff800000000000000007fffffffffffffffffffffffffffffffffffffffffffc000000000000000000000000000000000000000000000000000000
R0[127] <= 640'h4ffffffffffffffffffffffff7c0000000000000013fffffffffffffffffffffffffffffffffffffffffffd000000000000000000000000000000000000000000000000000000
R0[128] <= 640'h313fdffffffffffffffffffffffec00000000000003fffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000000
R0[129] <= 640'h200010fe7ffffffffffffffffffffffffb80000000000003fffffffffffffffffffffffffffffffffffffffffffff800000000000000000000000000000000000000000000000000000
R0[130] <= 640'h204030fe77ffffffffffffffffffffffff80000000000002fffffffffffffffffffffffffffffffffffffffffffffc40000000000000000000000000000000000000000000000000000
R0[131] <= 640'h4003ffe7fffffffffffffffffffffffc00000000000003fffffffffffffffffffffffffffffffffffffffffffffe40000000000000000000000000000000000000000000000000000
R0[132] <= 640'h37e7ffe7fffffffffffffffffffffff800000000000003fffffffffffffffffffffffffffffffffffffffffffffff1d00000000000000000000000000000000000000000000000000
R0[133] <= 640'h3ff7ffffffbffffffffffffffffff3e000000000000043fffffffffffffffffffffffffffffffffffffffffffffffffc0000000000000000000000000000000000000000000000000
R0[134] <= 640'h1fffff3ffffffffffffffffffffff04e0000000000004ffffffffffffffffffffffffffffffffffffffffffffffffffe4000000000000000000000000000000000000000000000000
R0[135] <= 640'h9ffff71fffffffffffffffffffffcffc6000000000000fffffffffffffffffffffffffffffffffffffffffffffffffffe800000000000000000000000000000000000000000000000
R0[136] <= 640'h8feffffefffffffffffffffffffffffee0000011c00063ffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000000000000000000000000000000000000
R0[137] <= 640'hcc080000f7ffffffffffffffffffffffffffffffc000011600067ffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000000000000000000000000000000000000
R0[138] <= 640'h200de00000277ffffffefffffffffffffffffffffffd8000fdf0076f7fffffffffffffffffffffffffffffffffffffffffffffffffffe30000000000000000000000000000000000000000000000
R0[139] <= 640'h10041c00000677fffffffffffffffffffffffffffffff8c00fee787ffffffffffffffffffffffffffffffffffffffffffffffffffffffe3c000000000000000000000000000000000000000000000
R0[140] <= 640'h4ff8c000e7bfff7ffffffffffffffffffffffffffffe00eec787fbffffffffffffffffffffffffffffffffffffffffffffffffffff7ff000000000000000000000000000000000000000000000
R0[141] <= 640'h847ffcc0033c3ffffffffffffffffffffffffffffffffe00fe2e9c7fffffffffffffffffffffffffffffffffffffffffffffffffffffffc010000000000000000000000000000000000000000000
R0[142] <= 640'h997ffe00031939ffffffffffffffffffffffffffffffff8f9f73fcffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000
R0[143] <= 640'h219efff000111119fcfffffffffffffffffffffffffffff079fe3c3fffffffffffffffffffffffffffffffffffffffffffffffffffffbf2e080000000000000000000000000000000000000000000
R0[144] <= 640'h93ffe8000c18127bfffffffffffffffffffffffffffff801773c77efffffffffffffffffffffffffffffffffffffffffffffffffffc9e9800000000000000000000000000000000000000000000
R0[145] <= 640'h23fe9000800806fdffffffffffffffffffffffffffff00363f1cfffffffffffffffffffffffffffffffffffffffffffffffffffefc898000000000000000000000000000000000000000000000
R0[146] <= 640'h37e0000000002f8fffffffffffffffffffffffffffc80b67fbc7ffffffffffffffffffffffffffffffffffffffffffffffffffc00010000000000000000000000000000000000000000000000
R0[147] <= 640'h660000000002f3effffffffffffffffffffffffffe80bffeff37ffffffffffffffffffbffffffffffffffffffffffffffffffe00010000000000000000000000000000000000000000000000
R0[148] <= 640'h2000000000003107ffffffffffffffffffffffffff0017cfff3fffffffffffffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000000
R0[149] <= 640'h61001fffffffffffffffffffffffff80b60ffe3dfffffffffffffffffff3c1feffffffffffffffffffffffffff80000000000000000000000000000000000000000000000000
R0[150] <= 640'h40001ffffffffffffffffffffffffc80173ffc1bffffffffffffffffffffc0049fffffffffffffffffffffffff00000000000000000000000000000000000000000000000000
R0[151] <= 640'hfffffffffffffffffffffffff8017ffe71ffffffffffffffffffff800061ffffffffeffffffffffffffff0e000000000000000000000000000000010000980000000000
R0[152] <= 640'h7ffefffffffffffffffffffffc046c7f93f7fffffffffffffffffff80008399fffffffffffffffffffff3c1000000000000000000000000000000663870c00000000000
R0[153] <= 640'h37fffffffffffffffffffffffe066c7bc07ffffffffffffffffffff800008fffffffffffffffffffffff000000000000000000000000000000000670060f00000000000
R0[154] <= 640'h3ff6fffffffffffffffffff8f6006c39c01b7ffffffffffffffffff8000003ffffffffffffffffffffff800c00000000000000000000000000000010040700000000000
R0[155] <= 640'h6fe0cfffffffffffffffffe872102f38c309bffffffffffffffffff8080807fffffffffffffffffffe7fc00f80000000000000000000000000000110004640000000000
R0[156] <= 640'h3f0c3fffffffffffffffff8601c770803098bfffffffffffffffff8c9003fffffffffffffffffffd73fe0000000000000000000000000000000001000c600000000000
R0[157] <= 640'h8003f0c3fffffffffffffffffcc00c37008018281fffffffffffffffffc0206ffffffffffffffffffff3fff00000fe000000000000000000000000001800ce00000000000
R0[158] <= 640'h7e0d1fffffffffffffffff9c8000010080008099fffffffffffffff80027ffffffffffffff9ffffffc7e00000fe000000000000000000000000000c00ce00000000000
R0[159] <= 640'h1e091fffffffffffffffff1e810001001800801ffffffffffffffff0b023bffffffffffff239fffe867c800089ff808000000000000000000000248004f80000000000
R0[160] <= 640'hf2087ffffffffffffffff3817260407980004263ffffffffffefc60c18dfffffffffffff07fffbcc03e00207fffffe7e00000000000000000000c0001400000000000
R0[161] <= 640'h672087ffffffffffffffffffb0e00066900000363fffffffffff0f60708ffffffffffffff9ffffbf033f0003fffffffffe00000000000000000000001b400000000000
R0[162] <= 640'h470c07ffffffffffffffffff9280003e9200003431feffffffff0f013003fffffffffffffbfffff3c1be0007ffffffffff000000000000000000000009600000000000
R0[163] <= 640'hf0c07fffffffffffffffff81780003f1e00000000fffffffffe800010017fffffffffffff3ffffef0fe810e7fffffffff000000000000000000000100700000000000
R0[164] <= 640'h4c0007fffffffffffffffff9b6d000ff1e01100001ff7fff7ffc049800017ffffffffffffffffffe3ff78018ffffffffff000000000000000000000000600000000000
R0[165] <= 640'h410106ffffffffffffffffffbe800cfbe2200000037c7fff7ffc00988001f7ffffffffffffffffff7fff7ce3ffffffffff800000000000000000000026c00000000000
R0[166] <= 640'h6ffffffffffffffffffbf0008f9c2380080003cffffffff8004040007fffffffffffffffffffffffeeffffffffffffc0000000000000000000026808000000000
R0[167] <= 640'h6fffffffffffffffffffe60191f36cc00800007dffffff8000406001efffffffffffffffffffffffffffffffffffffc40000000000000000000061c0000000000
R0[168] <= 640'h3ffffffffffffffffffe0018b73ff80001883e7ccfbfe40140000080feffffffffffffffffffffffffffffffffffe30c00000000000000000010000000000000
R0[169] <= 640'h13ffffffeffffffffffffc001307f830000c3b76f8ffae001000000019fe7fffffffffffffffffffffffffffffffff30c00000000000000000000000000000000
R0[170] <= 640'h3efefffffffffffffff90001307ff10004813767ff97e000000000010387ffe7fffffffffffffffffffffffffffffe0000000000000000000000000000000000
R0[171] <= 640'h3ffffffffffffffffff80c181207f80103087ee0ff9763400000010001e0927ffffffffffffffffffffffffffffffee000000000000000000000000000000000
R0[172] <= 640'h2fdb7ffffffffffffffc001802072000311d7ee76ff2e040000001000070801e6ffffffffffffffffffffffffffffff000000000000000000000000000000000
R0[173] <= 640'h7397ffff0fffffffffc80c3873fe00020c3fffee1f8f840000000000130000045ffffffffffffffffffffffffffffff80000000000000000000000000000000
R0[174] <= 640'h39c7fffe67ffffffff00081863fe00003c1fff8f8bb3900000000000300000005ffffffffffffffffffffffffffffffc0000000000000000000000000000000
R0[175] <= 640'hfdff7e30f7ffffffff10000803960030ffdbfff6cb3f90800000001c3c2000001ffffffffffffffffffffffffffffffc0000064000000000000000000000000
R0[176] <= 640'h6fffff33ffffffffff00001c082c01b9ffbffffb283200000010003673c0000008fffffffffffffffffffffffffffffc12146b9000000000000000000000000
R0[177] <= 640'h7fffff8e0cffffffff800010496f01bbffdffffb200600000000001678c0000009fffffffffffffffffffffffffffffd8c0ffff800000000000000000000000
R0[178] <= 640'h3fffffec30ffffffff800000ebe791ffffffffff0000000000080017fe0000003fffffffffffffffffffffffffffffffcceffffc00000000000000000000000
R0[179] <= 640'hffffff0308ffffffe000000cbf308fffffffe7e080000000000001fff8000000ffffffffffffffffffffffffffffffffffffffe08000000000000000000000
R0[180] <= 640'h100ffffff7000efffffc0000700330c8ffffffff6e000000000000003f91e000004fffffffffffffffffffffffffffffffffffffff98000000000000000000000
R0[181] <= 640'h100fffffee0017ffffffc000000338e8fffffffff9200000000000003e3e740010fffffffffffffffffffffffffffffffffffffffff8000000000000000000000
R0[182] <= 640'h17fffffc0017ffffffc006000b7ffffffffff7fb60000000000c0007ff84001dfffffffffffffffffffffffffffffffffffffffffe400000000000000000000
R0[183] <= 640'h37fffff80407effffef0200019effff7ffffbfef0000000000000007f1e4038ffffffffffffffffffffffffffffffffffffffffffe400000000000000000000
R0[184] <= 640'he7fffe90000ffffffe8806607bcfffffffffcff2000000000289737fff6067ffffffffffffffffffffffffffffffffffffffffffe700000000000000000000
R0[185] <= 640'h9ffffff8000003ffffe800046ffffffffffffff7c000000000298b37ffff03fffffffffffffffffffffffffffffffffffffffffffff00000000000000000000
R0[186] <= 640'hffffff0000007fffff0100cffffffffffffffffc000000000238fe7eefee7fffffffffffffffffffffffffffffffffffffffffffffe0000000000000000000
R0[187] <= 640'hf9fffc0000003ffffb0119ffffffffffffffffff000000000027fefeffc6fefffffffffffffffffffffffffffffffffffffffffffff0000000000000000000
R0[188] <= 640'h3f9fffc00000007ffb3e011ffffffffffffffffffc000000092e3fe7fffcffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000
R0[189] <= 640'h33dfffc0000000f7ff06013fffffffffffffffffec0000006b6ffff7ffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000
R0[190] <= 640'h1cfbf8000000046ff20607ffffffffffffffffff00000006b7bffffffffffefffffffffffffffffffffffffffffffffffffffffffff8000000000000000000
R0[191] <= 640'hc3b3980000000e6ef724ceffffffffffffffffffc000000ebffdffffffff7ffffffffefffffc7ffffffffffffffffffffffffffffff9000000000000000000
R0[192] <= 640'h1ec00000000083e6c007ffffffffffffffffff7000000737ffdff7fdffff7fffffffff9fffff7fe7fffffffffffffffffffffffff0000000000000000000
R0[193] <= 640'h198018ffffffffffffffffffffff800001f7fffffffffffffffffffff7fe7ffffffecfffffffffffffffffffffffff000000000000000000
R0[194] <= 640'h180018fffffffffffffffffffffe808019fffffffffffffffffffffff1f48effffffe7fffffffffffffffffffffffc000000000000000000
R0[195] <= 640'h1901cfefffffffffffffffffff900219fffffffffffffffffffffff822ce7ffffffefffffffffffffffffffffff8800000000000000000
R0[196] <= 640'h1000000017fffffffffffffffffffffb2399fffffffffffffffffffffffff2278ffbfcf7cfffffffffffffffffffffffe000000000000000000
R0[197] <= 640'h1077ffffffffffffffffffffe339dfffffffffffffffffffffffff323167ffdefff1fbfffffffffffffffffffc000000000000000000
R0[198] <= 640'h6007fc00000000000000000000000000000000000000000000fffffffffffffffffffffff3fbffffffffffffffffffffffffff980003fffffff3fffffffffffffffffffff8000000000000000000
R0[199] <= 640'h201e003fc0c0000000000000000000000000000000000000000016feffefeffffffffffffffffdfffffffffffffffffffffffffff83c001fffbf3e3fc7ffffffffffffffffffe600000000000000000
R0[200] <= 640'h3c3fe1fffc00010000000000000000000000000000000000000001ffeefffffffffffffffffffffffffffffffffffffffffffffffe06080efce9976ffffffffffffffffffffbe000000000000000000
R0[201] <= 640'h7ffff9fffc0001000000000000000000000000000000000000000277effffffffffffffffffffffffffffffffffffffffffffffffe66000cfc0f9777fffffffffffffffffffb6800000000000000000
R0[202] <= 640'h3ffffffffff180ff00000000000000000000000000000000000000637779ffffffffffffffffffffffffffffffffffffffffffffffffe1803f049fbf7ffffffffffffffffffff6f00000000000000000
R0[203] <= 640'hffffffffffffbeff0000000000000000000000000000008000000001ffffffffffffffffffffffffffffffffffffffffffffffffffffc9993b0f1b9bfffffffffffffffffffcb6000000000000000000
R0[204] <= 640'hffffffffffffbfffc000000000000000000000000000000000000000ffeffffffffffffffffffffffffffffffffffffffffffffffffffdff7ff9f0bfffffffffffffffffffffb7000000000000000000
R0[205] <= 640'hffffffffffffffff8000000000000000000000000000000000000000cedcffff7fffffffffffffffffffffffffffffffffffffffffffffbfff333ffffffffffffffffffffffcb2400000000000000000
R0[206] <= 640'hffffffffffffffff8000000000000000000000000000003e8000000006fcffffffffffffffffffffffffffffffffffffffffffffffffffffff3f3ffffffffffffffffffffff8b6e00000000000000000
R0[207] <= 640'hffffffffffffffffc40000000000000000000000000080c78000000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff36040000000000000000
R0[208] <= 640'hffffffffffffffffc40000000000000000000000000000cf300000031feffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fffffffffffffffffffffb3e3f0100010000000000
R0[209] <= 640'hffffffffffffffffe400000000000000008000000100810f70000000097fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7ff8000000000000000
R0[210] <= 640'hfffffffffffffffffc0000000000000000000000000087fff00000000f7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3ff8000000000000000
R0[211] <= 640'hfffffffffffffffffc000000000088008100000000031ffff88080007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefe0000000000000000
R0[212] <= 640'hfffffffffffffffffe7800000000db7f0700000001823fffff008000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff8100000000000000
R0[213] <= 640'hffffffffffffffffff7800000003effe870000000100ffffff010001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1c0800000000000
R0[214] <= 640'hffffffffffffffffffff80801fffffffff000000000fffffffff0033ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff81800000000000
R0[215] <= 640'hffffffffffffffffffffc3e73ffffffffff00000013fffffffffe73fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3c0c0080000000
R0[216] <= 640'hffffffffffffffffffffffff9fffffffffec000001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbdfdb8000000000
R0[217] <= 640'hfffffffffffffffffffffffffffffffffff0000033ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1200000000
R0[218] <= 640'hfffffffffffffffffffffffffffffffffff80002ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0240000000
R0[219] <= 640'hfffffffffffffffffffffffffffffffffffc0087ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa040000000
R0[220] <= 640'hfffffffffffffffffffffffffffffffffffc40b7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa000000000
R0[221] <= 640'hfffffffffffffffffffffffffffffffffffc013efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffffffc000000000
R0[222] <= 640'hfffffffffffffffffffffffffffffffffffc4ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffffffe000060000
R0[223] <= 640'hffffffffffffffffffffffffffffffffffffccfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff100000000
R0[224] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb93dffffd000200000
R0[225] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff159ffffd002249200
R0[226] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd94dfffec000441080
R0[227] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed4ddfffec000002480
R0[228] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed8d3fffec000002c80
R0[229] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4cc2fffec082244a80
R0[230] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe5907fffe00000ea40
R0[231] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff09a7fff608040a640
R0[232] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9827ffed000010608
R0[233] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2c646ffcd000000648
R0[234] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa4405ffe4801004c04
R0[235] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff99907ffe2808208400
R0[236] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd4923ffe2008232402
R0[237] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffce465fff2000000800
R0[238] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe6c45fff108001c300
R0[239] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeff24a5dfa108006c908
R0[240] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef726e5ffb100004c920
R0[241] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfb8460dfb1a000c5804
R0[242] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfd8441df90400365204
R0[243] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfc4043bfc2420388506
R0[244] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7e22061f82788422020
R0[245] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefb730465fc1bc8063212
R0[246] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe63b904a4fd03c046210a
R0[247] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2bd80031ffa1e0071828
R0[248] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9dec1061feb160061031
R0[249] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffbc7e12047ff99a80ec810
R0[250] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7ffffde7701037ffb8f47c8842
R0[251] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbffff6f19c0877ffe04cc02081
R0[252] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffefffffb74cc106fffd8681bb0e8
R0[253] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffeffffbb6244120bbfcc327a1028
R0[254] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffdff9fffb9265010063fc602709964
R0[255] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffeddffdf6d791ace2fe1a67648c0
R0[256] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffeddffcf4b0b90c93ff9976ccc80
R0[257] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfd7a7bfff5630f919387fc472da402
R0[258] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd7fff7bffd677cf910617ff02239040
R0[259] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5f7bfffff30c7d0c387ffc01f9390
R0[260] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffb1fffff986bc9924ffe702fc320
R0[261] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff77fff1ffff5b213c9b04fff592ec658
R0[262] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb3ff63cffbed099c11127ff7833440c
R0[263] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff76ff2cffcf5c38c24c0fff0b3b63bc
R0[264] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffdb2dffffddbe61be17fd81366794
R0[265] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9e5dfbb7ffffec1b69fa9bf7801e6c11
R0[266] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf67e9b5ffffeefd83f016f9c03f21b0
R0[267] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffef2579bdfffff6d9c7b83bfce43617b8
R0[268] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffff7df8b1effff3c8c7e83bfe3abb2691
R0[269] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefff77ffc0feffff545e1f219ff33b978b8
R0[270] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbd3d9dfffdf20fe0fc0dfbf818f95c
R0[271] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfbb7bcd3ddfefb63cbb1bdbdfcda46e4
R0[272] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeefff7d8d2fffffd6263fb3dbdfe1a5670
R0[273] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffb5fc19b3fffdbe63b2ce7dfc85bf7c
R0[274] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff37ffb5ec0b267ff6af276696ffff1d9f5e
R0[275] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb3fe35cc9b7cfffef9975a6dff5f99cfb6
R0[276] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbff8de899df6ffe1d8623613bf5939fe0
R0[277] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7eddec9b36fff33e44f7c33ffcc73dda
R0[278] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3fcef6c93b7ffb9f63fb0dbbfb47bded
R0[279] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbf7fe8f28b7a7fffdfa3fbed96eb437c2c
R0[280] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffbfeee453fcfffdefc7f1f7c7dfc76793
R0[281] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fed7ef6ce9fffff6e7e7d1dfefffc77ef1
R0[282] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefed8c09ebb7fe73f3e6e7e6ffc37f1c
R0[283] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedf8fe78c3d6fdfff53f6ce65edfbe17f9e
R0[284] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7dfb3e4e97fffffc967ef6edbffe27f7d
R0[285] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffceb77f3be90dbffff7df5ef6cdbfbe2df8c
R0[286] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefe6fdfe39e8d3ff9ffecf7ffe79dfee0f9c6
R0[287] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3f9bd3ee0c6ffdffba77b3e7003f30fbfc
R0[288] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdeddf7e6cceffeffbc277fde78ffd079fe
R0[289] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3dee9facccfff7fdf26feccfed7f0ef7a
R0[290] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffb9e69d8489edf3fdf05dfb6fa6f71878c
R0[291] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcfffd9dbbec48df77ffce03ff90737ff1f76e
R0[292] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6dccf9fe648ff7fdfff83ffb3ffbfc977be
R0[293] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffae265edf741beffcfffc3ffb3ff9ff0f3fa
R0[294] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb7bdf77d9f3017ddfefff47ef7bdfdff0f772
R0[295] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcff7d1fe59fbfff7ffc6bf7fffebf8dbe0
R0[296] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbaf9bbf1be08e7fffbffc3f8fdff67f8feec
R0[297] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf7d999cfd997fecfdfdc3f2fdff7778ff7c
R0[298] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffc59b8d893dfefeeefa3d9fffefbf8ffb6
R0[299] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ff0fec3e93bffffe77e3bbfeffd8f9ff78
R0[300] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfb7c282cfc5ffffff36e0e6ff7d3cf8dfbc
R0[301] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf40ae18ddfffffb6e38f7e6c7e78e790
R0[302] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecf36e778dfffeffcce16fff29ff39ff36
R0[303] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9619967dab1fffffe2e1dfcf3bffbdf36f
R0[304] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe6f6d9f1a23ffff6ff3e3bff73f9bd87c5c
R0[305] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdab35df2b63ffee1ff9e1bff8bfffe8fc5a
R0[306] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9938adb167fffb2ffce17ffcdfffe4fc4e
R0[307] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbc16e07b843f79ffffc60ffcf8deff0fcbf
R0[308] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4af7b9e63e2bddffd21f7ff8ffff8d877
R0[309] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffffff31fadce23fcffdffd81bdffcfdffc7869
R0[310] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffffffffffd9dfd4e643fbffdd3d81ffffb7f9fc3031
R0[311] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8fdfce466367ffbfb6e1ffff723ffcb831
R0[312] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffffffffffff7ffef6fef52e66ff7ffe4c1bfff5b37fcca74
R0[313] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda5f330e37fffffb2c0fffcdbcffce0de
R0[314] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffbfff7d3fbb9e3ef7f9f38e1fff9edbffc80ce
R0[315] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffbfffffffffff7e3fc8df1edffbefceb7ff3ec3bfcd246
R0[316] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffbffffffdfffff79fe4ce1cbf7bfff697ff7aefdfee260
R0[317] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffeffff39f7646243dabdfd09ffefef7fdee040
R0[318] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffded8f7b460836bbbfee9efdfef3fdec651
R0[319] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedfff7fffffffffffff633da48dbe89bfee17fb6773fee4602
R0[320] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5fff77fffffef3fffb619c20adb3cb7ffc17f2fa59ff89bb2
R0[321] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6ffffffffffefdfff9eccf021d9fe0fe7817a7ef7dffc3199
R0[322] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefeffffffdbeaf7ef91f861018e33dfe138fffddfec7249
R0[323] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffefffffffeb235c75987c680c17373fc933ffe5ef3c3ee0
R0[324] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee7ffffff63f69f39be3e6c1f7f237ec967ffe3e7fc4830
R0[325] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffffeeeefdfffff7bfbfffc7f9824ce3e3774c14ff7eda7fc7877
R0[326] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffefffe7ffffffffffbfdfffe3fc874c43f16f1c11dfedfc7fe36e7
R0[327] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffdffff7dfffffffff3ecd1ed8de6344e1f4dfbc91effd572fe6eef
R0[328] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfff7fdf7ffffdf7ed7ffd8d2b12275f62fb89367fbb5bfc588e
R0[329] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffbdffff7f7efffffcefff9ff1b19c1e376766f3c02f7f9bf9f838d6
R0[330] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffeffef7ffffffffeebfbcff81b9e081a0f37edc87bfd0be0fc66db
R0[331] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fff7fdffffffe4fbb67c907df0083270fedc87d3873f0ec76bb
R0[332] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffb7fffdfffff7f7ff1e2c667b2d9e2669fc83c3ff3fcf8676f
R0[333] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffdbbfffbffff73fffcf8ce13924c3277bfc1b1f6fffe76744f
R0[334] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffff3fdffdffff7ffffb3d0fc3000c2cb77c81d77efffb6e6e3f
R0[335] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefefdfbfff3f3fffffff7fefbf9dcff30c6628d3ff884ffefffb1c7cff
R0[336] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7efdbefff3b7ffdffffedffdee0e7fc8c600a65b9c867fefbfb3e787e
R0[337] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffdfe7ffbf7fedfff7edfffe6867fe0e60c22df98c37befffed63efe
R0[338] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffdfdf7bfbf7ffdffb77bffbe6d03fb8f30630dff0837fff7fdc61aff
R0[339] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb7ffba7ffdf7df7fffcf7dc3afc3338821db487bfff3f9ca327f
R0[340] <= 640'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfdff5bff9b7ffdefdb7bbffeddb1bfc11b0c62ca4839eff3f7ee333d
R0[341] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffbff9dfb9e7bffffef737ff76db039a21b63558ccc3dbfffeee62a7f
R0[342] <= 640'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf3ff9dff9e77fffff37bffb360723fc3191211ccc63efff3def21c1f
R0[343] <= 640'hefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffff2cffdeefddfffa4fef37807b9dc388d201f4863e3bf1bff23b6f
R0[344] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeefbef3dffdeffffbfff7f1fb7df3bc35084c00936c63f3ffe3ff83b7b
R0[345] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3fb7fffccfffffffd3bffedde99f9f998211006d61fb776ffd83f39
R0[346] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3fdbb7fcdffedfffe7befdcbe45fc7088201858861789f59fcc0f77
R0[347] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff93b7fbbffcdfbfdbffeddffdff480ae10c47430f00319886078243d67
R0[348] <= 640'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf33ff7dffd37ff5f7fe7eff1ffef2c120cc0c10723118820431363f27
R0[349] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddffffffffffffffffffffffffffe33df7e4f73f7f7f3fefdbf7ffe6bf4b04c480d181108b0606ff21f2b
R0[350] <= 640'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffffffffffffffffde33ff2f6ffbeffbfbfefdff7fff5d7e1803080d982000000277b41b2d
R0[351] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffffffeb3fcbfb7fbfffcfdf6f9fdf7ff7e3fc4030040e074010004ef661b3b
R0[352] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffffffffffffffffffffffffffffffffffefbf4ffbbfbbffdfffcfbfdf7ed67bfe08609217032c10025bd761dbf
R0[353] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffffffffffffffffffffffffffff3fd7fdbdbfff8fefdfdfffdef3f9bf8000135f676c1c0267f2c193e
R0[354] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7b7fffebdafff8fffceff7fef93fcefc060084fe76c280067f980d1b
R0[355] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffff73bbdfe7f9fffdff7cfbfdfeeb6de7fc0300026c120098047eb001af
R0[356] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedeffffffffffffffffffffffffffffffffffde7fedfd7fbfff5ff9d79fbff7f3f39f80002081c03012004f7b00824
R0[357] <= 640'hdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffffffffffffffffffffffffff7ef657effff1fffcffcf7bb7f89f3fb9ea0003481c630100007fd0030c
R0[358] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9f7fffffbf6ffffffffffffffffffffffffffff7e76efbf1befcfffdfb6fff8737ccca00002444130020006ec00980
R0[359] <= 640'hdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffffffbfeffffffffffffffffffffffffff7efe78ff9b3fffcfff1fbdfffe317dc42000030189000000003c01800
R0[360] <= 640'hffff7bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffbfffffffffffffffffffffffffffffe5efedfdf3ff7ddff87bbffff097f80800003000d800000000401800
R0[361] <= 640'hf3dbd6fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd7fbffffdfffffffffffffffffffffffffffefe59ff3fdf3dffcbff8fb7efff01fa40000000008cc00000001402c00
R0[362] <= 640'hde00fbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffff9ffffffffffffffffffffffffffff7ffbef7fef3dffdbffdf8fe7ffb10000000300808ec00040003420000
R0[363] <= 640'hec003f77ffffffffffffffffffffff03ffffffffffffffffffffffffffffffffff9fffffeffefffff7fffffffffffffffffdffbffb9e7fef3dfffeff971e77ff380000800100408e400000000240000
R0[364] <= 640'h98001fbffffffffffffffffffffffe03fffffffffffffffffffffffffffffffffddf5fffeffbffffffffffffffffffffffffffd77ffdfff73ffffbff9fbfff7e1c0000080000600f000000000600000
R0[365] <= 640'he000006ffcfffffffffffffffffffe03fffffffffffffffffffffffffffffffcfde7ffffe9fffffffffffffffffffffffffffff7ffe77ff3efffcbff9b3fedfe1c00004c01002007000000000000000
R0[366] <= 640'hc000003fefbfffffffffffffffffff02fffffffffffffffffffffffffffffffaf4fffffff1fbfffffffffffffffffffffffffff3eff77ff9feffcfff9e7ff9fe1800000201028007020000000000000
R0[367] <= 640'h87f9ffffffffffffffffffe03fffffffffffffffffffffffffffffffdfceffffffcfffffffffffffffffffffffffffff2df5f3ffc9fffcfff9d7cfdff1c0080020402c007000000000040800
R0[368] <= 640'h18ff3fffffffffffffffff02fffffffffffffffffffffffffffffffdffdffffffdffffff7ffffffffffffffffffffff3df3dbbfe5bffdfff9dffbdfe0c00d80c0000c004000000000001800
R0[369] <= 640'h39e37f9bffbffffffffb027ffffffffffffffffffffffffffffffbfedffffffdfcffff7fffffffffffffffffffdfff3f7dbfdf1f7fefff9e7ffdff0400e28e00002000000000000920000
R0[370] <= 640'h7fd5e7ffefffffffff03ffffffffffffffffffffffffffffffdcfdb7fffffdfcffff7bffffffffffffffffffefed3fffbdff1f7fefff9e77f6fd0001ce4700000000800000000000000
R0[371] <= 640'h23f8deffffffffffff00cfffffffffffffffffffffffffffffccfd9ffffffffcfffffbffffffffffffffffffffee3ffbdffb1fffcfff9e7ffffc2001fe8000000002a00000000040000
R0[372] <= 640'hcff3dfbffffffffe0071e3ffffffffffffffffffdfffffffe7fe9ffeffedfeffffffffffffffbffffffffffffc7cff4fff1efbefff9e5ffffe0000be1000000002200000000020000
R0[373] <= 640'h31feffffffffff0001fffffffffffffffffffcfffffffffc7ee9fff7ffdbdfffffffffffffffffffffffffbfd7cf69fff1effeffb9edff3fe0004780000000000404000000000000
R0[374] <= 640'h3effffffff00000fffff23ffffffffffffcffffffd8dd13bd7ff7fffbdffff7fffffffffdfffffffffdffc7bf75fffbe7feffdbf3fe1bf0000201800000000002000000200000
R0[375] <= 640'h17ffffffff00000fffffffffffffffffffdf3fffff05c032dbbedfffbcfbff7fffffffffffffffffffeff477fadfbfbe7fefffbe7fe17f0000323e00000100000000000000000
R0[376] <= 640'h7cfffff00000fffffffffffffffffffd77fffff058032db7cfe7c3cfbffffffffffffffffffffffe7f627fbcfff9effefffbeffc07c000f98db00000500000000000000000
R0[377] <= 640'h3ff7ff00001ffffffffffffffffff7dfdfffef4f403019f9fcfc7ef3ff7ffffffffff7ffffffffe7761effefff9f7fcfff1e6320df000fccdc00000000000000000000000
R0[378] <= 640'h63ff8c0001fffffffffffffffffffd89affd97f40000bff7ffe7cfbff3dffffffffffffffffffe27b1cffeff79fffcfff035ff0ff0008000c00000000000000000000000
R0[379] <= 640'h3ff80001ffffffffffffffffffcd99de7e86f01244ffffffe7af3ff9dfffffffffffffffffb803800117fff9effcc8196fff1fe0000c00400000000000000000000000
R0[380] <= 640'h1f7c0001ffffffffffffffffffcce07e740cd00b70f3dfffe7ce7ff7dffffffeffffffffffb000000003ffe1e47c1cfbf7ff0fe0003e08000000000000000000000000
R0[381] <= 640'h180001ffffffffffffffffffa4e1bf3019dcf020e7dfffc7fe7ffbffffffff7fffffffff800000000015c036fcfefbeffd07e2001e00000000000000000000000000
R0[382] <= 640'h1ffffffffffffffffff4c71f81016fc7831cfdfffe3dffffbffffffffdffffffffc000000000000f133fefffbe71f87e0000000000000000000000000000000
R0[383] <= 640'h1ffffffffffffffffffc6e0f800389e3896df9fffffeffffbbfffffffffffffffe000000000000001fbfefff3ef1f81e0000000000000000000000000000000
R0[384] <= 640'hf87ffffffffffffffff8c0f0600cdbdfc63ebfffffeffff9dfffffffffbfffff0000000000000000f9fcffb3ef9c06e0000000000000000000000000000000
R0[385] <= 640'hffffffffffffffffc48e4f1064d5f873f7fffe1ef7ff8dfffffffffbffffc00000000000000003cfefff3ee1f0760000000000000000000000000000000
R0[386] <= 640'h3fffffffffffffffc08f6d40258db83377ffff0fe7ff0dfffffffffbf3ba0000000000000000000000463ef7f87e0000000000000000000000000000000
R0[387] <= 640'h1fffffffffffffff708f010807197263f7ffbf43187e8ffffffffffbf8f80000000000000000000000001680c0300000000000000000000000000000000
R0[388] <= 640'h7fffffffffffc00780f8140779c3f33fffb6f60587f2cff97fffffffff0000000000000000000000000000000200000000000000000000000000000000
R0[389] <= 640'h1fffffffffff80000010201bbfb3f37f7fff660400804ebfffffffdffc0000000000000000000000000000000000000000000000000000000000000000
R0[390] <= 640'h7ffffffffe000000000002dbff7da7e7fb0800000f44fffffffffff000000000000000000000000000000000000000000000000000000000000000000
R0[391] <= 640'h1ffffff000000000000000e3fdff27f7f10000000780fffff3fff00000000000000000000000000000000000000000000000000000000000000000000
R0[392] <= 640'h7fffff00000000000000001641601cefe0000000000ef800000000000000000000000000000000000000000000000000000000000000000000000000
R0[393] <= 640'h17ffff00000000000000000093e07cff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[394] <= 640'h1ffe00000000000000000017fb7c9c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[395] <= 640'he310000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[396] <= 640'h0
R0[397] <= 640'h0
R0[398] <= 640'h0
R0[399] <= 640'h0
R0[400] <= 640'h0
R0[401] <= 640'h0
R0[402] <= 640'h0
R0[403] <= 640'h0
R0[404] <= 640'h0
R0[405] <= 640'h0
R0[406] <= 640'h0
R0[407] <= 640'h0
R0[408] <= 640'h0
R0[409] <= 640'h0
R0[410] <= 640'h0
R0[411] <= 640'h0
R0[412] <= 640'h0
R0[413] <= 640'h800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[414] <= 640'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[415] <= 640'h60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[416] <= 640'h18000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[417] <= 640'h7000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[418] <= 640'h800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[419] <= 640'h300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[420] <= 640'hc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[421] <= 640'h14000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[422] <= 640'h3000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[423] <= 640'hc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[424] <= 640'h780000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[425] <= 640'h60000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[426] <= 640'h1c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[427] <= 640'h0
R0[428] <= 640'h1f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[429] <= 640'hff000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R0[430] <= 640'h0
R0[431] <= 640'h0
R0[432] <= 640'h0
R0[433] <= 640'h0
R0[434] <= 640'h0
R0[435] <= 640'h0
R0[436] <= 640'h0
R0[437] <= 640'h0
R0[438] <= 640'h0
R0[439] <= 640'h0
R0[440] <= 640'h0
R0[441] <= 640'h0
R0[442] <= 640'h0
R0[443] <= 640'h0
R0[444] <= 640'h0
R0[445] <= 640'h0
R0[446] <= 640'h0
R0[447] <= 640'h0
R0[448] <= 640'h0
R0[449] <= 640'h0
R0[450] <= 640'h0
R0[451] <= 640'h0
R0[452] <= 640'h0
R0[453] <= 640'h0
R0[454] <= 640'h0
R0[455] <= 640'h0
R0[456] <= 640'h0
R0[457] <= 640'h0
R0[458] <= 640'h0
R0[459] <= 640'h6000000000000000000000000000000000000000000000000000000
R0[460] <= 640'h0
R0[461] <= 640'h0
R0[462] <= 640'h0
R0[463] <= 640'h0
R0[464] <= 640'h0
R0[465] <= 640'h10000000000000000000000000000000000000000000000000
R0[466] <= 640'h12038000000000000000000000000000000000000000000
R0[467] <= 640'h0
R0[468] <= 640'h0
R0[469] <= 640'h489000000000000000000000000000000000000000000000
R0[470] <= 640'h0
R0[471] <= 640'h0
R0[472] <= 640'h0
R0[473] <= 640'h0
R0[474] <= 640'h0
R0[475] <= 640'h0
R0[476] <= 640'h0
R0[477] <= 640'h0
R0[478] <= 640'h0
R0[479] <= 640'h0
end
always @(posedge vga_clk) begin
R1[0] <= 640'h0
R1[1] <= 640'h0
R1[2] <= 640'h0
R1[3] <= 640'h0
R1[4] <= 640'h0
R1[5] <= 640'h0
R1[6] <= 640'h0
R1[7] <= 640'h800000000000000000000000000000000000000000000000000000000000000000
R1[8] <= 640'h80000000000008000000000000000000000000000000000080000000000000000000
R1[9] <= 640'h4000000000000000000000000000000000000000000000000000000000000000
R1[10] <= 640'h4000000000000000000000000000000000000000000000000000000000000000
R1[11] <= 640'h30100000000000000000000000000000000000000000000000100000000000000
R1[12] <= 640'h20000001070104000000000000000000000000000000000000000000000000000000000000
R1[13] <= 640'h103400c000000000000000000000000000000000000000000000000000000000000
R1[14] <= 640'he008000000000100000000000000000000000000000000000000000000000000
R1[15] <= 640'h180800100803800690000000000c000000000000000000000000000000000000000000000000000
R1[16] <= 640'h6006000400381e0e130010680c48000000040000000000000000000000001000081000000000000
R1[17] <= 640'h6000000181e0c000000480048400000002000000000000000000000001000000000000000000
R1[18] <= 640'h20000601ff3ec0c360e603068c07008002000000000000000000000000000000000000000000
R1[19] <= 640'h3fc1ff3f1ec7206f00030407000000000000000000000000000000010000000000000000
R1[20] <= 640'h90000003cc0ff3ffffe016ff0630e030000c0000000000000000000000084000000000000000000
R1[21] <= 640'h800000010000009800ff7fff7c03eef8e6ff03000080000100000000000000000080000000000000000000
R1[22] <= 640'h6008880999effffff79fffefcceffff663001000100000000000000000000330000000000000000
R1[23] <= 640'h18000000000000000000000000000000000000002010099102138660098879fffffffce79ffff7f0e78ff66708900e000000000000000000020008001000000000000
R1[24] <= 640'h40010001cc38638373ffffffffeffffffffff66ffff01f0c43038000000000000000300c0180006000000000000
R1[25] <= 640'h4011803839992387fc7fffffffffffeffffff66ffff83e16671f080000000000000000000800000000000000000
R1[26] <= 640'h18000000000000000000000000000000000000000004079ec7c318f67bfef7ffffffffffffffffff7fffffffff73e3e78200c000000000000021c00080000000000000
R1[27] <= 640'he038000000000000000000000000000000000000000000ffcec7c7c3bff3ff7ffffffffffffffffffffffffffffff2f3e7fe008000000000002131800000000000000000
R1[28] <= 640'h3e0000000000000000000000000000000000000000001ffcf3fffe7fff3ff7fffffffffffffffffffffffffffffe638ff3c000c0000000000218e108001000000000000
R1[29] <= 640'h100fe3000000000000000000000000000000000000000001ffcf3fff7effffffffffffffffffffffffffffffffffff0e38fc3c040e0000000003008c38c000000000000000
R1[30] <= 640'h1b2fcffe00000000000000000000000000000000000000019ffffffff7efffffff7ffffffffffffffffffffffffffff2f7bfe388e380000000001808c00c020000000000000
R1[31] <= 640'h1b71efe0300000000000080000000000000000000000000b9ffffffffffbfffff7fffffffffffffffffffffffffffe777f7ff61ce7800000000c0cef8c00862200000000000
R1[32] <= 640'h171dbdfbffcfddc00001201000118000000000000000000000e7f7ffeffffffffffffffffffffffffffffffffffffff7efff89d7fff07c000000113694603400c38080000000000
R1[33] <= 640'h1013b7ffffffff3fb000010010000000000000000000000000cff7fffffffffffffffffffffffffffffffffffffffffffffffff9f7f7ef00300ff001169c603e00001000000000000
R1[34] <= 640'h1003f7ffffffff3f3000010000300200000000000000000000e7fffffffffffffffffbfffffffffffffffffffffffffffffffffdfff7ef81f71f03cf96dc77ffee383000000000000
R1[35] <= 640'hcfffeffffff7ffb80000300030060000000000000000006837ffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ff3f7b003ef96dfefffe71c0880000000000
R1[36] <= 640'h800cfffefffffffffcc03f030018180400000000000000010fc3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffe73ffcffffff9fef3efffe78f8000000000000
R1[37] <= 640'h8efffffffffffffccc3fb2c018088c000000000000000107fcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcde1fe79fefbcffbd7c3f010000000000
R1[38] <= 640'heffffffffffffffffcc83b0c0181f99000000000000000173feffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00ffdffffffffffcffb10010000000
R1[39] <= 640'h8000018cf3fffffffffffeffdc01b2c0c73f99300000000000016073fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffdffffffeff810030000000
R1[40] <= 640'h40003001800fffffffffffffffffeffffff3ff3ff00010000000000c71fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fffffffff7fffffffffff8ec3e301040000
R1[41] <= 640'hc66ffffffffffffffffffffffff7f3fffe0300000000000cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcfe0c100000000
R1[42] <= 640'h7fefffffffffffffffffffffffffefeffe03000000000107fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7cf840808000
R1[43] <= 640'he0c7fffffffffffffffffffffffffffffcfff00000000001007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7cffe0800000
R1[44] <= 640'hf03c3ffffffffffffffffffffffffffffffff88000000003007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000
R1[45] <= 640'h73cfffffffffffffffffffeffffffffdfffff8000000001007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3efe000000
R1[46] <= 640'h3077ffffffffffffffffffffffffffffffffff80c0000000008ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1fde180000
R1[47] <= 640'h7e17ffffffffffffffffffffffffffffffffff81c00000000f8fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffff8e3c0000
R1[48] <= 640'h300bfff3fffffffffffffffffffffffffffffbfff03f0000001883fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffffffffefffffffe010000
R1[49] <= 640'h331f7ffbfffffffffffffffffffffffffffffffff0e0008002000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000
R1[50] <= 640'h3dc9ffeffffffffffffffffffffffffffffffffe0c0008000003efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcff780000
R1[51] <= 640'h103dedffffffffffffffffffffffffffffffffffef001000000813ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefff00000
R1[52] <= 640'h1801009effeffffffffffffffffffffffffffffffffeff00000000c3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffffffffffffffffffffffc00000
R1[53] <= 640'h1800000fffe7fffffffffffffffffffffffffffffffffff8000018c3e7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffffc00000
R1[54] <= 640'he1ffff7fffffffffffffffffffffffffffffffffff0000099fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcc00000
R1[55] <= 640'h81000e317f7fffffffffffffffffffffffffffffffffffe3800018ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3cf00000
R1[56] <= 640'h36283fcfffbffffffffffffffffffffffffffffffff6f88e00303fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3800000
R1[57] <= 640'h20030ffffffffffffffffffffffffffffffffffffffec0000303ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800000
R1[58] <= 640'h11800010ffffffffffffffffffffffffffffffffffffffec000001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000
R1[59] <= 640'h309900fc7fffffffffffffffffffffffffffffffffffff1c00001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000
R1[60] <= 640'he39900fcff7fffffffffffffffffffffffffffffffffff1c00011ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000
R1[61] <= 640'hc380000fef7fffffffffffffffffffffffffffffffffff8040c11ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000
R1[62] <= 640'h3c704100fffffffffffffffffffffffffffffffffffffff8300c11ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000
R1[63] <= 640'h83014610fcffffffffffffffffffffffffffffffffffffff0c00781ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe300000
R1[64] <= 640'h37cf873fffffffffffffffffffffffffffffffffffffec00000007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ecc0000
R1[65] <= 640'h1fefc73fffffffffffffffffffffffffffffffffffffe8400000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0c000
R1[66] <= 640'h3000ff3fffffffffffffffffffffffffffffffffffffffff8f0000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff70fc00
R1[67] <= 640'hcff1ffffffffffffffffffffffffffffffffffffffffd8e0000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0fc00
R1[68] <= 640'hc1187f1ffffffffffffffffffffffffffffffffffffffffdfc00103fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffccf080
R1[69] <= 640'he1307f3fffff7ffffffffffffffffffffffffffffffffffffc00103fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffce4080
R1[70] <= 640'h70717cfcffffffffffffffffffffffffffffffffffffffffffe089ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcc6000
R1[71] <= 640'h3873fcf8fffffffffffffffffffffffffffffffffffffffffff081ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff71f830
R1[72] <= 640'h6fe7f89fffffffffffffffffffffffffffffffffffffffffffc066ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7cf7c0
R1[73] <= 640'h6667fc8bffffffffffffffffffffffffffffffffffffffffffc066fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcffc0
R1[74] <= 640'hf4679c81ffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffccfcc0
R1[75] <= 640'hf00e9c81ffffffffffffffffffffffffffffffffffffffffffff3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcc7cc0
R1[76] <= 640'hf818d99dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcffcc0
R1[77] <= 640'hd919db9fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7ff00
R1[78] <= 640'hff9fff9fffffffffffffffffffffffffffffffffffffffffffff9fffffffffffffffffffffffe11fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff71ff00
R1[79] <= 640'hffdbff9fffffffffffffffffffffffffffffffffffffffffffff9fffffffffffffffffffffffe038fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9ff00
R1[80] <= 640'hfefff0f7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00
R1[81] <= 640'h3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00
R1[82] <= 640'hffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcf00
R1[83] <= 640'hfe7fff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc40
R1[84] <= 640'hffffffffffffffffffffffffdffffffffffeffffffffffffffffffffffffffffffffffffffff00003ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc40
R1[85] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc40
R1[86] <= 640'hffffffffffffffffffffffffffffffffffefffffffffffffffffffffffffffffffffffffffff000001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefc0
R1[87] <= 640'hff7fffffffffffffffffffff63fffffffffffffffffffffffffffffffffffffffffffffffffe000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7c1
R1[88] <= 640'hdeffffffffffffffffffff630fffffffffffffffffffffffffffffffffffffffffffffffffff000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8fc0
R1[89] <= 640'hffffffffffffffffffffffffe7fffffffff7ffffffffffffffffffffffffffffffffffffffff000018fffffffffffffffffffffffffffffffffffeffffffffffffffffffffffffffffffffffffffffc0
R1[90] <= 640'hfffffffffffffffffffffeffc067ffffffcffffffffffffffffffffffffffffffffffffffffe00001c7ffffffffffffffffffffffffffffffffffefffffffffffffffffffffffffffffffffffffffbe0
R1[91] <= 640'hfffffffffffffffffffffe000367ffffffcffffffffffffffffffffffffffffffffffffffffe00000f7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9e0
R1[92] <= 640'hfffffffffffffffffffffe000167ffffffffffffffffffffffffffffffffffffffffff0ffffe000007ffffffffffffff3fffffffffffffffffffff1efffffffffffffffffffffffffffffffffffff9e1
R1[93] <= 640'hfffffffffffffffffffefc000080fffffcfefffffffffffffffffffffffffffffffffffffffe0000049fffffffffffff8fffffffffffffffffffff983ffffffffffffffffffffffffffffffffffff9e1
R1[94] <= 640'hfffffffffffffffffffffc000090fffff9007ffffffffffffffffffffffffffffffffffffffe0000003fffffffffffff87ffffffffffffffffffff080fffffffffffffffffffffffffffffffffffffc1
R1[95] <= 640'hffffffffffffffffffffc0000098ffff91017e7ffffffffffffffffffffff7fffffc7fffbeff0000003fffffffffffe31fffffffffffffffffffff0c07fffffffffffffffffffffffffffffffffffe61
R1[96] <= 640'hffcfffffffffffffffff8000000cffc038c11ffffffffffffffffffffffffffffff3cff9ffff60000dfffffefff3e0008ffffffffffffffffffffe420fffffffffffffffffffffffffffffffffffe7f8
R1[97] <= 640'hffffffffffffffffffff000000009e00000008feffffffffffffffffffffffff8f70873fffff6000093ffffffc7100008fffffffffffffffffffffe09ffffffffffffffffffffffffffffffffffff6ff
R1[98] <= 640'hffffffffffffffffffff000000000000000000787fffffffffffffffffffffff9f00031fffff00000001ffc7fc2000000ffffffffffffffffffffff8effffffffffffffffffffffffffffffffffffcc7
R1[99] <= 640'hffffffffffffffffffff0000000000000001003b7fffffffffffffffffffffff1c0001dfffff000000036ffc6600000003fffffffffffffffffffff8e7ffffffffffffffffffffffffffffffffff7eef
R1[100] <= 640'hfffffffffffffffffffe00000000000000000003ffffffffffffffffffffeffe980000ffffff000000016ff02700000000fffffffffffffffffffff966fffffffffffffffffffffffffffffffffffffe
R1[101] <= 640'hfffffffffffffffffffe00000000000000000003fffffffffffffffffffffffcc000000fffe00100000065c100000000037ffffffffffffffffffef9effffffffffffffffffffffffffffffffffffbfc
R1[102] <= 640'hfffffffffffffffffffe000000000000000000008ffffffffffffffffffffefc8000002fffc00000000060810000000002fffffffffffffffffffffc8ffffffffffffffffffffffffffffffffffff9ff
R1[103] <= 640'hfffffffffffffffffffe000000000000000000001cffffffffffffffffffeffe180000663fc00000000060000000000000fffffffffffffffffffffc811fffffffffffffffffffffffffffffffffffff
R1[104] <= 640'hfffffffffffffffffff60000000000000000001000fffffffffffffffffffffc4000001f49200000000000000000000000ffffffffffffffffffff8101fffffbffffbffbfffffffffffffffffffffff0
R1[105] <= 640'hfffffffffffffffffff60000000000000000000000ffffffffffffffffffff4800000007e90000000000000000000000001fffffffffffffffffff98000ffffffc7ffffffffffffffffffffffffffff0
R1[106] <= 640'hfffffffffffffffffff000000000000000000000017fffffffffffffffff7fc80400000f680000000000000000000000001ffffffffffffffffffff800007f9e8c1fffffffffffffffffffffffffffce
R1[107] <= 640'hffffffffffffffffffb90000000000000000000003ffffffffffffffffffffcc00000007090000000000000000000000001fffffffffffffffffffe000c0331e000fffffffffffffffffffffffffffce
R1[108] <= 640'hffffffffffffffffff9a000000000000000000000087ffffffffffffffffde4800000007000000c00000000000000000001fffffffffffffffffffe00001013000009fffffffffffffffffffffffffce
R1[109] <= 640'hffffffffffffffffffba80000000000000000000001c7fffffffffffffffce6c00000000000000000000000000000000000fffffffffffffffffffe00000012000001fffffffffffffffffffffffffcf
R1[110] <= 640'hfffffffffffffffffff6800000000000000000000008e7ffffffffffffff8ecc000000000000000000000000000000000007ffffffffffffffffffe00000000000007fffffffffffffffffffffffffff
R1[111] <= 640'hfffffffffffffffffff6000000000000000000000003c0ffffffffffffffc7c0000000000000000000000000000000000007ffffffffffffffffffe0000100080000ffffffffffffffffffffffffffff
R1[112] <= 640'hfffffffffffffffffffc800000000000000000000002019fffffffffffffdf7c000000000000000000000000000000000003ffffffffffffffffffc00000000080003ffffffffffffffffffffffffffc
R1[113] <= 640'hfffffffffffffffffffc800000000000000000000000011fffffffffffffff60000000000000000000000000000000000003ffffffffffffffffffd1000000000000fffffffffffffffffffffffffffc
R1[114] <= 640'hffffffffffffffffffff000000000000000000000000003fffffffffffffe740000000000000000000000000000000000007ffffffffffffffffff80000000000000cffffffffffffffffffffffffffe
R1[115] <= 640'hfffffffffffffffdffff00000000000000000000000000fffffffffffffffec0000000000000000000000000000000000007ffffffffffffffffff800000000000001fffffffffffffffffffffffffff
R1[116] <= 640'hfffffffffffffffffff800000000000000000000000001fffffffffffffffc48000000000000000000000000000000000003fffffffffffffffffff40000016000003ffffffffffffffffffffffffff3
R1[117] <= 640'hfffffffffffffffffffc00000000000000000000000001ffffffffffffff3c08000000000000000000000000000000000000ffffffffffffffffffe00000006000007ffffffffffffffffffffffffffb
R1[118] <= 640'hffffffffffffffffffff00000000000000000000000000fffffffffffffffc00000000000000000000000000000000000000ff1fffffffffffffffe60000180000003fffffffffffffffffffffffffff
R1[119] <= 640'hffffffffffffffffffe1c0000000000000000000000000ffffffffffffffe000000000000000000000000000000000000000001ffffffffffffffffffc12010000007fffffffffffffffffffffffffde
R1[120] <= 640'hfffffffffffffffffffc80000000000000000000000000ffffffffffffffc700000000000000000000000000000000000002227fffffffffffffffffffcfc63800013ffffffffffffffffffffffffcff
R1[121] <= 640'hffffffffffffffffffe3000000000000000000000000001fffffffffffffe00000000000000000000000000000000000000200ffffffffffffffffffffffefe00001ffffffffffffffffffffffffffff
R1[122] <= 640'hfffffffffffffffffff300000000000000000000000003ffffffffffffffe00000000000000000000000000000000000000000fffffffffffffffffffffffff0003fffffffffffffffffffffffffffff
R1[123] <= 640'hffffffffffffffffffff00000000000000000000000007ffffffffffffff7000000000000000000000000000000000000000023fbffffffffffffffffffffff8c17fffffffffffffffffffffffffffff
R1[124] <= 640'hfffffffffffffffffffe0000000000000000000014c31fffffffffffffff7000000000000000000000000000000000000000003f9ffffffffffffffffffffffe00fffffffffffffffffffffffffffffb
R1[125] <= 640'hffffffffffffffffffff0800000000000000000000037ffffffffffffffff000000000000000000000000000000000000000003817ffffffffffffffffffffffffffffffffffffffffffffffffffffff
R1[126] <= 640'hfffffffffffffffffff71800000000000000000000007ffffffffffffffff800000000000000000000000000000000000000000003ffffffffffffffffffffffffffffffffffffffffffffffffffffff
R1[127] <= 640'hfffffffffffffffffffb00000000000000000080000083ffffffffffffffec00000000000000000000000000000000000000000002ffffffffffffffffffffffffffffffffffffffffffffffffffbffe
R1[128] <= 640'hffffffffffffffffffcec02000000000000000000000013fffffffffffffc0000000000000000000000000000000000000000000007fffffffffffffffffffffffffffffffffffffffffffffffffffff
R1[129] <= 640'hfffffffffffffdfffef01800000000000000000000000047ffffffffffffc0000000000000000000000000000000000000000000007fffffffffffffffffffffffffffffffffffffffffffffffffffff
R1[130] <= 640'hfffffffffffffdfbfcf01880000000000000000000000007ffffffffffffd0000000000000000000000000000000000000000000003bffffffffffffffffffffffffffffffffffffffffffffffffffff
R1[131] <= 640'hfffffffffffffffbffc0018000000000000000000000003fffffffffffffc0000000000000000000000000000000000000000000001bffffffffffffffffffffffffffffffffffffffffffffffffffff
R1[132] <= 640'hfffffffffffffffc8180018000000040000000000000007fffffffffffffc00000000000000000000000000000000000000000000000e2ffffffffffffffffffffffffffffffffffffffffffffffffff
R1[133] <= 640'hfffffffffffffffc0080000004000000000000000000c1fffffffffffffbc00000000000000000000000000000000000000000000000003fffffffffffffffffffffffffffffffffffffffffffffffff
R1[134] <= 640'hfffffffffffffffe00000c0000000000000000000000fb1ffffffffffffb000000000000000000000000000000000000000000000000001bffffffffffffffffffffffffffffffffffffffffffffffff
R1[135] <= 640'hfffffffffffffff600008e00000000000080000000030039ffffffffffff00000000000000000000000000000000000000000000000000017fffffffffffffffffffffffffffffffffffffffffffffff
R1[136] <= 640'hffffffffffffff701000010000000000000000000000011fffffee3fff9c00000000000000000000000000000000000000000000000000001fffffffffffffffffffffffffffffffffffffffffffffff
R1[137] <= 640'hfffffff33f7ffff080000000000000000000000000000003ffffee9fff9800000000000000000000000000000000000000000000000000001fffffffffffffffffffffffffffffffffffffffffffffff
R1[138] <= 640'hffffdff21fffffd8800000010000000000000000000000027fff020ff89080000000000000000000000000000000000000000000000000001cffffffffffffffffffffffffffffffffffffffffffffff
R1[139] <= 640'hfffeffbe3fffff988000000000000000000000000000000073ff0118780000000000000000000000000000000000000000000000000000001c3fffffffffffffffffffffffffffffffffffffffffffff
R1[140] <= 640'hffffffb0073fff184000800000000000000000000000000001ff113878040000000000000000000000000000000000000000000000000000800fffffffffffffffffffffffffffffffffffffffffffff
R1[141] <= 640'hffff7b80033ffcc3c000000000000000000000000000000001ff01d163800000000000000000000000000000000000000000000000000000003fefffffffffffffffffffffffffffffffffffffffffff
R1[142] <= 640'hffff668001fffce6c60000000000000000000000000000000070608c0300000000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffff
R1[143] <= 640'hfffde61000fffeeeee60300000000000000000000000000000f8601c3c0000000000000000000000000000000000000000000000000000040d1f7fffffffffffffffffffffffffffffffffffffffffff
R1[144] <= 640'hfffff6c0017fff3e7ed84000000000000000000000000000007fe88c388100000000000000000000000000000000000000000000000000036167ffffffffffffffffffffffffffffffffffffffffffff
R1[145] <= 640'hffffffdc016fff7ff7f9020000000000000000000000000000ffc9c0e3000000000000000000000000000000000000000000000000000103767fffffffffffffffffffffffffffffffffffffffffffff
R1[146] <= 640'hfffffffc81fffffffffd0700000000000000000000000000037f4980438000000000000000000000000000000000000000000000000003fffeffffffffffffffffffffffffffffffffffffffffffffff
R1[147] <= 640'hffffffff99fffffffffd0c10000000000000000000000000017f400100c800000000000000000040000000000000000000000000000001fffeffffffffffffffffffffffffffffffffffffffffffffff
R1[148] <= 640'hffffffffdfffffffffffcef800000000000000000000000000ffe83000c000000000000000000000000000000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffff
R1[149] <= 640'hffffffffffffffffffff9effe00000000000000000000000007f49f001c20000000000000000000c3e01000000000000000000000000007fffffffffffffffffffffffffffffffffffffffffffffffff
R1[150] <= 640'hffffffffffffffffffffbfffe00000000000000000000000037fe8c003e4000000000000000000003ffb60000000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffff
R1[151] <= 640'hfffffffffffffffffffffffff00000000000000000000000007fe80018e000000000000000000007fff9e0000000010000000000000000f1fffffffffffffffffffffffffffffffeffff67ffffffffff
R1[152] <= 640'hfffffffffffffffffffffffff80010000000000000000000003fb93806c0800000000000000000007fff7c66000000000000000000000c3effffffffffffffffffffffffffffff99c78f3fffffffffff
R1[153] <= 640'hfffffffffffffffffffffffffc8000000000000000000000001f993843f8000000000000000000007ffff700000000000000000000000fffffffffffffffffffffffffffffffff98ff9f0fffffffffff
R1[154] <= 640'hfffffffffffffffffffffffffc0090000000000000000000709ff93c63fe480000000000000000007fffffc00000000000000000000007ff3ffffffffffffffffffffffffffffffeffbf8fffffffffff
R1[155] <= 640'hfffffffffffffffffffffffff901f300000000000000000178defd0c73cf640000000000000000007f7f7f800000000000000000001803ff07ffffffffffffffffffffffffffffeefffb9bffffffffff
R1[156] <= 640'hffffffffffffffffffffffffffc0f3c0000000000000000079fe388f7fcf67400000000000000000736ffc000000000000000000028c01fffffffffffffffffffffffffffffffffefff39fffffffffff
R1[157] <= 640'hfffffffffffffffffffffff7ffc0f3c0000000000000000033ff3c8ff7fe7d7e000000000000000003fdf900000000000000000000c000fffff01ffffffffffffffffffffffffffe7ff31fffffffffff
R1[158] <= 640'hffffffffffffffffffffffffff81f2e00000000000000000637ffffeff7fff7f660000000000000007ffd8000000000000006000000381fffff01fffffffffffffffffffffffffff3ff31fffffffffff
R1[159] <= 640'hffffffffffffffffffffffffffe1f6e00000000000000000e17efffeffe7ff7fe0000000000000000f4fdc4000000000000dc6000179837fff76007f7fffffffffffffffffffffdb7ffb07ffffffffff
R1[160] <= 640'hfffffffffffffffffffffffffff0df780000000000000000c7e8d9fbf867fffbd9c00000000001039f3e720000000000000f8000433fc1ffdf800000181ffffffffffffffffffff3fffebfffffffffff
R1[161] <= 640'hffffffffffffffffffffffffff98df780000000000000000004f1fff996fffffc9c00000000000f09f8f7000000000000006000040fcc0fffc0000000001ffffffffffffffffffffffe4bfffffffffff
R1[162] <= 640'hffffffffffffffffffffffffffb8f3f80000000000000000006d7fffc16dffffcbce0100000000f0fecffc0000000000000400000c3e41fff80000000000fffffffffffffffffffffff69fffffffffff
R1[163] <= 640'hfffffffffffffffffffffffffff0f3f8000000000000000007e87fffc0e1ffffffff00000000017fffeffe80000000000000c000010f017ef18000000000fffffffffffffffffffffeff8fffffffffff
R1[164] <= 640'hffffffffffffffffffffffffffb3fff8000000000000000006492fff00e1feeffffe0080008003fb67fffe80000000000000000001c0087fe70000000000ffffffffffffffffffffffff9fffffffffff
R1[165] <= 640'hffffffffffffffffffffffffffbefef9000000000000000000417ff3041ddffffffc8380008003ff677ffe080000000000000000008000831c00000000007fffffffffffffffffffffd93fffffffffff
R1[166] <= 640'hfffffffffffffffffffffffffffffff900000000000000000040fff7063dc7ff7fffc3000000007ffbfbfff800000000000000000000000110000000000003ffffffffffffffffffffd97f7fffffffff
R1[167] <= 640'hfffffffffffffffffffffffffffffff9000000000000000000019fe6e0c933ff7ffff820000007fffbf9ffe100000000000000000000000000000000000003bffffffffffffffffffff9e3ffffffffff
R1[168] <= 640'hffffffffffffffffffffffffffffffffc0000000000000000001ffe748c007fffe77c18330401bfebfffff7f0100000000000000000000000000000000001cf3ffffffffffffffffffefffffffffffff
R1[169] <= 640'hfffffffffffffffffffffffffffffffec00000010000000000003ffecf807cffff3c489070051ffefffffffe6018000000000000000000000000000000000cf3ffffffffffffffffffffffffffffffff
R1[170] <= 640'hffffffffffffffffffffffffffffffffc1010000000000000006fffecf800efffb7ec89800681ffffffffffefc780018000000000000000000000000000001ffffffffffffffffffffffffffffffffff
R1[171] <= 640'hffffffffffffffffffffffffffffffffc0000000000000000007f3e7edf807fefcf7811f00689cbffffffefffe1f6d800000000000000000000000000000011fffffffffffffffffffffffffffffffff
R1[172] <= 640'hffffffffffffffffffffffffffffffffd0248000000000000003ffe7fdf8dfffcee28118900d1fbffffffeffff8f7fe19000000000000000000000000000000fffffffffffffffffffffffffffffffff
R1[173] <= 640'hfffffffffffffffffffffffffffffffff8c680000f00000000037f3c78c01fffdf3c00011e0707bffffffffffecfffffba0000000000000000000000000000007fffffffffffffffffffffffffffffff
R1[174] <= 640'hfffffffffffffffffffffffffffffffffc63800019800000000fff7e79c01ffffc3e00070744c6fffffffffffcfffffffa0000000000000000000000000000003fffffffffffffffffffffffffffffff
R1[175] <= 640'hfffffffffffffffffffffffffffffffff020081cf0800000000effff7fc69ffcf0024000934c06f7fffffffe3c3dfffffe0000000000000000000000000000003fffff9bffffffffffffffffffffffff
R1[176] <= 640'hfffffffffffffffffffffffffffffffff900000cc0000000000ffffe3f7d3fe4600400004d7cdffffffefffc98c3ffffff7000000000000000000000000000003edeb946ffffffffffffffffffffffff
R1[177] <= 640'hfffffffffffffffffffffffffffffffff80000071f3000000007fffefb690fe4400200004dff9ffffffffffe9873ffffff600000000000000000000000000000273f00007fffffffffffffffffffffff
R1[178] <= 640'hfffffffffffffffffffffffffffffffffc0000013cf000000007fffff14186e0000000000fffffffffff7ffe801ffffffc000000000000000000000000000000033100003fffffffffffffffffffffff
R1[179] <= 640'hffffffffffffffffffffffffffffffffff000000fcf70000001ffffff340cf70000000181f7ffffffffffffe0007ffffff000000000000000000000000000000000000001f7fffffffffffffffffffff
R1[180] <= 640'hfffffffffffffffffffffffffffffffeff0000008fff1000003ffff8ffccf370000000091ffffffffffffffc06e1fffffb00000000000000000000000000000000000000067fffffffffffffffffffff
R1[181] <= 640'hfffffffffffffffffffffffffffffffeff0000011ffe80000003ffffffcc7170000000006dfffffffffffffc1c18bffef000000000000000000000000000000000000000007fffffffffffffffffffff
R1[182] <= 640'hfffffffffffffffffffffffffffffffffe8000003ffe80000003ff9fff4800000000008049ffffffffff3fff8007bffe2000000000000000000000000000000000000000001bffffffffffffffffffff
R1[183] <= 640'hfffffffffffffffffffffffffffffffffc8000007fbf81000010fdfffe610000800004010fffffffffffffff80e1bfc70000000000000000000000000000000000000000001bffffffffffffffffffff
R1[184] <= 640'hffffffffffffffffffffffffffffffffff1800016ffff000000177f99f843000000000300dfffffffffd768c80009f9800000000000000000000000000000000000000000018ffffffffffffffffffff
R1[185] <= 640'hfffffffffffffffffffffffffffffffff60000007fffffc000017fffb90000000000000083fffffffffd674c80000fc000000000000000000000000000000000000000000000ffffffffffffffffffff
R1[186] <= 640'hffffffffffffffffffffffffffffffffff000000ffffff800000feff300000000000000003fffffffffdc70181101180000000000000000000000000000000000000000000001fffffffffffffffffff
R1[187] <= 640'hffffffffffffffffffffffffffffffffff060003ffffffc00004fee6000000000000000000ffffffffffd80101003901000000000000000000000000000000000000000000000fffffffffffffffffff
R1[188] <= 640'hfffffffffffffffffffffffffffffffffc060003fffffff8004c1fee0000000000000000003fffffff6d1c01800030000000000000000000000000000000000000000000000007ffffffffffffffffff
R1[189] <= 640'hfffffffffffffffffffffffffffffffffcc20003fffffff0800f9fec0000000000000000013ffffff9490000800000000000000000000000000000000000000000000000000007ffffffffffffffffff
R1[190] <= 640'hffffffffffffffffffffffffffffffffffe30407fffffffb900df9f8000000000000000000fffffff9484000000000010000000000000000000000000000000000000000000007ffffffffffffffffff
R1[191] <= 640'hffffffffffffffffffffffffffffffffff3c4c67fffffff19108db310000000000000000003ffffff1400200000000800000000100000380000000000000000000000000000006ffffffffffffffffff
R1[192] <= 640'hffffffffffffffffffffffffffffffffffffe13fffffffff7c193ff80000000000000000008ffffff8c8002008020000800000000060000080180000000000000000000000000fffffffffffffffffff
R1[193] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffe67fe700000000000000000000007ffffe080000000000000000000008018000000130000000000000000000000000ffffffffffffffffff
R1[194] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffe7ffe700000000000000000000017f7fe600000000000000000000000e0b7100000018000000000000000000000003ffffffffffffffffff
R1[195] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffe6fe30100000000000000000006ffde6000000000000000000000007dd31800000010000000000000000000000077fffffffffffffffff
R1[196] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffefffffffe80000000000000000000004dc660000000000000000000000000dd8700403083000000000000000000000001ffffffffffffffffff
R1[197] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffef88000000000000000000001cc620000000000000000000000000cdce980021000e0400000000000000000003ffffffffffffffffff
R1[198] <= 640'hffff9ff803ffffffffffffffffffffffffffffffffffffffffffff00000000000000000000000c040000000000000000000000000067fffc0000000c0000000000000000000007ffffffffffffffffff
R1[199] <= 640'hfdfe1ffc03f3fffffffffffffffffffffffffffffffffffffffffe90100101000000000000000020000000000000000000000000007c3ffe00040c1c03800000000000000000019fffffffffffffffff
R1[200] <= 640'hfc3c01e0003fffefffffffffffffffffffffffffffffffffffffffe0011000000000000000000000000000000000000000000000001f9f7f103166890000000000000000000041ffffffffffffffffff
R1[201] <= 640'hf8000060003fffefffffffffffffffffffffffffffffffffffffffd881000000000000000000000000000000000000000000000000199fff303f068880000000000000000000497fffffffffffffffff
R1[202] <= 640'hc0000000000e7f00ffffffffffffffffffffffffffffffffffffff9c88860000000000000000000000000000000000000000000000001e7fc0fb604080000000000000000000090fffffffffffffffff
R1[203] <= 640'h4100ffffffffffffffffffffffffffffff7ffffffffe00000000000000000000000000000000000000000000000000003666c4f0e4640000000000000000000349ffffffffffffffffff
R1[204] <= 640'h40003fffffffffffffffffffffffffffffffffffffff0010000000000000000000000000000000000000000000000000020080060f400000000000000000000048ffffffffffffffffff
R1[205] <= 640'h7fffffffffffffffffffffffffffffffffffffff3123000080000000000000000000000000000000000000000000004000ccc000000000000000000000034dbfffffffffffffffff
R1[206] <= 640'h7fffffffffffffffffffffffffffffc17ffffffff903000000000000000000000000000000000000000000800000000000c0c00000000000000000000007491fffffffffffffffff
R1[207] <= 640'h3bffffffffffffffffffffffffff7f387ffffffff80000000000000000000000000030000000000000000800000000000000000000000000000000000000c9fbffffffffffffffff
R1[208] <= 640'h3bffffffffffffffffffffffffffff30cffffffce01000000000000000000000000600ff000000000081ff00000000000000060000000000000000000004c1c0fefffeffffffffff
R1[209] <= 640'h1bffffffffffffffff7ffffffeff7ef08ffffffff68000000000000000000000000fffff7f000000feffffc000000000000000000000000000000000000018007fffffffffffffff
R1[210] <= 640'h3ffffffffffffffffffffffffff78000ffffffff0800000000000000000000001ffdffffff80000ffffffe60000000000000000000000000000000000000c007fffffffffffffff
R1[211] <= 640'h3ffffffffff77ff7efffffffffce000077f7fff80000000000000000000000003fbfffffffc0001fffffffe0000000000000000000000000000000000000101ffffffffffffffff
R1[212] <= 640'h187ffffffff2480f8fffffffe7dc00000ff7fff00000000000000000000000003ffffffffffef03ffffffffe0000000000000000000000000000000000001007effffffefffffff
R1[213] <= 640'h87fffffffc100178fffffffeff000000fefffe0000000000000000000000003ffffffffffffefffffffffff8000000000000000000000000000000000000000e3f7fffffffffff
R1[214] <= 640'h7f7fe000000000fffffffff000000000ffcc0000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000000000007e7fffdfffffff
R1[215] <= 640'h3c18c0000000000ffffffec00000000018c000000000000000000000608c7fffffffffffffffffffffffffe000000000000000000000000000000000000000c3f3ff57ffffff
R1[216] <= 640'h1800000000000000600000000013fffffe000000000000000000000000000000000010fffffffffffffffffffffffffffff00000000000000000000000000000000000000420247ecdffffff
R1[217] <= 640'h1cc080000000000000000000000fffffcc000000000000000000000000000000000007fffffffffffffffffffffffffffff2000000000000000000000000000000000000000000ece5ffffff
R1[218] <= 640'h11c07c00000000000000000000007fffd000000000000000000000000000000000003c7fffffffffffffffffffffffffffffe800000000000000080000000000000000000000000fdb7ffffff
R1[219] <= 640'h3ff1ff80000000000000000000003ff78000000000000000000000000000000000000cffffffffffffffffffffffffffffffff800000000000000c30000000000000000000000005f96ffffff
R1[220] <= 640'hfffcfc0000000000000000000003bf480000000000000000000000000000000000008efffffffffffffffffffffffffffffffc000000000304003fe000000000000000000000005fc6ffffff
R1[221] <= 640'h8fffefc0000000000000000000003fec10000000000000000000000000000000000041ffffffffffffffffffffffffffffffffec00000240700787fe100000000000000040000003fb6ffffff
R1[222] <= 640'h8fffffe0000000000000000000003b0000000000000000000000000000000000000071ffffffffffffffffffffffffffffffffff0f800668f87feffe100000000000000040000001fb279ffff
R1[223] <= 640'h40c0fffffff00000000000000000000003300000000000000000000000000000000000003ffffffffffffffffffffffffffffffffffffff0067ffefffff7c00000000000000000000000eb27fffff
R1[224] <= 640'hbfffffffcc300000000000000000000000000000000000000000000000000000000000feffffffffffffffffffffffffffffffffffffffeffffffffffff8000000000000046c200002f925ffffd
R1[225] <= 640'h1ffffffffeff0000000000000000000000000000000000000000000000000000000000037fffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000ea600002f145b6dfd
R1[226] <= 640'h3ffffffffffff0f000000000000000000000000000000000000000000000000000c0000c7ffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000026b200013f922bef7d
R1[227] <= 640'h1fffffffffffffffe0000000000000000000000000000000000000000000000000188303e7fffffffffffffffffffffffffffffffffffffffffffffffffffff00000000000012b2200013f486fdb7c
R1[228] <= 640'h3fffffffffffffffe000000000000000000000000000000000000000000000000000c37ffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000001262c000139fa2cd37d
R1[229] <= 640'h183fffffffffffffffe0000000000000000000000000000000000000000000000000c1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000b3390001393908b579
R1[230] <= 640'h3e3fffffffffffffffff800000000000000000000000000000000000000000000100ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000086b800018eb6d15bd
R1[231] <= 640'hffffffffffffffffffffe000000000000000000000000000000000000000000001467ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000f658000964a0919bc
R1[232] <= 640'hff7ffffffffffffffffff00000000000000000000000000000000000000000003003fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0000000000027c800122f068f9f0
R1[233] <= 640'hfffffffffffffffffffff80000000000000000000000000000000000000000002003fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000f0b2980328f93bf934
R1[234] <= 640'hffffffffffffffffffffff0000000000000000000001000000000000000018000101ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3ca000005fb6a005b07a33b368
R1[235] <= 640'hffffffffffffffffffffffe000000000000000000001000c0080000000003c00effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee00080e689900195735b7bb6
R1[236] <= 640'hfffffffffffffffffffffff80100000000000000000307fffcc0003f0000fc00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8e2886fe5c0019d24044bf0
R1[237] <= 640'hfffffffffffffffffffffff90300000000000000000007ffffe31fffc000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff648830f3a0009639ebf7bf
R1[238] <= 640'hfffffffffffffffffffffff967e0000000000000000001fffffffffff01efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc401a3be080af590ebcbd
R1[239] <= 640'hfffffffffffffffffffffffff8f8200000000000000800ffffffffffc01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec1065a5e615af194936c6
R1[240] <= 640'hfffffffffffffffffffffffff3fc00000000000000000fffffffffff80ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe430ac418044cfb40b36cf
R1[241] <= 640'hffffffffffffffffffffffffffff000800000000001e1ffffffffffd80ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc4e173a97a2405f033a7fb
R1[242] <= 640'hfffffffffffffffffffffffffffffafc00000000003fbfffffffffffc3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe4d3379aea26ebf909bf7b
R1[243] <= 640'hfffffffffffffffffffffffffffffffe00000000003f9ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff46139bcd5718f59437ab1
R1[244] <= 640'hffffffffffffffffffffffffffffffffc0800003843ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd9fffe0397d1c9eb7d0102ddfd7
R1[245] <= 640'hffffffffffffffffffffffffffffffffe18c017fc63ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffd9fff7145be788b738014fd4ded
R1[246] <= 640'hfffffffffffffffffffffffffffffffff3feffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffff9fff75fe59315b5ad81ca9def1
R1[247] <= 640'hfffffffffffffffffffffffffffffffffbfffffff37ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffff9fff46d53c99ceec4a0458c397
R1[248] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc9fbf72e21b2c9fcde3b609ef0e
R1[249] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffafff91fff2d3c7e91bb5c59d43536cf
R1[250] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbffdbfffb6889bbb9b1c478ac75c1d
R1[251] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5b3cf7b3f3b066b90201e96f07f9460
R1[252] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f3ed333f348be387941e6187610c01
R1[253] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbd765237fecbcb1a5b54dbec165abc4
R1[254] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff26fb4ebffe7d93bb6dbc9f76ccf6483
R1[255] <= 640'hfeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa725c12affb09386a1457bf315cdad35
R1[256] <= 640'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee16a90baffbab5b50b1ac3fcc8d73a7a
R1[257] <= 640'h83ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff644f9dddf90a0f78a16e78efb05358f1
R1[258] <= 640'hc3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff72906495fffb080252bfcaf8e55aedb8
R1[259] <= 640'hf7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe993abc4179888f29855c5e7f37707968
R1[260] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff564156f97881624484e7267f9b1534d0
R1[261] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff77aa2f8f879db0ded855be972e659b585
R1[262] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb1ffcfff3d9dbb74eace7cf9c8f0cf3bb
R1[263] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddcfbfc297dbb78aef7593e5c4f4472543
R1[264] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedf7c14fbf7bbcd8a10ced1ace63b09882b
R1[265] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefbfdecd8277af0dbe5219555fe7927c3ee
R1[266] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedbffdcf78ad6e2c7a3f9b8fb7fed92dc7f
R1[267] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffcbbfee86e6643a3a8365762fe18baa43
R1[268] <= 640'h3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff77e7b3738fec5f2e6d6b167cd7d50d9d6c
R1[269] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffb123d5dd9be67e2a2dcf42d81f8d55
R1[270] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe79d973e263dcba9ef6af69514ec3b746aa
R1[271] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4fefcb53f3aa7d0bbf67ee33ffe007fb1a
R1[272] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddf18abed79277bb95ed909a7ebcd7e3bc
R1[273] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffba6fddeb2dffebfc6486325367a8b5fdbbb
R1[274] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfe7443d79b7bfe67f2f1f8ce7d9c8bf9a7
R1[275] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7e6f4fb6ce2e67b01fe2bd1e3db4029949
R1[276] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa7337e9edd4e38fff67ee3decffd2acea93f
R1[277] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7bd3fcef141f9cc7f1ee3f033f9f2d3f325
R1[278] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdd33fc71cc13fda5e51d61fee69e74e11a1e
R1[279] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdefeb95fcd45bff7fcebf7e666f75d8da3d3
R1[280] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb6479d40e977deecce6663af2deb6b3c48
R1[281] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef993f4db08c359d3dc761bd29c37fa30f0f
R1[282] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff719d33677cd53d2ffaf765c199edf9ec79e9
R1[283] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfbdcf17583fbe37fab6167e7d7fc4ed460
R1[284] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeb6fe6f605e97c7e2ff33f7d835d3e9e4d6a0
R1[285] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefb96678244c9b7b3fec8a6c0b709fff271f4
R1[286] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fe9b3d72485b5ffbf36f285254973f263bd
R1[287] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffee7ff4fdee44c5f766bffd621f9b6cc6c13533
R1[288] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7eee32fea5610df4fffdf53af997671e48671
R1[289] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff37fcd7f77f105be0fefb7236db7a8e3e17485
R1[290] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fb3b9af5fbf57efb7effa26ae8c4f7df37ffb
R1[291] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbbdab07660dfbfbaf7b011e62ce8e1b08fd
R1[292] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffde7de7f361bd701fe49fe0c0bf6b6f96f0ba74
R1[293] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6d74becfe8917daf3fd885658e6bb7f87e5c
R1[294] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6e72fada7fedafbbb67cba71e477fab78cacf
R1[295] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff33d32e3b038be5ccf369855e99f345583cdf
R1[296] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb157f868d7f590fe0e9ede5df3b773978797a
R1[297] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3a9af661d390ceffc9e7a7e5deeee6bc7bad
R1[298] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffef482244cb789b07e94f4d799fc5ec6fcf95d
R1[299] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb09455b6c6417ff6e6fd8751f77ccfc89987
R1[300] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6eb49ad76f0886ed2fb796777ce3afdcd69e3
R1[301] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff02ef27dde007f7aef9be177a313fe7df9bc
R1[302] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fffffffffff718d6b634f98bcf3feb9b22eb99def9ac31ec
R1[303] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3fff3ffffffffffffffffffffffffffffffffffffffffffff1ffffffffffffe6fdb9bc168cece463f5f2dbbf96b598be7c
R1[304] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1ff007fffffffffffffffffffffffffffffffffffffffffffdffffffffffffd73210546740bdee3ffa71de6bb3efdcf9fb
R1[305] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc01f8037ffffffffffffffffffffffffffffffffffffffffffb1fffffffffff3c630f8a96627bb5f2db1733ffbd5afcc59e7
R1[306] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe003f003ffffffffffffffffffffffffffffffffffffffffffff3fffbfffffedbf0df16d2260273ddce3063e9eba5e7f0fb3b
R1[307] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff900ff003fffffffffffffffffffffffffffffffffffffffffff9214a2ffffff6ffc2634609664fefb9b6f327bbf07fff1da04
R1[308] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe403e0003fffffffffffffffffffffffffffffffffffffffffff98dfffffffff6fff9257319861b75f896ff0ff3fce6ef8ee82
R1[309] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff803f00011fffffffffffffffffffffffffffffffffffffffffff9ffff3ffffffb9ffbaec7840138ffd9679a04bffb7adf8e4f6
R1[310] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1fe04000fffffffffffffffffffffffffffffffffffffffffff9fffdfffffffffff397c9ece8337fb9bb2c0b2fb359ffc6cff
R1[311] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0180007fffffffffffffffffffffffffffffffffe3fffffffb5ffffffffffdfff76cdeceec6fff3db5791ceffdfd8fddcfc
R1[312] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff860037fffdfffffffffffffc3fffffffffffffffe3ffffffff8bffbfffff7bbe7ee486626e2bfff9563b39ffef6eaf87c18
R1[313] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000c007ffffffffffffffffffffffffffff043fffffffd8fff3fffffcbbfb5fb8c739a1a7bfdf6fc37fdfef3f7c36a7
R1[314] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7c00000000801ffffffffffffffffffffffffffff8387fffffffcbdff3fffffc9fd9fecc5118e37629fb7bc0fedfd94fbc50f7
R1[315] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffff800fe3fdfffffe01fffcfffffffffffffffffffffffffffffffffffefff77ffffffbdcffa5349d8a18f65d7cce2ceff3d678e6ce9
R1[316] <= 640'hffffffffffffffffffffffffffffffffffffffffe3ffffffffffffffffffffffffff000ffffffffffffffffffffffffffffffffffffffff6ff37ffffffbcffdab25ce8b254cf50e04a9df7793ef46d16
R1[317] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0007ffd3fffbfffffffffffffffffffffffffffffff5fff77fffef5ffbfdb0ee2e059cb73bf8c3d85fc63eec4ca9
R1[318] <= 640'hfcf03effffffffffffffffffffffffffffffffffffffffffffffffffffffffe773ffc07fc0fff80ffffffffffffffffffffffffffdf3fafffff79c77bfacab32e3dcb41fffa97ede953bec48ca
R1[319] <= 640'hf7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffff048f887ff0017ffffffffffffffffffffefff6dbfdfffff76726ffda6990909fc7b7f7cbed59a9bfd49b3c
R1[320] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff17ff00fe0007ffffffffffffffffffffbefee99bff7fff9b7bbbd0b33e8119ff62bf601b3519bbff67679
R1[321] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffa00f0000fffffffffffffffffbfffdffff47ad3fffe9eb7e5cd67b002979e78ff409f1db89fe878f5
R1[322] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800ff00ff3fffffffffffffffbffbdfb2efcdf3ffff25df6bc5209860b6773db3803d77f66ede2ceb
R1[323] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1b7fff7ff91ffffffffffff7eeed5fbe5af5b3fffc30d6ebaa4c885406ee62b281217f4f4ef656d5
R1[324] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffffc7ffffffffff93febffe9a157f7bfff6bf817f904b047c2cb4532781637f712cd8fed7
R1[325] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb39686b7cd5f7efbffffa7914f9f1bc65c94ff366e035b7bd347d662a2
R1[326] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb3a6e373ff6ccd89fffe7773ee2c54fe2413170c2e811afff9af143642
R1[327] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff874c0fb880ffffffffa3f6ab1bf64f9b33dff7bf3e33f766737a21d200dc08b35daae5f854cc
R1[328] <= 640'he3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0bffffffffffff51ff9ddfbc3c2afbdfdee9de68a3d2913e42906dd6408fd35db1fa1d49
R1[329] <= 640'hfffffffffffffffff8f0fff8fffffffffffffffffffffffffffffffffffff9e3fffffffffffffffffffffffffffffffffffffffbdb5b9fdc39cdfbd6fffbdbbfcbe27e121219776ec83da7b6f9fc6fe9
R1[330] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffb0fdff42451e7d7ed57f7ccd3357f12977add7a502562917d6272f5
R1[331] <= 640'h3fffcfffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff4bf60ecff638ef899f7ffdf2e77fc9ebac710a71de403a47e199f05b9f
R1[332] <= 640'h3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed3ef0b0bff2d97b9bffedbe7fbdd9d491295b737ddc12afe7d484c7ab7
R1[333] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe5bef3d9bff7f8f9dfbfbaf5b4b5fdf9d98cbc7927c003b2f737a7c6ebb
R1[334] <= 640'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe8ecd5703fef1bbab7ff9a35f1e6cefec9c6c6049bf00bfeff9fe243ed3
R1[335] <= 640'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed5fb6bc7bf7db7c87de8da77ddb8a3f9840e31ec7dc42b7ff1fdae6a35
R1[336] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6ef3ff7ff9bdbfcee6b17a63b5e5ef3c8627d6deff804f3f9dfdb459b7
R1[337] <= 640'hf7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff2fe0ed7fef0b3a77ffbcbb69add0b776063104ecb588677fcbfb3e4b1b
R1[338] <= 640'h1fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebe687adfed2b4ebbfdcfdd4dff2c5a743570ae6518c77bcedbcfe3a59
R1[339] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf83e508ebd6d7bddbafb4d23cfeba25d763184dfe6c587bfdfddfec3cb3
R1[340] <= 640'h800001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdec6e7aaeff7fc7977dfff956ec5a8f3f3e293c035b1cc7d3cfdecc6267e
R1[341] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffefe44d257b9fe96739cf7abfcf3bd074de44b10c22ef467ee571f5f77d3c
R1[342] <= 640'h800001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefcb7b7e6ef3f8ff586ffefcef5facc9740230e90ded867fdbddaff77b6c
R1[343] <= 640'h1500001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3ffffffffffffffffffffffedc85a15b5ffd8a7fef0cf5f877fc70332b811ca409278a1d4cff5ef31f1e
R1[344] <= 640'h40001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffffffffffffffffffffffccbf7f4f3cefd484eeddffc88f9fba0a0fda9c9bb27a19f1db8714a13367e
R1[345] <= 640'h30000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffe764dcddb47cbf4dfdbddbb78d9ebfc7d3c9119c835c9f259bf9383c1a6f
R1[346] <= 640'h20001ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fffffffffffffffffffffff4ff25f9f1ea6b89dfface59f35af61fa78e9d8f83cb40f2e7e3abb78302e
R1[347] <= 640'h30003ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfffe6ffffffffffffffffffb70773bf5d1fb15fb769ec7b6eb5fb7c562cc2e819321016771bb7e20b1e
R1[348] <= 640'h3000000c1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8ff9fff9cfffcebffffffffffffffffff6f0db1efec6e4cb7f3bfaf95efffeee0060086029b90e8675734eee197b
R1[349] <= 640'h30000000000ffffffffffffffffffffffffffffffffffffffffffffff9fffffff9b82fffffaadfff7bbffffffffffffffffcf97caa6a7fec02ffb7fdf7a7f8fb33d7f50ce1c92b32e94c201972c28fd
R1[350] <= 640'h80000000000ffffffffffffffffffffffffffffffffffffffffffff7f0fff0feb93d77ffffc2ffffdbbffffffffffffffff85afdfdcd7b7516f7677fd73eeedffaea7c8561c62c45f8ff011ee6235fb
R1[351] <= 640'hc0000000007ffffffffffffffffffffffffffffffffffffffffffffffffffff45f0b7fffff412ffe4f9ffffffffffffffff9bcf5d3bd369629fe9dbfdf8efac2bce57a884062bdc22427873189c1def
R1[352] <= 640'h37fffffffffffffffffffffffffffffffffffffffffffffffffbe64747efffff61fffa6f9ffffffffffffffff49e1956f95d735f79cb57ffd7e7b9bb913d041933ef86503d84ece28694f
R1[353] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffb692f29fffffb7fffeef9ffffffffffffffff7bd83d7b9ef7e8b7dff7be6bfe6df9b19dd8078a8d0843828311beda0e91
R1[354] <= 640'h7efffffffffffffffffffffffffffffffffffffffffffffffbff4c9ffffff9cfffffffffffffffffffffff9ded9799d7576593df7ef759febde66a4dec090743ad29014b228e64322d
R1[355] <= 640'h3ffffffffffffffffffffffffffffffffffffffffffffff7fcdf7eefffccfffffffffffffffffffffff4efd8f7c9bbbc6bbe77db977ebff741f69626503b1be1be32103cddc3e1c
R1[356] <= 640'h381fffffffffff0001ffffffffffffffffffffffffffffffff7dabdafffbecffffd7fffffffffffffffffeceebcdfcfb4f0ddeff7eef7dda0a39ed3860381d96a6842118fd8f8377e
R1[357] <= 640'h200000000000001fffffffffffe000083fffffffffffffffffffffffffffffff7a91bccff9a7e7ffdb7fffffffffffffffffff7effe5612e3ddd9df7dedc83f61a342550200b4ee26023086c9bc3e30
R1[358] <= 640'hf01ffffffe0000000ffc003ffffffffffffffffffffffffd9e7ebccffd9fe7ffd7bffffffffffffffffb7a6ced9bb752bdfdfdf635ff67b7ac9f5350202461ae4301002336e7c31
R1[359] <= 640'h2000000000000000000001b9c00000000000e381ffffffffffffffffffffffdf3a47f597efc7ffff35bffffffffffffffffff98ddedfcbff2ff3fdfde7ee23f5eec2aa100014624c9f033019e742500
R1[360] <= 640'h2084000000000000000000000000000000007fffffffffffffffffffffffcc594bfdffef68fbff5bbfffffff7fffffffffeda7fd7f69accdfbebfdbf9d6a7386f866700c2c03c90303300eff26000
R1[361] <= 640'hc2429000000000000000000000000000000007fffffffffffffffffffffffee4ac3f9dec282f3ff37f7ffffff7ffffffffbe7e7ff9fff6ebb6bdfbed7fc71caf227a0e80601814d03026604e864000
R1[362] <= 640'h210004000000000000000000000001000000007ff877fffffffffffffffffff5312f3bddcf60e7ff377fffffff7ffffffffdfc8a713fb7796fdbecfe97341bac6afff0fc1407415163002c410e43e00
R1[363] <= 640'h100000880000000000000000000000040000000001fffffffffffffffffffff9d9ff4bf9f1f3f2fd3f7ffffffffffffffdfff7e67ee7fdf7debdc37fdfbdfeb8c5991d3c1e0ea017a3004c003c31200
R1[364] <= 640'h70003040000000000000000000000000000000001ffffffffffffffffffffffcca27ff96d574f7fd737ffffffffffffffeffbfeef3427faeecee47f1d35cbedda6230cf40b07909622000c018260008
R1[365] <= 640'h300000d0030000000000000000000204000000001ffffffffffffffffffffe778e1e7fd1f7ebb7fdff7ffffffeffffffffeefec237fca6de385e776fde665ee5bf0100300a03d00ba0000c000200000
R1[366] <= 640'ha00000601040000000000000000000070000000000769ffffffffffffffffffd8f4fffb36eefb2ff4bfffffff6fffffffeff3fde37666dc72c9f773dd9b667c3ee006168000140198000040c0020203
R1[367] <= 640'h180000014806000000000000000000104000000000006c7ffffffff7fffffffebd796704f6bd9f7f64bfdbfffff7fffffff7db7696afbf5b26cbfbcbfd9cf26ece88170810901a810920000003821061
R1[368] <= 640'h2740c000000000000000000500000000000e11ffffffffbfffffffdb68a47987eed8d9feeff8ffffff7f7fff7f7d93ee2fff667a3e7fabdfd369677df283a29f0c47281be00000000fe00e8
R1[369] <= 640'h469c80640040000000040780000000000000ffffffe72ffffffbdc2bb319a7fa9fe93eb9d8fffff7ffffffffffbec9d5a6df7e26fe474fc5a237b85a031d450005d01fc8000000131388c
R1[370] <= 640'h8c2a1800100000000006000000000000000fffffe33fffffddeb2e1b45059a9fe9fe9f7dffffff4fffffffeffd1eb25edfab0ffcc6efdf3e3ddaf8237182800070005800000017720e0
R1[371] <= 640'hc0005c272100000000000003300000000000000ffffffa5fffff9cf7d4f0cd1fe01fcdbe5dfdffffffbffffbfe6db6d968dfbed79e6ddfe7dbe1c43f9439df57800040054060000006200e8
R1[372] <= 640'h400000302c20400000000c00ae1c0000000000ffffffce27ffeedf58c9f29d6db295c58ecbfffffffff7f7f9b6fbf9e32fffbb6b9f7f0bd79faf827334985fb000000005114000000340008
R1[373] <= 640'h1c0000008010000000000800200000000000000ffffffc87feed8d3071f6b2f3e256cffe199cfffff79667ddfffe7fea0b6f7bf9bf77dfbfb73bcedd000a4f3800000002a1a000000620002
R1[374] <= 640'h3e000000451000000008000000000dc00700f3fffffb497feff722ec62e22edf846896c9b7dfffff9fffffbdfbe21f6c6dafff90fe7dfff96e1fe7e0c9fd9268000238301d00000040000c
R1[375] <= 640'h3f00000029000000000000000000000000fffffffca2e57ff8fa3d8d24ed6cf97fcd76c87f7ffffdefdfffff3d95ebc8f76e5d17ebd7ed9db8deb80c0fc4800001028001a02000002000d
R1[376] <= 640'h107e00000100b00000000000000000000ffdfffffe6a8dfff8fa778c25efd9bbfbe5f449367ffffee3bffdbe3f1ce9dcbdbf86b35cd5968b7ebb8200945f2c00000280018000000000009
R1[377] <= 640'hfe00000060080080000000000001ffffffffe8e82a6cd0b4a7cfaa7ebb3b916fdeedf67fffffefffffdeff18b9e576d180baaff31eb3dcd0380000981b003005c0004000000000008
R1[378] <= 640'h1fc000021d8078000300000001ffffffffff0277d42e686a7de5dc0a93dd3d57afeeeffffff67ffff7e339534214f7c3cee7bef8c3ca463fe1866c81780300440000000000000000
R1[379] <= 640'hef0003fc00001400c000100000007ffffffffffb364b3a57908a8a1b4466dfdd4f7b7ff6ffffdfb77ffbff3761491c8aa47a9df32bfe3b5fa27fd87d208b80000000000000000000000
R1[380] <= 640'h37fc0011f0000208800013000007fffffffffffb33f812bf3adf027bd69e7dcbdbf7a6ffffffffd7ff7bff1c800008000779b1be2e3d92e36f4dfc35844400000000000000000000000
R1[381] <= 640'h603fe0007e000114000130087fffffefffffff5b3000f764a51fdfbb3996fb89ff971efffffffd3ffedff160000000006ae9c9ff7dd6051ee8d5e26608000000000000000000000000
R1[382] <= 640'h19007f0000c000000001ffff7ffff7ef013ffeb38847ebe906858c7f372ddce46fc51cb7ffffae3ffffff200000000000100ffdd7e5549fc48dfe06200000000000000000000000000
R1[383] <= 640'hf80066dc00178000003fff7fffeee7010efffb91657eec761cf659e7fb320527da45d6e7fffe72f6f7ddc0000000000007b31bf7d7c06e25ed7600000000000000000000000000000
R1[384] <= 640'h4f000003c0007000001bcbff8800c3c02ffff873d0f9afb243833dd5f77e11613c6bd7e3ffff36f7f78c000000000000001ddfffdd81c63c91f000000000000000000000000000000
R1[385] <= 640'h307fc000000640fc000001ffc00000483fffb9bb15b0cf9b8af4ae4be2cfe16a7c72dfffffffe5e7f020000000000000001e65b5a8c17e2ea9e000000000000000000000000000000
R1[386] <= 640'h1f01ff8000000f000000007360000063fff6b8361892bfda72f64eb9a396f21a2cd2c3bfffffb5ac55000000000000000000e7f7b967c8d1b18000000000000000000000000000000
R1[387] <= 640'h3800fff8000003818dc000edf0000fffffe828b45ffe7f8e6ad343be7623ce79f50e0ff7f24046736000000000000000000000003287f3d6e0000000000000000000000000000000
R1[388] <= 640'hfe0001effff00b8c89c6837ffff3fffffb8793945aaface3d27677f6d29fa798d3c068032fb3fda800000000000000000100000000003c100000000000000000000000000000000
R1[389] <= 640'h6fe0000000ff81f0000800dffffff3ff8000398ed5fe5704d0236fc0099eb1f7f9d506fff5ffe5b0000000000000000000000000000000000000000000000000000000000000000
R1[390] <= 640'h31fff8000000fe00260400bffffffff90000000004052549ab7bdf94f6220010bb67bfe3f7f58e00000000000000000000000000000000000000000000000000000000000000000
R1[391] <= 640'h1c01ffe8f9940bf98199002ffffffe7000000000000b5c421e808a0ee40000187f4e9ccce00fc000000000000000000000000000000000000000000000000000000000000000000
R1[392] <= 640'h7c00fcfe7fff80e7f00000bffffe0000000000000003a99e90eb181e000001ffd147c0000000000000000000000000000000000000000000000000000000000000000000000000
R1[393] <= 640'hf800100000fff001e800028ffff0000000000000000046cfbdf9ce0000000000ce000000000000000000000000000000000000000000000000000000000000000000000000000
R1[394] <= 640'h3f8000000001ffe3e07c006e901000000000000000000e8e49a670000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[395] <= 640'hffcc00cc300ffff008000118000000000000000000005186c840000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[396] <= 640'h3fffffffff038ffc00100000000000000000000000000340000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[397] <= 640'h3c07fffffedffd803fe0410000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[398] <= 640'hfe07ffffc00fff8c07f988018000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[399] <= 640'h1fce3000f0001bffe07741800000000000000000001bc0000000000000000000000000000000000000000000000000003000000000000000000000000000000000000000000
R1[400] <= 640'hfffffccffff801fff6000000000000000000000000410000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[401] <= 640'h33ffffffffffe0006f800000000000000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[402] <= 640'h381ffffffffffff806df0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[403] <= 640'hf86ffffff003ffffc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[404] <= 640'h3fe00e30000003ffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[405] <= 640'hfffff00707000000ffc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[406] <= 640'h3ffffffffffffc0007fe00800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[407] <= 640'h3fffffffffffffff43b30200000000000000000020000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000
R1[408] <= 640'h11fffffffffffffffde00040000000000000000000000000000000000000000000000000000000000000000000000000001900000000000000000000000000000000000
R1[409] <= 640'he0fffe81c3003fffffe0000000000000000000000000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000000
R1[410] <= 640'h79788381e3ff0071fff8e3c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[411] <= 640'h3ffffffefffffef93f00f06000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[412] <= 640'h7ffffffffffffffffe0180018000000007800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[413] <= 640'h1ffffffffffffffffffdc0400000000001600600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[414] <= 640'h707fffff8ce60fffffffe3800000000006c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[415] <= 640'h3f7124c00fefc7ff3c2e8060000000000090000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[416] <= 640'h1ffffffffffffffffffe3818282000000024000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[417] <= 640'h3fffffffffffffffffffffe780000000008800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[418] <= 640'h7fffffffffffffffffffff780000000003700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[419] <= 640'h1ffffffe01fe7ffffff99080000000000cc0180000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000
R1[420] <= 640'hc80073effffffffffff7ef80000000000130060000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[421] <= 640'h7ffdffffffffffffffffff8000000000006a01c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[422] <= 640'h3ffffffffffffffffffffff000000000001c806000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[423] <= 640'h7ffffffffffffffffffffbc000000000007300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[424] <= 640'h1ffffffffe7ffffffffffff000000000001840000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[425] <= 640'h30ffffffffffffffffffffe00000000000398000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[426] <= 640'h147ffffffffffffffffffff000000000000e2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[427] <= 640'hfffffffffffffffffffffffff8700000003f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[428] <= 640'h3fffffffffffffffffffffffffe0f8000004000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[429] <= 640'hffffe9ffffffffffffffffbffff00ff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[430] <= 640'h1ff3fe77fffffffffffffffffffffc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[431] <= 640'h201ffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[432] <= 640'h3ffffffffffffefffffffff00c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[433] <= 640'hffffffffffffffffffffff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[434] <= 640'h3ffffffffc3fffffffffe000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[435] <= 640'h7fff00833fffffffff00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[436] <= 640'h2e01ffffffffeff0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[437] <= 640'h681fffffffffc000000000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000
R1[438] <= 640'h1ffffffffe100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[439] <= 640'hffffff180000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[440] <= 640'h3efc00800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[441] <= 640'hfc300000000000000000000000000000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[442] <= 640'h78000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R1[443] <= 640'h0
R1[444] <= 640'h0
R1[445] <= 640'h4000000000000000000000000000000000
R1[446] <= 640'hc000000000000000000000000000000000
R1[447] <= 640'h0
R1[448] <= 640'h7f0380000000000000000000000000000000000
R1[449] <= 640'h180000000000000000000000000000000602000000000000000000000000000000000000
R1[450] <= 640'h80000000000000000000000000000000003800000000000000000000000000000000000
R1[451] <= 640'h80000000000000000000000000000000000000000000000000
R1[452] <= 640'h180000000000000000000000000000000000000000000000000000000000000
R1[453] <= 640'hc000080000000000000000000000000000000000000000000000000000000000000
R1[454] <= 640'h1800000000000000008000000000000000000000000000000000000000000000000
R1[455] <= 640'h60000000000effffc3000000000000000000000000000000000000000000000000
R1[456] <= 640'h1c000038f3e1820000000000000000000000000000000000000000000000000000
R1[457] <= 640'h200000000000000000100000187ffc00d0370020001000000000000000000000000000000000000000000000000
R1[458] <= 640'h6000700c08000000000000000000000000000003c000025000000000000000000000000000000000000000000000000
R1[459] <= 640'h9f30040800000000000000000000000000000000000000000000000
R1[460] <= 640'h3fffc64800000000000000000000000000000000000000000000000
R1[461] <= 640'h8001ffffe5800000000000000000000000000000000000000000000000
R1[462] <= 640'hff8003fffff7eb6000000000000000000000000000000000000000000000
R1[463] <= 640'h1000000000000000000000000018c0001fffff7ef7f00000000000000000000000000000000000000000000
R1[464] <= 640'h24008000000000000000000000000000000000200000007ffff7ef7fc0000000000000000000000000000000000000000000
R1[465] <= 640'h10000000007ffe3ef3fe0000000000000000000000000000000000000000000
R1[466] <= 640'hfff3ee1fc6000000000000000000000000000000000000000000
R1[467] <= 640'h4000000000000000000000000000000000000000000
R1[468] <= 640'h100000000000000000000000000000000000000000000000000000000000000000000000000000000007f9dfbfe7c00000000000000000000000000000000000000000
R1[469] <= 640'h40000000000000000000000000000000000000000000200000000000000000000000000000000000000001d972ffff80000000000000000000000000c00800000000000
R1[470] <= 640'h2000000000000000000000000000000000000000000000004c000000000000000000000000000000000000000004b9ffffc000000000000000000000007f800000000000000
R1[471] <= 640'h20000000000000000000000000000000000000000000000003c0000000000000000000000000000000000000000001fffff00000000000000000000003f70e0300000200000
R1[472] <= 640'h400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001fff800000180000000001c08fffb0f13c0026000000
R1[473] <= 640'hff8000000000000000000000ff810000006000000007f38ef88000800010000000
R1[474] <= 640'h8000000000000000000000000000000000000000000000000000000000000080000000000000000000000080000000000000000000000001c0000000000000000ef00c01f000000000000000
R1[475] <= 640'h60000000000000000000000000000000000000000000000003800000000000000000000010000000000000000000000000000c0000000003f3ffff007ffe000100000000000
R1[476] <= 640'hc00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007ffbfd1168fc000040e0000000000
R1[477] <= 640'h200000001c0001f0000000000000000000000000000000000000000000000000e13f0f9a00fec000b000060040000000
R1[478] <= 640'h20000000000001800000000000000000000000000000000000000000000000000125f8800ff00010000000004e040004
R1[479] <= 640'h2200000000000000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000000000000000000000000000ff000000000000000000e0400
end
always @(posedge vga_clk) begin
R2[0] <= 640'hffffffffefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[1] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[2] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[3] <= 640'h7fffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[4] <= 640'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[5] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[6] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[7] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[8] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffff7ffffffffffffffffffffffffffffffffff7fffffffffffffffffff
R2[9] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[10] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[11] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcfefffffffffffffffffffffffffffffffffffffffffffffffeffffffffffffff
R2[12] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffef8fefbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[13] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefcbff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
R2[14] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1ff7fffffffffeffffffffffffffffffffffffffffffffffffffffffffffffff
R2[15] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7f7ffeff7fc7ff96ffffffffff3fffffffffffffffffffffffffffffffffffffffffffffffffff
R2[16] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9ff9fffbffc7e1f1ecffef97f3b7fffffffbffffffffffffffffffffffffeffff7effffffffffff
R2[17] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9ffffffe7e1f3ffffffb7ffb7bfffffffdfffffffffffffffffffffffeffffffffffffffffff
R2[18] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffff9fe00c13f3c9f19fcf973f8ff7ffdffffffffffffffffffffffffffffffffffffffffff
R2[19] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc03e00c0e138df90fffcfbf8fffffffffffffffffffffffffffffffeffffffffffffffff
R2[20] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6ffffffc33f00c00001fe900f9cf1fcffff3fffffffffffffffffffffff7bffffffffffffffffff
R2[21] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffeffffff67ff00800083fc11071900fcffff7ffffeffffffffffffffffff7fffffffffffffffffff
R2[22] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9ff777f66610000008600010331000099cffefffeffffffffffffffffffffccffffffffffffffff
R2[23] <= 640'hfffffffffffffffffffffffffffe7ffffffffffffffffffffffffffffffffffffffdfeff66efdec799ff6778600000003186000080f18700998f76ff1fffffffffffffffffffdfff7ffeffffffffffff
R2[24] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbffefffe33c79c7c8c0000000010000000000990000fe0f3bcfc7fffffffffffffffcff3fe7fff9ffffffffffff
R2[25] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbfee7fc7c666dc780380000000000010000009900007c1e998e0f7fffffffffffffffffff7fffffffffffffffff
R2[26] <= 640'hffffffffffffffffffffffffffe7fffffffffffffffffffffffffffffffffffffffffbf861383ce70984010800000000000000000080000000008c1c187dff3fffffffffffffde3fff7fffffffffffff
R2[27] <= 640'hffffffffffffffffffffffff1fc7ffffffffffffffffffffffffffffffffffffffffff003138383c400c008000000000000000000000000000000d0c1801ff7fffffffffffdece7fffffffffffffffff
R2[28] <= 640'hfffffffffffffffffffffffffc1ffffffffffffffffffffffffffffffffffffffffffe0030c00018000c0080000000000000000000000000000019c700c3fff3ffffffffffde71ef7ffeffffffffffff
R2[29] <= 640'hffffffffffffffffffffffeff01cfffffffffffffffffffffffffffffffffffffffffe0030c00081000000000000000000000000000000000000f1c703c3fbf1fffffffffcff73c73fffffffffffffff
R2[30] <= 640'hfffffffffffffffffffffe4d03001fffffffffffffffffffffffffffffffffffffffe60000000081000000080000000000000000000000000000d08401c771c7fffffffffe7f73ff3fdfffffffffffff
R2[31] <= 640'hfffffffffffffffffffffe48e101fcffffffffffff7fffffffffffffffffffffffff4600000000004000008000000000000000000000000000188808009e3187ffffffff3f31073ff79ddfffffffffff
R2[32] <= 640'hfffffffffffffffffe8e242040030223ffffedfefffee7fffffffffffffffffffff180800100000000000000000000000000000000000000810007628000f83ffffffeec96b9fcbff3c7f7ffffffffff
R2[33] <= 640'hfffffffffffffffefec4800000000c04ffffeffefffffffffffffffffffffffff300800000000000000000000000000000000000000000000000006080810ffcff00ffee9639fc1ffffeffffffffffff
R2[34] <= 640'hfffffffffffffffeffc0800000000c0cffffeffffcffdffffffffffffffffffff1800000000000000000400000000000000000000000000000000020008107e08e0fc306923880011c7cffffffffffff
R2[35] <= 640'hfffffffffffffffff3000100000080047ffffcfffcff9ffffffffffffffffff97c800000000000000000000000000000000000000000000000000000000800c084ffc106920100018e3f77ffffffffff
R2[36] <= 640'hffffffffffffff7ff3000100000000033fc0fcffe7e7fbfffffffffffffffef03c0000000000000000000000000000000000000000000000000000000018c0030000006010c100018707ffffffffffff
R2[37] <= 640'hffffffffffffffff710000000000000333c04d3fe7f773fffffffffffffffef8030000000000000000000000000000000000000000000000000000000000000321e018601043004283c0feffffffffff
R2[38] <= 640'hfffffffffffffff10000000000000000337c4f3fe7e066fffffffffffffffe8c010000000000000000000000000000000000000000000000000000000000000000ff00200000000003004effefffffff
R2[39] <= 640'hffffffff7ffffe730c0000000000010023fe4d3f38c066cffffffffffffe9f8c0000000000000000000000000000000000000000000000000000000000000000000001000020000001007effcfffffff
R2[40] <= 640'hfffffbfffcffe7ff000000000000000001000000c00c00fffeffffffffff38e00000000000000000000000000000000000000000000000000000000000006000000000800000000000713c1cfefbffff
R2[41] <= 640'hfffffffffffff39900000000000000000000000080c0001fcfffffffffff30000000000000000000000000000000000000000000000000000000000000000000000000000000000000301f3effffffff
R2[42] <= 640'hfffffffffffff8010000000000000000000000000101001fcfffffffffef80000000000000000000000000000000000000000000000000000000000000000000000000000000000000008307bf7f7fff
R2[43] <= 640'hffffffffff1f38000000000000000000000000000003000ffffffffffeff800000000000000000000000000000000000000000000000000000000000000000000000000000000000000083001f7fffff
R2[44] <= 640'hffffffffff0fc3c0000000000000000000000000000000077ffffffffcff800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fffffff
R2[45] <= 640'hfffffffffff8c300000000000000000001000000002000007ffffffffeff800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c101ffffff
R2[46] <= 640'hfffffffffcf8800000000000000000000000000000000007f3fffffffff7000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e021e7ffff
R2[47] <= 640'hfffffffff81e800000000000000000000000000000000007e3ffffffff070000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000071c3ffff
R2[48] <= 640'hffffffcff4000c000000000000000000000000000004000fc0ffffffe77c0000000000000018000000000000000000000000000000000000000000000000000100000000000000000100000001feffff
R2[49] <= 640'hffffffcce08004000000000000000000000000000000000f1fff7ffdfff00000000000000088000000000000000000000000000000000000000000000000000000000000000000000000000001ffffff
R2[50] <= 640'hfffffffc236001000000000000000000000000000000001f3fff7fffffc1000000000080008000000000000000000000000000000000000000000000000000000000000000000000000000030087ffff
R2[51] <= 640'hfffffefc212000000000000000000000000000000000010ffeffffff7ec000000003080000800000000000000000000000000000000000000000000000000000000000000000000000000001000fffff
R2[52] <= 640'hffe7feff6100100000000000000000000000000000000100ffffffff3c0000000000180001780000000000000000000000000000000000000000000000000001000000000000000000000000003fffff
R2[53] <= 640'hffe7fffff00018000000000000000000000000000000000007ffffe73c180000001801f003716066000000000000000000000000000000000000000000000000000000000000000000008000003fffff
R2[54] <= 640'hfffffff1e0000800000000000100608000000000000000000fffff6600000000000e037003677e66186000000100000000000000000000000000000000000000000000000000000000000000033fffff
R2[55] <= 640'hff7efff1ce808000000000000101608000000000000000001c7fffe70000000000010301f3e77f067c66c0000000000000180000000000000000000000000000000000000000000000000000c30fffff
R2[56] <= 640'hfffc9d7c03000400000000831101ff300000000000000090771ffcfc000000000000fce7ffff9ff9de00803100008000000000000000000000000000000000000000000000000000000000000c7fffff
R2[57] <= 640'hffffdffcf0000000000000008018733800000000000000013ffffcfc000000000018037fffffbfffdd00283b0000000000000000000000000000000000000000000000000000000000000000007fffff
R2[58] <= 640'hfee7fffef0000000000000100118730e00000000000000013fffffe000000000000003bfffffffffff3c7eff780000000000000000000000000000000000000000000000000000000000000000ffffff
R2[59] <= 640'hffcf66ff03800000000000201c00ff8e8000000000000000e3ffffe0000000000080f79ffffffffffffcfffefc0000000000000000000000000000000000000000000000000000000000000000ffffff
R2[60] <= 640'hff1c66ff0300800000000001fc00fff0f800000000000000e3fffee0000000000083fe9fffffffffffffffde800000000000000000000000000000000000000000000000000000000000000001ffffff
R2[61] <= 640'hff3c7ffff010800000000000c21cfefb10000000000000007fbf3ee000000000000c1fbfffffffffffffff9f800000000000000000000000000000000000000000000000000000000000000003ffffff
R2[62] <= 640'hfc38fbeff00000000000001c073ffe3f00400000000000007cff3ee000000000001f1fffffffffffffffffffc00000000000000000000000000000000000000000000000000000000000000001ffffff
R2[63] <= 640'h7cfeb9ef03000000000000cc62c77ffff966848000000000f3ff87e0000000000003ffffffffffffffffffffe08006000080c00000000000010000008000000000000000000000000000000001cfffff
R2[64] <= 640'hfffc83078c000000000078dc819efebff780e000000000013fffffff800000000439fffffffffffffeffffffdf0e0182000080000000000100000000000000000000000000000000000000008133ffff
R2[65] <= 640'hfffe01038c0000000004c39fc3feffffffffe000000000017bfffff0000000000719ffffffffffffffffffffde00011200000000000000000000000000000000000000000000000000000000000f3fff
R2[66] <= 640'hcfff00c000000000000007bffffffffffffff8100000000070ffff00000000007fdffffffffffffffffffffffef0801200080000000000000000000000000000000000000000000000000000008f03ff
R2[67] <= 640'hfff300e00000000000003efffffffffeffffd8000000000271ffff0000000000ffdffffffffffffffffffffffc18801200f00000000000000000000000000000000000000000000000000000000f03ff
R2[68] <= 640'h3ee780e0000000000000fffffffffffffffff9800000000203ffefc000000000ffdfffffffffffffffffffffec1000820220000000100000000000000000000000000000000000000000000000330f7f
R2[69] <= 640'h1ecf80c0000080000023c3fffffffffffffffd800000000003ffefc000000000ffffffffffffffffffffffffec700082030200000010000000800000000000000000000000000000000000000031bf7f
R2[70] <= 640'h8f8e8303000000000033e7fffffffffffffffe8000000000001f760000000020ffffffffffffffffffffffffff700080003f0000001000000780c3310000000000000000000000000000000000339fff
R2[71] <= 640'hc78c03070000000000333fffff7ffffffffffe8000000000000f7e000000011ffbfffffffffffffffffffeffff30009000fc3c00000000068f8cc33160000000000000000000000000000000008e07cf
R2[72] <= 640'h901807600000000000c7fffffffffffffffff9e08c000000003f9900000000c7fcfffffffffffffffffffff7e3898c01864e018000180000007000fee00000000000000000000000000000000083083f
R2[73] <= 640'h9998037400000000070ffeffffffffffffffffe083000000003f9900000031fffffffffffffffffffffffffffc980000007e800000001820e0c3fffe800000000000000000000000000000000003003f
R2[74] <= 640'hb98637e000000000c0fffffffffffffffffffdec00000000000800000007fffff7fffffffffffffffffffff7ef8000c087bc0000481fff1ff27ffff000000000000000000000000000000000033033f
R2[75] <= 640'hff1637e000000008063fffffffffffffffffefe300000000000c0000000ffffff7ffffffffffffffffffffff3fc00001e73c0000081c37fff3fffff000000000000000000000000000000000033833f
R2[76] <= 640'h7e726620000000003e7ffffffffffff7ffffefd38000000000000000000ffffffffffffffffffffffffffffffff800103f7c0002000c73fffffffffe00000000000000000000000000000000030033f
R2[77] <= 640'h26e62460000000001c67fffffffffffffffffff9c0000000000000000001ffffffffffffffffffffffffffff7fbf800103efc00031043e3fffe7fffff0000000000000000000000000000000003800ff
R2[78] <= 640'h600060000000001c7fffffffffffffffffffffcf000000000060000001ffffffffffffffffe11fffffffff7fff00030ffee00001047efffffffffffc000000000000000000000000000000008e00ff
R2[79] <= 640'h24006000000000067effffffffffffffffffce1e0000000000600000037fffffffffffffffe038fffffffff3fc110e3ffee2060406c3ffff7fffffff000000800000000000000000000000000600ff
R2[80] <= 640'h1000f080000000003fffffffffffffffffffffffde08000000000000001ffffffffffffffffc000ffffffffffff0063dffffc660e7f7f7ffffffffffc620000000000010000000000000000000003ff
R2[81] <= 640'hc00000000000000038ffffffffffffffffffffffff408000000000000001ffffffffffffffff8000ffffffffffff1839ffffff67317f7ffffffffffffee00000000000000000000000000000000003ff
R2[82] <= 640'h80000000011bffffffffffffffffffffffff020000000000000003ffffffffffffffff00000fffffffffef3c7fffffff99317f3fff7fffffffffd10000000000300000000000000000000030ff
R2[83] <= 640'h18000800000000007ffffffffffffffffffffffff010800000000000007fffffffffffffffe00000fffffffffffbff77fffffd81ef03ff03fffffffff9900000080003c0000000000000000000023bf
R2[84] <= 640'h18ffffffffdffffffffffeffffffd00640000000000007ffffffffffffffff00003fffffffffffe7ffffffffd98ec31fe03fffffffffd90000008007ff8000000000000000000003bf
R2[85] <= 640'h3ffffffffffffffffffffffffff9e680000000000007ffffffffffffffff00000fffffffffffe7ffffffffffcec78ef83ffffffffff90000000683fe8000000000000000000003bf
R2[86] <= 640'h13fffffffffffffffffeffffffffffe80000000000003ffffffffffffffff000001fffffffffffffffffffffffcfe8efc2fffffffffff783fc60ffffec8000000000000000000103f
R2[87] <= 640'h80000000000000ffffffff63fffffffffffffffffffee0000000000003fffffffffffffffe000007ffffffffffffffffffffff71fe8e7c3f7fffffffffff3fe7fcffdefcc00000000000000000383e
R2[88] <= 640'h2100000000000000ffffff630fffffffffffffffffffff98000000000007ffffffffffffffff000007ffffffffffffffffffffff9bc00e3003bfffffffffe7cffcf3fffefff80000000000000000703f
R2[89] <= 640'hfffffffffe7fffffffff7ffffffffffd000000000000fffffffffffffffff000018ffffffffffffffffffffffffff0ffe03fffeffffffe7df3ffbffffff9c0000000000000000003f
R2[90] <= 640'hffffffeffc067ffffffcffffffffffff100000000001ffffffffffffffffe00001c7ffffffffffffffffffffffffffffe00fffeffffffffffffffffffffff0700000000000000041f
R2[91] <= 640'h7fffffe000367ffffffcffffffffffff000000000001ffffffffffffffffe00000f7ffffffffffffffffffffffffffffe00bfffffffffffffffffffffffff0f60000000000000061f
R2[92] <= 640'h107fffffe000167fffffffffffffffffff80000000000ffffffffffff0ffffe000007ffffffffffffff3ffffffffffcfffe0cffff1effffffffffffffffffff7e46000000000000061e
R2[93] <= 640'h7fffefc000080fffffcfefffffffffffc0000000000fffffffffffffffffe0000049fffffffffffff8ffffffffffcfbfe8effff983ffffffffefffffffffffc47000000000000061e
R2[94] <= 640'h1ffffffc000090fffff9007ffffffffffc00000000023ffffffffffffffffe0000003fffffffffffff87fffffffffef3fb8effff080ffffffffeffffffffffff98000000000000003e
R2[95] <= 640'h1fffffc0000098ffff91017e7fffffff7f00000000027ff7fffffc7fffbeff0000003fffffffffffe31fffff3fe7ff717b87ff7f0c07ffff7ffffee7ffffffffb8000000000000019e
R2[96] <= 640'h3000000000018fffff8000000cffc038c11fffffffffd80000000000fffffffff3cff9ffff60000dfffffefff3e0008fffffffc7ccf77e84fffe420ffffffffffefeffffffbffc0900000000001807
R2[97] <= 640'h201fffff000000009e00000008fefffffffd0000000003ffffff8f70873fffff6000093ffffffc7100008fffffffff8ee166847fffe09ffffffffffffffffffffffd1100000000000900
R2[98] <= 640'h303fffff000000000000000000787ffffffc00000000037fffff9f00031fffff00000001ffc7fc2000000ffffffff78f03e3003ffff8efffffffffffffffffffffff0000000000000338
R2[99] <= 640'h303fffff0000000000000001003b7ffffffc0000000031ffffff1c0001dfffff000000036ffc6600000003fffffec00e07c3003ffff8e7ffffffffffffffffffffff0000000000008110
R2[100] <= 640'h8fffffe00000000000000000003fffffffe000000007bffeffe980000ffffff000000016ff02700000000ffffdfc03c01800067fff966ffffffffffffffffffffff6000000000000001
R2[101] <= 640'h3fffffe00000000000000000003fffffffe000000007ffffffcc000000fffe00100000065c100000000037ffffff838f0180087fef9efffffffffffffffffffffff6000000000000403
R2[102] <= 640'h3ffffffe000000000000000000008fffffff380000007ffffefc8000002fffc00000000060810000000002fffffffc00f098000ffffc8fffffffffffffffffffffff6200000000000600
R2[103] <= 640'hfffffffe000080000000000000001cfffffe7c800000ffffeffe180000663fc00000000060000000000000ffffff18031f88000efffc811fffffffffffffffffffff6600000000000000
R2[104] <= 640'h7ffffff60000000000000000001000fffffcffc00000fffffffc4000001f49200000000000000000000000ffffffc0310d80007fff8101fffffbffffbffbffffff7de30000000000000f
R2[105] <= 640'h7ffffff60000000000000000000000ffffffffc00003ffffff4800000007e90000000000000000000000001fffff80010dc0403fff98000ffffffc7ffffffffffffff10000000000000f
R2[106] <= 640'h3ffffff000008000000000000000017fffffffe000016fff7fc80400000f680000000000000000000000001fffff08c70d0041c3fff800007f9e8c1fffffffffffff7800000000000031
R2[107] <= 640'hbfffffb90000880000000000000003fffffffff000006fffffcc00000007090000000000000000000000001fffff1c8ec80101c17fe000c0331e000fffffffffffff7800000000000031
R2[108] <= 640'hfbffff9a000098000000004400000087fffffff8011f6fffde4800000007000000c00000000000000000001fffffdc1ce87001c03fe00001013000009fffffffff9ee180000000000031
R2[109] <= 640'hffffffba80007800000001ec0000001c7ffffffc0f83efffce6c00000000000000000000000000000000000fffffc03c4d60080e7fe00000012000001fffffffff9ec180000000000030
R2[110] <= 640'h80007ffffff680006000000001dc00800008e7fffffe87c0cdff8ecc000000000000000000000000000000000407ffff84214d03088e7fe00000000000007fffffffff9f2000000000000000
R2[111] <= 640'h38007ffffff60000600000000d9903800003c0fffffec37ec9ffc7c0000000000000000000010000001811888407ffff0e417cc000c83fe0000100080000ffffffffc68b3010000000000000
R2[112] <= 640'h8660007ffffffc80001880000c1fd9f6640002019ffffcce67ffffdf7c00000000000000000000c000000040003003fffff33bdc0081301fc00000000080003ffffff80f1c0c30000000000003
R2[113] <= 640'h10400fffffffc8000008000049ffffffe0000011ffffedf67ffffff60000000000000000002400000000009f00003ffffff309f0800013fd1000000000000fffffff00020c120000000000003
R2[114] <= 640'h310400ffffffff000003810000fffffffe0000003fffe787cfcfffe74000000000000000000340000000047db20007ffffffe0f10800803f80000000000000cffffec000614100000000000001
R2[115] <= 640'h310000fffdffff0000070000013fffffff030000ffffe7efd97ffffec00000000000100000024000000004ff903007fffffcf0f0c800003f800000000000001fff7e0000003000000000000000
R2[116] <= 640'hf70007ffffff80000073000017fffffff90c001fffffffff97bfffc48000000000c1800000080001c0001fd907003ffffffff1ec800003ff40000016000003fff26000000080000000000000c
R2[117] <= 640'h8ff1007ffffffc00000080000087fffffff3e001fffffffff97bff3c08000000000c98000000c8000e0003ff90f000ffffffc7de4800000fe00000006000007ffe200000048000000000000004
R2[118] <= 640'h10000fff100ffffffff00000080000007fffffff34000fffffffffcfffffc00000000000ef8000003fc88006007ff838000ff1ffe84e40900000fe60000180000003ff8000000000000000000000000
R2[119] <= 640'h3fff900ffffffe1c000de0c00000efffffff20000ffffff7fdecfffe000000000007ffc000003fd8004608e7fc08000001fffc46748000c0ffffc12010000007ff1800000003000000000000021
R2[120] <= 640'h1dffd807ffffffc80003e0ff10e07ffc9ffe00000ffffffffffffffc700000000007e3f880001ff300e9c67ffc00002227fffcf7f4000011fffffcfc63800013ff0000000000000000000000300
R2[121] <= 640'h10001ffff80ffffffe30000070f3d0007ff0038f800001fffffffffffffe000000000003f7f80001fff601e9e7f7fc0000200ffffef7f4000018fffffffefe00001ffe0000000000000000000000000
R2[122] <= 640'h3ffff84fffffff30000031efc9e07fe0000280003ffffffffffffffe0000000000007ffc0003fffe00f9f7fffc0000000ffffffffc00001c7fffffffff0003fffe0000000000000000000000000
R2[123] <= 640'h1fffff80ffffffff000018c0ffff0ffe0000000007ffffffffffffff7000000000001ffff1817fffc00fbf7fffc00000023fbffffecc00001ffffffffff8c17fff80000000000000000000000000
R2[124] <= 640'h1103fcfffff8fffffffe000019c07ff0ef8f400014c31fffffffffffffff700000000007ffffff99ffffc00fffffffc00000003f9ffffffe20003ffffffffffe00ffff00000000000000000000000004
R2[125] <= 640'h107c7fffff87fffffff080001e37fff07efcfce00037fff3f9ffffffffff00000003247fffffe3fffffc0ffffff7ec00000003817fffffe6090e7ff7c7fffffffffff00000000000000000000000000
R2[126] <= 640'h800f8fffffff3ffffff7180001e17cff07feffff00007fff7fbffffffffff800013833eefffffef9ffffe0fffffffee00000000003ffffcc6081ffc1203ffffffffffe80000000000000000000000000
R2[127] <= 640'hefffcfffffffffffffb000000000701837fff7f200083fffffbffff7fffec00010113effffffff97fffe3cfffffc7e00000000002ffffcc20013c80002efffffffff680000000000020000000004001
R2[128] <= 640'he799fffffffe7fffffcec0200000096e63bffffff000013fffffffffffffc000061c3effffffff9e7efffffeffff630600000000007ffeee7c9804000062efffffffe480000000000381000000000000
R2[129] <= 640'h1efffffffffefdfffef01800000009fec7ffffffff800047ffffffffffffc000060fb77fffffffdfffffe79f3fff703e00000000007ffffe6c81e0000022fefffffffc00000000000081000000000000
R2[130] <= 640'hffff9ffffffffdfbfcf0188000000fffffffffffff800007ffffffffffffd000001f837fffffffffffffe7fe37ffd07e80000000003bffffedc100080022fe9fffff1c00000000030000000000000000
R2[131] <= 640'hfffffffffffffffbffc0018000000ffffffffffffe00003fffffffffffffc00000ff16fffffffff3ffffc6f83fffc1ff00000080001bffffeffb000400226fbfffff800000001007003c000000000000
R2[132] <= 640'hfffffffffffffffc8180018000006fbfffffdfff9e00007fffffffffffffc00c1fffffffffffffe3fffffe31b7ff81ff000001c00000e2fffffddc80382226bffff8c00000001900016e000000000000
R2[133] <= 640'hfffffffffffffffc0080000004007fffffff8ffe1e00c1fffffffffffffbc00cfffffffffffffee0fffffe71bb7e3bff800003c08000003ffffddec138ff70bffff8c0000000001880c6210000000000
R2[134] <= 640'hfffffffffffffffe00000c0000001fffffff86fe8200fb1ffffffffffffb0047fffffffffffffee018ff7ef012647fff80001f268080001bffff9ff3fbff709bff9b00000000c43ff0cfe10000000000
R2[135] <= 640'hfffffffffffffff600008e0000000fffff7ffeff83830039ffffffffffff00c7fffffffffffffee0001f20c010fc7ff70001ff3f078000017ffff3f9f7ff2089fe800000000106ef3c9cc40000000000
R2[136] <= 640'hffffffffffffff7010000100000007ffffff7efec7c0011fffffee3fff9c001ffffffffffffffec0040f626018197fff0001ff0f19c740001ffffbffffffc03f676e80000061017ec6f3c08200000000
R2[137] <= 640'hfffffff33f7ffff080000000000007bfffffe7fe86c00003ffffee9fff98000ffffffffefffff6c00600f2400000fff10007fffb0fffe0401ffffffffffec0fc62e01800000dc3efe7f3070200000000
R2[138] <= 640'hffffdff21fffffd8800000010000011fffffef7e0e4800027fff020ff8908007ffffff3c7ffff7000000b6400001fff00007fff30fffdc601cffffffffff80e000060000000cfffffffeff3600000000
R2[139] <= 640'hfffeffbe3fffff988000000000000118fffffffe1ec0000073ff011878000103fffefc803fffff00000316c00003ffe00007fff307ffdb001c3fffffff3f00c1091c000000c4fffffffefcb600000000
R2[140] <= 640'hffffffb0073fff184000800000000199ffffffbeffc0000001ff113878040107ffffe0803ffefe00000016c00000ff000003ffc737fff100800ffffffffc0003093800000001fffffffffca600000000
R2[141] <= 640'hffff7b80033ffcc3c00000000000000fffffff96ff78000001ff01d16380081fffff01003ffe900000801ec0000739000003ff8e39fff000003feffffffd000300c020000038ffffdfffffa640000000
R2[142] <= 640'hffff668001fffce6c60000000000000fffffffb23ff800400070608c0300001ffff901003bfd8000000012c0000710000003ffc43bff600000ffffffffbf3c00c48300000178ffffffffffb660000000
R2[143] <= 640'hfffde61000fffeeeee60300000000003ffffff7303f8600000f8601c3c00001ffff931013bd9b000000000c00040f920000ffff09fff80040d1f7ffffff87c3046980000810ffffffffffffe60000000
R2[144] <= 640'hfffff6c0017fff3e7ed8400000000001fffffe9866ffc100007fe88c388100fff7fe910311fc00000000000000007e80006f38e43fff00036167ffffffffe6fc60008e00624f3cffffffffe3c3000000
R2[145] <= 640'hffffffdc016fff7ff7f90200000000001ffffe9b7e7fc90000ffc9c0e300003ffffcf000116000000000000000063f000001b2e037f80103767fffffffff07ce20001c00647efcffffffffff70800000
R2[146] <= 640'hfffffffc81fffffffffd07000000000007fffff3ffffec80037f49804380000ffff874000000000000000000000400000000e08003c003fffefffffffffff6cf000088003c7edffffffffffff8800000
R2[147] <= 640'hddffffff99fffffffffd0c100000000000fffff7dfffec80017f400100c8000ffffd268000400040000000000000800000000000038601fffefffffffffffcdf8600800108ff8fffffffffffc0000000
R2[148] <= 640'hffffffffdfffffffffffcef80000000003fffe7fffffec0000ffe83000c00007ffff00000000000000000000000000000000000001c000ffffffffffffffffff8e00000001fffffffffffffff0000000
R2[149] <= 640'hffffffffffffffffffff9effe000000003ffbf7fffffec00007f49f001c200e7feff00000000000c3e0100000000000000000000007c007fffffffffffffffff86001c0001bfffffffffffff3c000000
R2[150] <= 640'hd97fffffffffffffffffbfffe000000000ef33fbafffc800037fe8c003e400febef30100000000003ffb60000000000000000000003e00ffffffffffffffffff8000180009fffffffffffffffcc00000
R2[151] <= 640'hd17bfffffffffffffffffffff0000000038e33837fffc800007fe80018e00000b3f7998100000007fff9e0000000010000000000000000f1ffffffffffffffff0000c100187bfffeffff67ffe3600000
R2[152] <= 640'hc399fffffffffffffffffffff800100000121e80fefc3000003fb93806c080017e7c9002808000007fff7c66000000000000000000000c3efffffffffffffffefc1ce0000fffff99c78f3fffff600000
R2[153] <= 640'h9bfffffffffffffffffffffc80000000801ee0fec10000001f993843f800003fc70002060000007ffff700000000000000000000000fffffffffffffffffffc09ec0000fffff98ff9f0fffffd00000
R2[154] <= 640'h20bb7ffffffffffffffffffffc0090000080c6003fc00000709ff93c63fe480000840001030000007fffffc00000000000000000000007ff3fffffffffffffffe7fec000effffffeffbf8fffffcc0000
R2[155] <= 640'he0773ffffffffffffffffffff901f3000010e2023b00000178defd0c73cf640000000001000640007f7f7f800000000000000000001803ff07ffffffffffffffffcec0003bffffeefffb9bffffdc0000
R2[156] <= 640'he3277ffffffffffdffffffffffc0f3c0001000800000000079fe388f7fcf67400000000000020000736ffc000000000000000000028c01fffffffffffffffffffffe070c3bfffffefff39ffffff00000
R2[157] <= 640'he020c7fffffffffd7ffffff7ffc0f3c0008000004000000033ff3c8ff7fe7d7e000000000002000003fdf900000060000000000000c000fffff01ffffffffffffefe01003ffffffe7ff31ffffff00000
R2[158] <= 640'h37efefffffc017fffffff81f2e00080000fc0000000637ffffeff7fff7f660000000000000007ffd8000070700000006000000381fffff01ffffffffffffffe0000ffffffff3ff31ffffffc0000
R2[159] <= 640'h400f0bc6fffffffc01ffffffffe1f6e00010001fc4000000e17efffeffe7ff7fe0000000000080000f4fdc4023787380000dc6000179837fff76007f7ffffffffffce003cfffffdb7ffb07fffffe0000
R2[160] <= 640'he10738897f7ffffc01fffffffff0df780000001801000000c7e8d9fbf867fffbd9c00000000001039f3e7200f7fff900000f8000433fc1ffdf800000181fffffff7ee639ff7ffff3fffebfffffe40100
R2[161] <= 640'h3807b31d3cfffffc00bfffffff98df780000000000000000004f1fff996fffffc9c00000000000f09f8f7001fffff9c0c006000040fcc0fffc0000000001ffffffff6ee3ffffffffffe4bfffffee0000
R2[162] <= 640'h3807937d6cfffffc00bfffffffb8f3f80000008080000000006d7fffc16dffffcbce0100000000f0fecffc003ffffc80800400000c3e41fff80000000000ffffffff7ee3fffffffffff69ffffffe0000
R2[163] <= 640'h40834fc67ffffe00fffffffff0f3f8000000000000000007e87fffc0e1ffffffff00000000017fffeffe8016fffc000c00c000010f017ef18000000000ffffffffff3ffffffffffeff8fffffff0000
R2[164] <= 640'h8170024f8e7fffff00bfffffffb3fff8000000000000000006492fff00e1feeffffe0080008003fb67fffe80008ffc101800000001c0087fe70000000000ffffffffff3cffffffffffff9fffffff0000
R2[165] <= 640'h83e026f1c66ffffc01bffffffbefef9000000000000000000417ff3041ddffffffc8380008003ff677ffe080003fcf020000000008000831c00000000007fffffff38efffffffffffd93fffffff0000
R2[166] <= 640'h1804226d20667fddc001fbfffffffff900000000000000000040fff7063dc7ff7fffc3000000007ffbfbfff800000000000000000000000110000000000003ffffffffffffffffffffd97f7fffff0000
R2[167] <= 640'h880002e1e32f7ffc00037ffffffffff9000000000000000000019fe6e0c933ff7ffff820000007fffbf9ffe100000000000000000000000000000044000003bffffffffffffffffffff9e3fffffe0000
R2[168] <= 640'h4100003e38998ffc001d7fffffffffffc0000000000000000001ffe748c007fffe77c18330401bfebfffff7f0100000000000000000000000000980000001cf3ffffffffffffffffffeffffffffc0000
R2[169] <= 640'h6c0000392001e3f36001fffffffffffec00000010000000000003ffecf807cffff3c489070051ffefffffffe6018000000000000000000000000088000000cf3fffffffffffffffffffffffffffc0000
R2[170] <= 640'h180000318007312100016fffffffffffc1010000000000000006fffecf800efffb7ec89800681ffffffffffefc7800180000000101001f0000008080400001fffffffffffffffffffffffffffffe0000
R2[171] <= 640'h88b000118006210000003fffffffffffc0000000000000000007f3e7edf807fefcf7811f00689cbffffffefffe1f6d8000000001f118fffc000000000000011fffffffffffffffffffffffffffff0000
R2[172] <= 640'h81b0009c0000000000003cbfffffffffd0248000000000000003ffe7fdf8dfffcee28118900d1fbffffffeffff8f7fe190000002fc11ffff000000040000000fffffffffffffffffffffffffffff0000
R2[173] <= 640'hd000c9c00000080000003fffffffffff8c680000f00000000037f3c78c01fffdf3c00011e0707bffffffffffecfffffba00000efc17ffff4000200e800000007ffffffffffffffffffffffffffe0000
R2[174] <= 640'h4c0208df00000000000001fffffffffffc63800019800000000fff7e79c01ffffc3e00070744c6fffffffffffcfffffffa000006ffff7fffc000c000000000003ffffffffffffffffffffffffffe8000
R2[175] <= 640'h608600c3800000000000001ffffffffff020081cf0800000000effff7fc69ffcf0024000934c06f7fffffffe3c3dfffffe000007ffff7fffe2388000000000003fffff9bffffffffffffffffffcf8000
R2[176] <= 640'h2841888c100000000000067fffffffff900000cc0000000000ffffe3f7d3fe4600400004d7cdffffffefffc98c3ffffff70000ef77efffc78000000008000003edeb946fffffffffffffffffffbf800
R2[177] <= 640'h408603899800000000000067fffffffff80000071f3000000007fffefb690fe4400200004dff9ffffffffffe9873ffffff60000ff7ffffc00080000000800000273f00007ffffffffffffffffff93800
R2[178] <= 640'hc087c7191c00000000000003fffffffffc0000013cf000000007fffff14186e0000000000fffffffffff7ffe801ffffffc000007f7ffffc00000000000000000033100003fffffffffffffffffff0000
R2[179] <= 640'h477fff39dd00000000000018ffffffffff000000fcf70000001ffffff340cf70000000181f7ffffffffffffe0007ffffff00000033fffc000000000000000000000000001f7fffffffffffffffff8040
R2[180] <= 640'h2e7fff70df00000000000000fbfffffeff0000008fff1001003ffff8ffccf370000000091ffffffffffffffc06e1fffffb00000033fff800000000000000000000000000067ffffffffffffffff8c000
R2[181] <= 640'h7c7fc7701c0000000000000007fffffeff0000011ffe80000003ffffffcc7170000000006dfffffffffffffc1c18bffef0000000031cf080000000000000000000000000007ffffffffffffffffc7c00
R2[182] <= 640'h26ffffe61c000000000000000f7ffffffe8000003ffe80000003ff9fff4800000000008049ffffffffff3fff8007bffe2000000002093000000000000000000000000000001bffffffffffffffff3c00
R2[183] <= 640'h7c7fcc6c700000000000000183ffffffc8000007fbf81000010fdfffe610000800004010fffffffffffffff80e1bfc700000000008100000000000000000000000000e0001bfffffffffffffff7c100
R2[184] <= 640'h19feff7bb900000080000000007fffffff1800016ffff000000177f99f843000000000300dfffffffffd768c80009f9800000000000000000000000000000000000067600018ffffffffffffffdf6400
R2[185] <= 640'hffffffe3ff00000000000000002ffcfff60000007fffffc000017fffb90000000000000083fffffffffd674c80000fc0000000000000000000000000000000000000fffc0000ffffffffffffffdd4000
R2[186] <= 640'hfffffff3ff000000000000000003f8ffff000000ffffff800000feff300000000000000003fffffffffdc70181101180000000000000000000000000000000000cff7fff18001fffffffffffffd8c000
R2[187] <= 640'hffffff7eff0000000000000000193fffff060003ffffffc00004fee6000000000000000000ffffffffffd80101003901000000000000000000000000000000001effffffc0000ffffffffffffff8c000
R2[188] <= 640'hffffffffffe000000000000000193ffffc060003fffffff8004c1fee0000000000000000003fffffff6d1c0180003000000000000000000000000000000000001effffffe30007fffffffffffffc6000
R2[189] <= 640'hffffffffffe0000000000000000067fffcc20003fffffff0800f9fec0000000000000000013ffffff949000080000000000000000000000000000000000000080ce7ffffff8007fffffffffffff40000
R2[190] <= 640'hffffffffffe0036030000000000067ffffe30407fffffffb900df9f8000000000000000000fffffff948400000000001000000000000000000000000000000000083cffffc8007fffffffffffde40000
R2[191] <= 640'hfefffffffffc4060b000000000046effff3c4c67fffffff19108db310000000000000000003ffffff140020000000080000000010000038000000000000000000083fffffc0006ffffffffffffc00000
R2[192] <= 640'hfffffffffffc39b39000000000003f73ffffe13fffffffff7c193ff80000000000000000008ffffff8c80020080200008000180000600000801800000000000000006ffffec00ffffffffffffff11800
R2[193] <= 640'hfffffffffffff9301800000000003b73ffffffffffffffffe67fe700000000000000000000007ffffe08000000000000000080000801800000013000000000000001ffff9c0000ffffffffffffe10000
R2[194] <= 640'hfffffffffffffdbe18000000000078e7ffffffffffffffffe7ffe700000000000000000000017f7fe6000000000000000031e0000e0b7100000018000000000000006ffe180003ffffffffffffe00000
R2[195] <= 640'hfffffffffffffffff800000000001fffffffffffffffffffffe6fe30100000000000000000006ffde600000000000000003fe00007dd3180000001000000000000004df80000077fffffffffff380000
R2[196] <= 640'hfffffffffffffff7e000000018000ffffffffffffffffefffffffe80000000000000000000004dc660000000000000000c3f700000dd8700403083000000000000000d70000001fffffffffffcf80000
R2[197] <= 640'hfffffffffffffffff000000000800c3fffffffffffffffffffffef88000000000000000000001cc62000000000000000033ffe0000cdce980021000e0400000000000000000003fffffffffffcc00000
R2[198] <= 640'hffff9ff803ffffffff00000081800c3fffffffffffffffffffffff00000000000000000000000c040002800002400000837fff800067fffc0000000c0000000000000000000007ffffffffffffc00000
R2[199] <= 640'hfdfe1ffc03f3ffffff00000001810f037ffffffffffffffffffffe901001010000000000000000200000f3389e4000001dffff98007c3ffe00040c1c03800000000000000000019fffffffffffdc0000
R2[200] <= 640'hfc3c01e0003fffefff3001000660043fffffffffffffffffffffffe00110000000000000002000000003ffff7fe00003cfffffe6001f9f7f103166890000000000000000000041fffffffffffbf80000
R2[201] <= 640'hf8000060003fffefffe0c00006e6e07fffffffffffffffffffffffd88100000000000000000000000007ffffffe80007ffffffff00199fff303f068880000000000000000000497ffffffffffff10000
R2[202] <= 640'hc0000000000e7f00ffe30000c7fff8ffffffffffffffffffffffff9c88860000000008000000c000003ffffffffc000ffffffffec0001e7fc0fb604080000000000000000000090ffffffffffe910000
R2[203] <= 640'h4100fff30f00ff9f78ffffffffffffffff7ffffffffe000000000000000000064000007ffffffffe003fffffffffe0003666c4f0e4640000000000000000000349fffffffffffe010000
R2[204] <= 640'h40003ff9f80cffff7fffffffffff3fffffffffffffff0010000000000000070e04040fffffffffff81ffffffffffe000020080060f400000000000000000000048ffffffffff3fe00000
R2[205] <= 640'h7ff9f03fffffffffffffff7f7fffffffffffffff312300008000180e37ff8006ffffffffffffc1ffffffffffe000004000ccc000000000000000000000034dbfffffffff3fe00080
R2[206] <= 640'h20000000000007fffffffffffffffffffff7fffffffc17ffffffff903000000001c8fffffd90fffffffffffffffffffffff7ff800000000c0c00000000000000000000007491fffffffff9fe00080
R2[207] <= 640'h38020000000003bfffffffffffffffffffef1ffff7f387ffffffff80000000001c78fffffff9bffffcfffffff7ffffffff7fffc0000000000000000000000000000000000c9fbffffffff9ff66000
R2[208] <= 640'h6800f200000003bffffffffffffffffffe798ffffff30cffffffce010000000008fdfbfffe7fffff9ff00ffffffffff7e00ffff0000000000060000000000000000000004c1c0fefffeff97ffc300
R2[209] <= 640'hfc31c000001bffffffffffffffff7f7fdffeff7ef08ffffffff680000000006ffffffffffffff0000080ffffff0100003fff000000000000000000000000000000000018007fffffff87fffc00
R2[210] <= 640'h1bfeffe0000003fffffffffffffffffffd9fffff78000ffffffff0800000001077fffffffffffe0020000007ffff00000019ffce000000000000000000000000000000000c007fffffff87fffc00
R2[211] <= 640'h1efffff7020003ffffffffff77ff7efff9fffffce000077f7fff80000000003b7fffeffffffffc0400000003fffe00000001ffff000000000000000000000000000000000101fffffff98fffffc0
R2[212] <= 640'h11effffffffc00187ffffffff2480f8fffffffe7dc00000ff7fff00000000007ffffffffffffffc000000000010fc000000001ffee00000010003e23be30000000000000001007efffffd1fffe7e0
R2[213] <= 640'h187ffffffffe00087fffffffc100178fffffffeff000000fefffe000000000027ffffffffffffc0000000000001000000000007ffe08000096007ffffffc100000000000000000e3f7fff03fffff8
R2[214] <= 640'h3fffffffff000007f7fe000000000fffffffff000000000ffcc00000000f07fffffffffffffc0000000000000000000000000fff1000199fc3ffffffffb0000000000000000007e7ffea1ffffff
R2[215] <= 640'h33fffffffffb80003c18c0000000000ffffffec00000000018c0000000007c7fffffffff9f73800000000000000000000000001ffff739dffefffffffffef88000000000000000c3f3fe29ffffff
R2[216] <= 640'h1fffe7fffffe80000000600000000013fffffe0000000000000000000000cfffffffffffef000000000000000000000c0000000fffffffffffffffffffffe608c0000000000004202477a6ffffaf
R2[217] <= 640'h7ffe33f7fff0000000000000000000fffffcc0000000000000000000020fffffffffffff8000000000000000000001f0000000dfffffffffffffffffffffeff010000000000000000e9deffffe7
R2[218] <= 640'h3e003ffee3f83ffff0000000000000000007fffd000000000000000000000070fffffffffffc38000000000000000000001ff80000017fffffffffffffff7fffffff870000000000000000f80c7fff65
R2[219] <= 640'h3f807ffc00e007fffc000000000000000003ff7800000f0e000000000000001fffffffffffff30000000000000000000000ff800000007ffffffffffffff3cfffffffbc0000000000000005e2dfffff7
R2[220] <= 640'hfff9ffff000303ffff800000000020000003bf480000039ff80000000000003fffffffffffff710000000000000200000003fc80000003fffffffffcfbffc01ffffffc80000000000000005f9dffffb3
R2[221] <= 640'hfffffff7000103ffffe00000000738000003fec1000023fdf8000000000000fffffffffffffbe00000000000000600000007fc000000013fffffdbf8ff87801efffffe18c00000040000003f093fff93
R2[222] <= 640'hfffffff7000001ffffff9001000fff800003b000000077fbfc0c0006710083fffffffffffff8e0000000000000e78004000fff000000000f07ff99707801001effffff9ccc3c00040000001d3db9ffd9
R2[223] <= 640'hfffbf3f0000000fffffff801f88e8ec00000330000063fffc69c03effb81fffffffffffffffc00000000000001e7c08e0107ff00c000000000ff980010000083ffffffc7ffe7080000000004cfbfffc9
R2[224] <= 640'hfffff4000000033cffffff77ff079e00000000000003fffffffffffffff9fffffffffffffff01000000000000f03200f3e3ffffc8000000000010000000000007ffffffbffffb046c300002bdb95ffeb
R2[225] <= 640'hffffe00000000100ffffffffffffde00000000000001fffffffffffffffbfffffffffffffffc80000000000005c0009fbffffffc0000000000000000000000003fffffffffffb08687e00027e9c86de3
R2[226] <= 640'hfffc000000000000f0ffffffffffff0000000000001ffffffffffffffffffffffffff3ffff3800000000000002c03bfffffffffe0000000000000000000000001fffffffffffb4b4f70001b3edb8ef62
R2[227] <= 640'hffe0000000000000001fffffffffff8000000001003fffffffffffffffffffffffffe77cfc1800000000000000a03ffffffffffe7000000000000000000000000fffffffffffffea221a2163ffdc1973
R2[228] <= 640'hffc0000000000000001fffffffffffe00000000f03ffffffffffffffffffffffffffff3c8000000000000000201ff8dfffffffff78000000000000000000000007ffffffffffef67081aeb6f4ed75052
R2[229] <= 640'he7c0000000000000001fffffffffffe00000001fffffffffffffffffffffffffffff3e000000000000000000780ff0fffffffffef8000000000000000000000003fffffffffffef8354feb7c5253b456
R2[230] <= 640'hc1c000000000000000007ffffffffff80000003ffffffffffffffffffffffffffeff00000000000000008000f8077bfffffffffee0000000000000000000000000fffffffffffe7eafcfea57dc761592
R2[231] <= 640'h1ffffffffff80000003ffffffffffffffffffffffffffeb98000000000000000800cf8833ffffffffffce00000000000000000000000000ffffffffffe4b41cffa9875bf590b
R2[232] <= 640'h8000000000000000000ffffffffffc6000077fffffffffffffffffffffffffcffc000000000000000cfc001967ffffffffffffe000000000000000000000000001fffffffffe6c350ff12ccf9a98d7
R2[233] <= 640'h7fffffffffff8001fffffffffffffffffffffffffffdffc0000000000000003fc00197fffffffffffffe000000000000000000000f0000003ffffffff5b0b87e75a13646887
R2[234] <= 640'hfffffffffffe823ffffffeffffffffffffffffe7fffefe0000000000000103f800017effffffffffffe000000000000000000000fc000000c35fffff38afdfe17d5a6ca3b3
R2[235] <= 640'h1ffffffffffff37ffffffefff3ff7fffffffffc3ff10000000000000000101fc00013effffffffffffe0000000000000017880c3fe080000011fff7db6670fe54ae4852b67
R2[236] <= 640'h7feffffffffe3fffffffcf800033fffc0ffff03ff00000000000000000000fec01e3e7ffffffffffff0000000000000013ce0fbfc38000000071d66b24d7ff547f5d8960d
R2[237] <= 640'h6fcfffffffff7fffffffff800001ce0003fff000000000000000000000000fee03e363fffffffffffe0000000000000001f9cfffffc000000009b669719ddf4d5c535df40
R2[238] <= 640'h6981ffffffffffffffffffe00000000000fe10000000000000000000000001c0066061ffffffffffee00000000000003083fffffbfe0000000003ae910acf77e80ffe0e4e
R2[239] <= 640'h707dffffffffffffff7ff00000000003fe0000000000000000000008081000067071fffffff7fffe00000000000003881fffffdff00000000137e4e94bbc5dcae370d79
R2[240] <= 640'hc03fffffffffffffffff000000000007f000000000000000000000000008fc1820083fffffffffef00000000000000100fffffc5ae00000001b1fd3b66da00af3e3dc9e
R2[241] <= 640'hfff7ffffffffffe1e000000000027f00000000000000000000000001ce9e8c0003ffffffffff20000000000000020ffffffcdbe000000038130d5ef9c0e44df6d224
R2[242] <= 640'h503ffffffffffc04000000000003c00000000000000000000000001801c2c0001ffffffffffe8000000000000061ffffffff9b24100001850b40be3d48b52a889c1
R2[243] <= 640'h1ffffffffffc0600000000000000000000000000000000000000900100e2000ffffffffff18000000000000063ffffffff9b34180020b88fe5f098bdad34772c8
R2[244] <= 640'h3f7ffffc7bc0000000000000000000000000000000000000009c00e007a0000fffefffff78000000000000061ffffffff9b3da60021ffeb6077e4c38751f560b
R2[245] <= 640'h1e73fe8039c0000000000000000000000000000000000000008c03f103e00003ffffffff3800001e000000013fffffffff93de60008f0593b39e89f4240bc2a0
R2[246] <= 640'hc0100000080000000000000000000000000000000000000079c03f303e000003fffff0e7c00000000007803fffffffffe93d4a020ca1d86b96f266eae1f5875
R2[247] <= 640'h40000000c800000000000000000000000000000900000000788017f1ce000003ffffe003c00000003007803fffffffffe93d0b522f0b6af74f512d6f7aa6ded
R2[248] <= 640'h2100ff880000007ffffc800f000000003f00073cffffffd45343b9608a41ace2a333d89af928c4
R2[249] <= 640'h8040000000000000ff80000000ffffff0e0f8000000f3f000f81ffff7fee9b67b121deab14bb40a3664d509b7a
R2[250] <= 640'hc00000000000000000000000000000000000000000000000000000000000000000000429e00000000000007ffc000000ffffffbc0fc000003fc2000fc3ffffff49f281882086b6a500c4c3c40212b7b0
R2[251] <= 640'hf00000000000000000000000000000000000000000000000000000010000000080000c3de000e000388001bffe001c01fffffffce0c000001fe2020fe7fffffecc7df7dfe0acd8d3778fa17f8353cf1e
R2[252] <= 640'hf000000000000000000000000000000000000000000000000000000380000000bf00133c403ffc20fefcc1ffff007f83fffffffce0c000010c0003ffffffffbee5de402f6926c918ea8aa13edaa5c3d6
R2[253] <= 640'h3380000003ffc3ffbdeffffc71feffe1ffcf003ecffffffffff8c00381c0000fffffffffbea1babd67a15543bbf87ed0078f9de4d7
R2[254] <= 640'hfe00000000000000000000000007300000003bfe3fff9fffffffbf87ff1ffeffffffffffffffffdfe0b238000bffffffffffe8a964cf261b6f0bfa532cd2b37c98658
R2[255] <= 640'h1000000000000000000000001fef000000000000000000000000071200000023fe3fff3ffffeff3e2fff807fffffffffffffffffffff803c003fffffffffff6e1de7a3b08dc969e4534d41e5b8896d2
R2[256] <= 640'h80000000000000000000000000fee8000000000000000000800000793000000e3fffffffffffffffff7f63fffffefffffffffffff7ffc401c003fffffffffffb1e45592c68f898dede66e2167d1b1145
R2[257] <= 640'h7c000000000000000000000001fefc4000000000000000000000017bf800001f1fffffffffffffffffffc3fffffffffffffffffffffff001ffffffffffffffbad76adc8a66ee9d93708d9196aac34bb8
R2[258] <= 640'h3c000000000000000000000607fffdffc00000000000000000000331f800001fcffbfffffffffffffffe8ffffffffffffffffffffffff1fffffffffffffcdf34839f5e92493bf1b035f4bd419fcd12c7
R2[259] <= 640'h800000000000000000080071fffffffe0000000000001800000037bf800fe3fffffffffffffffffffff1efffffffffffffffffffffff9afffffffffffffcfadc65a7f389e9b4c347aa87286ee86c6ef
R2[260] <= 640'hfc0fe3f03ff3ffffc000000000003c0000000ffe000b8ff7ffefffffffffffffffffffffffffffffffffffffffffaafffffffffffffffb6e3b3f6aaf9ce17fd6fe875c3e5d8a8cd
R2[261] <= 640'hfc1ffff03ff3fffff000000000003e0c00000ffc000e2ff7fffffffffffffffffffeffffffffffffffffffffffffffffbffffffffffffdb2d2f53cccd2ac1007a07975ea8921a2a
R2[262] <= 640'he1ffffe3ffffffff000000020003c0c00000ff8f009bff7ffffffffffffffffffffffffffffffffffffffffffffffff7fffffffffffea5a8e3792b4f71a9b1d2a99efb62f9a865
R2[263] <= 640'h8ffffe3fffffffe18000003801fc17800007fe7e8fe3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaa91ad6275fdba2925a1f9de2b3b849aa0
R2[264] <= 640'hfffffffffffffff80000001000382000001efe0fce0ffffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffff5d0a83aef94da6127e542a2db6374c2976b
R2[265] <= 640'h1ffffeffffffffffc0000000000200800001efc07ebfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffed57bb6efcf847ee98b3e7a2e2da07eb1de3
R2[266] <= 640'hfc0000000ff00a7fffbffffff800000100000180000087807ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff6cbc8398c78fbcc5466daefabd736f55eea
R2[267] <= 640'h3e800000000006fffffffffffa00000000c031c000000f003e3fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbb6178cd83f1dee6239fe302935efe4d6677
R2[268] <= 640'hc0000000fff000000000018ffffffffffffec3000000c03be0000000001e3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff72db7ee8f5f76b3d67768e1892b7851cb2a
R2[269] <= 640'hc0000000ffe0000000000fffffffffffffffffff0000fe7fe0000000003ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff320bffe353b02c378edf66bbae4ece7ff73
R2[270] <= 640'h3fce01f00003fffffffffffffffffffff8000dfffe00000081cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb05bfbb2e7980ce13d9ad522ae5475040fcb
R2[271] <= 640'h780003f00003fffffffff7fffffffffff80000fffc00000083efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9cef75df9ef6fefb1d8dd69135a5b47d161
R2[272] <= 640'h30000138000007ffff3ffffffffffffffb00000ffff0000007ffff83fffffffffffffffffffffffffffffff3ffffffffffffffffffffffffffffff9477e7e2f54bd48d59d83506fd30594aa9f3
R2[273] <= 640'hc6ff00000f03ffffffffffffffffff000007f9f0000007ffffe7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff97f674dbcc001640ed87bdceb6ae6c3a04a0
R2[274] <= 640'h1fef70083ff9fffffffffffffffffffe00003f8e0000007ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff59b7dabbb0d7efd5cb8fe0a578244091a1b8
R2[275] <= 640'h7c7813ee3fffffffffffffffffffffff000803000800003ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcdfb67ebb581bf747d5723a3ac0ba8c33e62
R2[276] <= 640'h3817ffcfffffffffffffffffffffffc00c00000000003fffff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff3c59e6f2cd2873fffb917f1e76528ede2c
R2[277] <= 640'h7fffffceffffffffffffffffffffffe04c00000000000ffffc3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb9aadf8be24e013b8e9fe1bb8e217bce3b9c
R2[278] <= 640'hffffffeffffffffffffffffffffffff8ee00000000000e7ffc3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff1cadf54fa1c362a7996bf7d359c5d34d7bbd
R2[279] <= 640'hffff7effffffffffffffffffffffffffffdff10400000000e7ff87ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbf63a95542536026dbadb2567efa1e65581c
R2[280] <= 640'h7ffffffffffffffffffffffffffffffffe3ff8800000000107ffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeed2f9e5ff0e2de27fb3e78ffc5ee88398fe
R2[281] <= 640'h7ffffffffffffffffffffffffffffffffefffe8000000003073fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbf94b2d47bd66d8ea9faefffa18d8396bf4f
R2[282] <= 640'h7fffffffffffffffffffffffffffffffffffff80000000030f1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffada7fb3b9f473541dbab5fd997ff2528e93
R2[283] <= 640'h7fffffffffffffffffffffffffffffffffffff80000000031f07ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc9dedbce2fdede542f91fb23bf29797f36e07
R2[284] <= 640'h880003f7ffff7ffffffffffffffffffffffffffffff80000000073f00ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddcc46c8fe3fcef1ab7cd5bfbee66799bfb3e3
R2[285] <= 640'hcc0003ffffff7ffffffffffffffffffffffffffffff8000000007ff00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcb1d2ef8d55c7d77cdefcd4fe046fb1eff3ff
R2[286] <= 640'hfff0003ffffff7ffffffffffffffffffffffffffffff8000000003fff8ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffe7f3aa25da9f7b3f735ee377c8ba375df39
R2[287] <= 640'heffff0803ffffffffffffffffffffffffffffff7ffffff8000800003ffff1f3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe5795fbe2975e37eef77be4ffa7bd76bedc53
R2[288] <= 640'hfffff8801fffffffffffffffffffffffffffffffffffffc00001000707ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5fbefca3e8cee3ef9eefbc332dbb9a22c679
R2[289] <= 640'hfffff8003fffffffffffffffffffffffffffffffffffffc000e000001fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff77a65f877e80b95ebedffeb37ed51fb9fe66cd
R2[290] <= 640'hffffffff7fffffffffffffffffffffffffffffffffffffc0000f00c1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbe7f735df2f4fc9fbbc4ff9ab7f54d94b9f75f
R2[291] <= 640'hffffffffffffffffffffffffffffffffffffffffefffffc0000ff0c3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff9fedbfd9d9dfec26b8b9e584f87f806f134ffe
R2[292] <= 640'hffffffffffffffffffffffffffffffffffffffffe7ffffc080ceffcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffaffdc6eec1f82ead777fdc057c24233fd2f36d
R2[293] <= 640'hfffffffffffffffffffffffffffffffffffffffffffcffc0c00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc25cdfba71f04c3fdbafcdc7bd11d54e0c3637
R2[294] <= 640'hfffffffffffffffffffffffffffffffffffffffffff0ffc0e00f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdfee565666e1c5cf89f7ad84738aa017c163d9
R2[295] <= 640'hfffffffffffffffffffffffffffffffffffffffffcc1ffc0fc711ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff231bf3b8b391cf37f73ab630e925bb6c53df3
R2[296] <= 640'hfffffffffffffffffffffffffffffffffffffffffe81fffff0731ffffffffeff7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdf5e7fed99b0df1cdf361e7bf75f3e3f9a751
R2[297] <= 640'hffffffffffffffffffffffffffffffffffffffffffc1fffff8733ffffffff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbd872eec89af83e5fe29e6f6be7c7e6391ef6e
R2[298] <= 640'hffffffffffffffffffffffffffffffffffffffffffe1fffffefffffffffff3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff55d3ff7f4ffbfbf6fdf4cfedfc937b501b70
R2[299] <= 640'hfffffffffffffffffffffffffffffffffffffffffff9ffffffffffffffffbefffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffed794a8d29ef67ef97636787e52f85bd547c07
R2[300] <= 640'hfffffffffffffffffffffffffffffffffffffffffffdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7ffffffffffffacffb62c0a875f73edf1f2cf1e97466d2596
R2[301] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffffffffffffffffffffffffffffe1ffffffffffcef3ec8df4c0ace8b6bfda3124759d79e369df
R2[302] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe3fffffffffffffffffffffffffffffffffffffffffffffff67bfffffffffec95b5ff79a669861873fe7290f3427ffffeff
R2[303] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc1ffecfffffffffffffffffffffffffffffffffffffffffff2f9ff3fffffff06a72ef89bbe07eca3f28219dc85f79d25c94
R2[304] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff82f8ffbffffffffffffffffffffffffffffffffffffffffff35b9fbfffffed32abc9e3e656ca1f6b9b271fdb71e0dc9a30b
R2[305] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa02f43c9ffffffffffffffffffffffffffffffffffffffffff7d2efbfffffed683557f6e334f617ecefd317effc1476dd913
R2[306] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc09cf83d9ffffffffffffffffffffffffffffffffffffffffffbd7ee2000001a5ffb8c5cf2a28be11dd9b737de8a56339b8cd
R2[307] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff50360bfdffffffffffffffffffffffffffffffffffffffffffefddb79000fffeb1edfef9696b9e6d0a1b9b3d9fcca76fcf9ce
R2[308] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe795f411bfceffffffffffffffffffffffffffffffffffff3f00003696b2ffffff2339a3e0f4d5741f4faf33a0ee1dd1f4f1c99b
R2[309] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffc07fc6fffee3fffffffffffffffffffffffffffffe00003ff7ffffdacede7fffff33fe5d5cbd6b04ab618557736bffadfcb8eca3
R2[310] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffff800e1f7bfff3ffffffffffffffffffffffff20c00007fc3fffffffd9be72ffffff999fffad85a35445faf8f94873fb8e9ef9e5bd
R2[311] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffc010fe7fffb7f1fffffffffff00000003fe7ffffffffdd87fffff78bfd8ffffff230a7ea940d6e07ff9d71981c73f7edfc499b2
R2[312] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff83e079ffc81fe27fff0000000003dffffffffffffff0dc0ffffff55dedfffffdffde75fab342967e7eeb6ddf2dedaf24260990f
R2[313] <= 640'hffffbffffffffffffffffffffffffffffffffffffffffffffffffffffefe000fffe336387e08008ffffff1fffffffffffffcfbc8ffffffbc0bb9cfffdfdbe94672c3b6eaef3788f6623ecfd8837cf958
R2[314] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffc00083ffcfffff63e3ff1ffffffffffffffffbfffffff6c7bdfffffffeffb9dfffffedfc3fc3e9bcd1acebeafce8d74dff377ebe8e
R2[315] <= 640'hffffffffffbfffffffffffffffffffffffffffffffff000000000007ff01c0201c1c1fe78733fffffffffffffff1fffffff07cfffffdfe909e3dbfffefd1fa2eef77cee08ee73b7a417f73efff77c87c
R2[316] <= 640'hffffffffffffffffffffffffffffffff800000001c00000000000fffffffff800000fff0c380fffffffffffffffbfffffffffffffffcfe4dbafdbfffdff79eed75fc49a0cfbe1cf903272fd01fde73fe
R2[317] <= 640'hfffffffffffc00000000000000000000000000ffffffffffffffff7e0331ff000000fff8302c3ff4e7ff1ffffffffffffffffffffffefe5af337ffffffd2dfa9de736cd68d347dfb087ccabeef7d3af2
R2[318] <= 640'hffffff030fc1000000000000000ffffffffffffffffffffffffff8f8e03b0ff8cf00188c303f8f3f71f773fffffffffffffffffffffe6f69fb837fffe562ecbfb551b0fa0be5d9fd126e292fdfa579ee
R2[319] <= 640'h800000fffffffffffffffffffffffffffffffffffffffffffffffffe0bf7fff1ff8010000fb7677806ffebfffffffffffffffffffff49bdf1baf5fffaccbe6f247c3a8bc391f73201f788f1f7f5bfc8
R2[320] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffc1c30ffffe3fffc000000e800ff01fff8ffffffffffffffffffff65c6ffe7bebffffd2f4d644f0c6485f9f68e20299dd5f379f74fa
R2[321] <= 640'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000e0fe03ffc00000008005ff0ffff01fffffffffffffefcfdb7bfbfd7777ffd9eeb88e769a2033b96d12ef617edf3f35ce666e
R2[322] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff000387fe33f8c0180000007ff00ff00c03fffffffffffe7ccf97f7efdfdd7ffde75f779dd6e78725d7910fac5bbfecfc704f7d4
R2[323] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffef8003cefe13fbcc000000000e480008006e7ffffffffffff94dafe9f6cdbffefefc74ffa77b3f2814f781ae7d27fb9dbdef073ba
R2[324] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffe037fefc1ffffef3000000002000000003bffffffffffbf9cc45fd8a78fdf2485bd9b9cc75f1ea0caca37ad7cbe5ccebdf211e7
R2[325] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8ffffcffffffc00c00000000000000000ffffffffffbfedb27e1fbc560a25cef1fd1fe1b26d6cb95e5afbc808ffcf4da8b186
R2[326] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffff8e3f801000000000f2c8000ffffffffcddd8f9fe2de75acddd9be0d25df9df06db2b6cd36dbabf4513204593e
R2[327] <= 640'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffffe180078b3f0477f3fffffffddaddb7d6bcccdfbedd8a7f45eb6be772666762e9e00b7def9b3fe0b27
R2[328] <= 640'h1c00000000003f07ffffffffffffffffffffffffffffffffffffffffffffffffff0000001000000000000000f400ffffcffffe0795b97fbbcc7f73daf6be7b8071e5d7152a3a172a05f77cbdb9fc2e37
R2[329] <= 640'hc000000000000000070f0007000000000000000000000000000000000000061c000003fefffffff807e0000000000007fffffebf4bee978fb6c7f9da5fea5dc266ee8d0ab5362dc5c07c8c624bde3887
R2[330] <= 640'hffffffffffffffffffff00000000000000000000000000000000fffffffffff9fffffff800000018070000feffff8000fffffeb3ff1c1fde9f0ce94f76efd3f9ef992c1c02a35d7c182dbcf670dabbdf
R2[331] <= 640'hc3803000008000000000ffffffffffffffffffffffffffffffff0080800003f800c000000000fffffffffffffffffffc3ffffe31effb2b939bd35b5de6fe7e9fbf783d3891def73dec48ff76220e1e5c
R2[332] <= 640'hfcffc000000000000000000000000000000000000000000000000000003fffffffffffffffffffffffffffffffffffffffffffc797fdebffc8a7f1a35262e6a7f3e8ff900a788d789cf74ef779da7c25
R2[333] <= 640'hffc7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff23d70fc36b7ff7d50fdffa5efefe346125bcb83c343185f21fffb02b77
R2[334] <= 640'h3fe03ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbc9edb7afa63e3f2be10b247dfedffdef8ac737e9bfc45bf9d6f7367036
R2[335] <= 640'hcff9f3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb9dacd13e5fcaeec7f57a92ed4db4bb53c8c8556b918c075bd39fdaf3bf3
R2[336] <= 640'h7f01cfffffffc7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdc29f25dd58ffe28727eee36fceddb27b85e32937cde841cff77fffe6ecf
R2[337] <= 640'hfff08ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffea9fda32cc9bfcef4ae6b77cd80b3b4e09d24e157de884ffcd5346e495b
R2[338] <= 640'hffffe07f3ef7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddefffaa3fc9ab2f9fb7bb0f656353edc5210afc98bf4c69acebde8b777b
R2[339] <= 640'h3ffff07fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec5be42853a6976c7ddaf9b83bfcb43377c4895a8c688e2128fff9a76be5
R2[340] <= 640'h81003e007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffaf497a2f235333a7fbdae27bdb62e71294eefc2f7f65de6fb47ff3fd6faf
R2[341] <= 640'h80033c1fffe7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff97ffffffffff9ffbf4efabf79bfffdfb7334bcd0ee13f7432d9532f1c335db9d67bc383f
R2[342] <= 640'hb003fe0fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe7ffffffffffffeaad539de5c3efbfd72c9a5ca83b111f229e74b296cd0ca37ec13d2efe
R2[343] <= 640'h1900bfe7f3ffffe7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdffffffffffffffff1fffc37fbdf38ce907079367f67fdd951fe3fcfdfb0d9eb4abbc76d9dfb9f0d1c7f
R2[344] <= 640'h2007e000fff99fcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5fffffffff7ffff7ffffff9bb41f3de5a643aaed7dd5783735f8125eeaf200f70058d31ed537f8c63b35
R2[345] <= 640'h7f0038fe9fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcdfffffffc3ffef00f7e7ffe92e0ddfda7af88ee68c6eb6c06b6b366ec70d1709eb38e1fd83412ac69c3
R2[346] <= 640'h1007e000c077fffffffffffffffffffffffffffffffffffffffffffffffffffffa7fffffffecdfffffffc3003fcffff03fcb7087cdec24efe99b654ffe6f3c358db5f65df57ab33731699d1cea00972
R2[347] <= 640'hfc000003663fffffffffffffffffffffffffffffffffffffffffffffffffffcdbffbffffdfc01fbbff7fffffc1fff7ff4edafff41c56bcbda7fff9aab44bf5364720a7a01f6cdc1a4ed7675a1a94
R2[348] <= 640'h18ffff3e00001fffffffffffffffffffffffffffffffffffffffffffd86ffffa89b7f6ffff9c00b553ffffffffe001bfff02f72cffbbcfc8faff7fe5c8fedfc7ddbe98179e1ec6941bfcdec9c24d91
R2[349] <= 640'h201e7ffffff003ffffffffffffffffffffffffffffffffffffffffcfe6000fffbafdd786fff20c32cdd03ffffffffffbffe0177a5789f7ad97edc7bf9fedfbb7fce4beceb1d46f7c80bddde40509171
R2[350] <= 640'ha000001ffff003f83fffffffffffffffffffffffffffffffffffffc80f000f111f7aa9f07f0bbf0b2dd1bc0ffff7ffffffe2f7b270a9f39e9b7e8c9daec93b6e7fcf70c2ecf91f1440c9f8cf9dc3f3b
R2[351] <= 640'hfff8001f9ffffffffffffffffffffffffffffffffffffffe07000000ee9bde07c1bb0f1f1b9bfe31ffffc7fffffe50a11b4b5bbdb5873f77ac27f257528f83685d8395e62b8f842f30d6355d
R2[352] <= 640'hffc813fe77fffffffffffffffffffffffffffffffffffffffe00043c928f52ea1f9a4b86592003ffffffffffef8d2fb402e7b95c2bffa7cbf3348eb5f3f7f7819968fee4bb3271d18847e30
R2[353] <= 640'h400000003fff00f7ffffffffffffffffefffffffffffffffffffffffffff184d452ffffbef8efffe5cdfffffffffffffffda5659eefe615bcdf95ddfe59e2eb64d4bc5c2c564a052dbf3d2964586d6d
R2[354] <= 640'h400000001ffff8101fffffffffffffffffffffffffffffffffffffffffffff57bfff3f63e7e7fffe5f9fffffffffffffffd7ef412fa6b6fb3f3edce71e9e51e1059fdb1658e718037e5f5d96ca20afc
R2[355] <= 640'h4000000003ffffffc0bf906fffff803fffffffffffffffe3ffffffffffffffbe189f6bf7d1b6f6ff57ffffffffffffffffdf1a4ffa46f458bfdeda79f9dfa07763bbdb40a865de4e742404a8f467b71
R2[356] <= 640'h37ffc7e00c007ffe78fff6ffffffffffffffc08e7feff8fff7eff799d76dcfdde7f1fcbbffffffff9ffffffffee5ede32683ae57ffaabc8ebd776c253f5dd05053cacddb2f4000b55358b
R2[357] <= 640'h200000000073bfe0000003fffc1ffff7dffc0c7ffffffffedf7be1fc7fffffcb0f82d9ff33b4f9fcb78effffff9fffffffee6a490facf23fee3cbe7fcfdcc4729de7c8705008255baf3a40fb0d61062
R2[358] <= 640'hc00000000000033f0fe019ffc1effffff003ffc1fffffffffffbe1fff7efffde7e9bdabff7fbbafebeddffffffbfffffffeff44ace2b7f7a79dbeda6e59254febaeba8d0601ffadab4173538754362e
R2[359] <= 640'h6000000000000014e67ffe463fffff9fffff1c7effffffffffffe3ffe7f3ffb112a692b8f4fdf6f94effffffff3fffffefba6ec55ff70f9bdda3f75aebbdbb3921231bd0286af877e38f739e80b2497
R2[360] <= 640'h5e84000000000003effffffffbca15ffffff83fffffffffff7eecf7ff81fefa9c1159af4e679fc677ffffffffffffffe60ff58cfbc77dfbb3fae5f47d9f48270c5d378335cb13e6d8c620139e0f0e
R2[361] <= 640'hcfa7ed000000000000007fffff0ec0f89fcfff8ffc03dffdf98fefcf0079877fff45d9fdbaede3fb6b3fffffff7ffffff6f7f68be5fbb6e5cbc3f8fdb69a7033ad8455f40e87f81aa30d497b333db4d
R2[362] <= 640'h1a601040400000000000000c0000f80020000ff800788dffff70cf1bfe03fc3df645fe59dd6f6fbfabba7ffffff6ffffff3dbfab4d5dafb5bcfddcef72a6e1b1b74ad097c2c997894012e8be0fd9c108
R2[363] <= 640'h19c0036880000000000000000000e0b0278007ffffe00ffffff087139fb9f01d9b8732f9fdd35fff97b6ffffffe4ffffff66fbfca77ed5fc6ab9447fd3afbadfddef7a46a2311c978034ca3519cc1308
R2[364] <= 640'he80001c000000000000000000000030688003fffe00e3ff7ffe019b8799f026c7ffae2fdd38d82fd27fdbffffa7fffffff6cfe82d7db66bbcf3fcd7fb33e44f35df0d1e21d90a02ed1c5c9f03d77b04
R2[365] <= 640'h150003890030000000000000000000002b0000fffe00009ef3ff7bbe03c07d3fb019dbdbe7751536e33effffff6dffffffcdff7db65c37cd91fcbd76393f332d26532fb7a159c123f0600d0497df032f
R2[366] <= 640'h1c000001f90400000000000000000020520000e3fff89600f0ffff379fe3ffc947b263b3bb6dcb7c8bf6effffff6bbffffefbf796166f96f485e37fbfbf724ff1d783969e9f1b732b25000a001b4167c
R2[367] <= 640'h80000383f76000000000000000000306980003fffff9380043fffad9ffffffde51d77763930e04cdf27efffff3673fffffe193579faf3765f9bf86bfeb8f777e825f2a7c08d850894d012c0441a028e
R2[368] <= 640'h806da6c0000000000000006207212003fffff1ee00123ff749fdffffc354f3c17b696c676387efaffff377fffffb85fefb7f13b7fdbfffcadee443cec70d45d5520401143b500000007052245
R2[369] <= 640'h800935c806400400000000e019030007fffffff0003c3dfd5bdfbdd9d6030e7ac838f5b73dfff7fffef3f7fee7b5f9ff96cb3f7eafaf7516e7ed79f72a8e50449c442c82930c0000326c3072
R2[370] <= 640'h70010702a38001000000002011820007f3ffffff001f3dde31d7bbebfcf5ab7b9c00f5fbffd9fffff9ea77ffffd5f9fb37c14d6f7aafada87eafd2dfa4f16aca90085a91fa0400001b88051d
R2[371] <= 640'h1200011df2100000000000339f07e0007fffffff000ffc302b948fee24fbfc6d94cb561e76d7f3fff9f1ff3ffff77d095fcdf6cf98ed8bfccbd6c37bfdad79deb00023901d2413009b9a0714
R2[372] <= 640'hb0000127dd2040000000714c4e1c32318f8fff00007fe275b079be0d8595f33af73958f77d473fffc7ff7bccd91d738bd8eece79e6c771b7f77672bdf873faee00034007d3b020088de13f7
R2[373] <= 640'h230000006c50000000010c007f00000ffffffff000ffb51ffddac8ab35d3a8e4d352d179cf7f4ffffbf7f8c91e7babb2cbbf9d9bf6db65f3dfefeca2fefa1d4e80013e890c30000063503b9
R2[374] <= 640'hc1000000a2d600000014000180000dc0f8ff0c3fffc7e9e7dcbc8ede839ab73d0fefaf3d03e7fffffefcfff7f75b9a9952ac59dc7bf5f392e73f67c9146465d40111c4a727060000570292
R2[375] <= 640'h1c0f000001a9c0000038000180007e0003f003fff1b2684e4d8c8a3cc1554f2087237ebfefdffcefbcdbfff9cbb32bc03fdc1f3df1f7eedc573a2f8a2530855c000fcc346704000439024d
R2[376] <= 640'h2f81e000028e70008580000f000c3fffb002107fe1ef2c53c88f28f3399c1f9ce2683b28efdfffffb7ff2fdc7cb8ec7bfdeccc5653befe15493c89be03a6c6807198408260800013f01c6
R2[377] <= 640'hfff01f000005dc80180002f07e3fffe1ff81fe618c0be93dba6bf83c7c647360cdd7f9a2effffbeef7fad3c0e9ae36181e6fe5374efffe3fd873aecfc632e80c81e2009b180001000065
R2[378] <= 640'hffffe03c0005b640e80001befffffe070300ff6086e477e46829e7de1e6fde63d0effc1f5ffffffb7fd8db6ec5ba0ce07f6188d7f7c97e8fc8d18ea9ded1b004808a008f180000000028
R2[379] <= 640'h310fffc0380003f60000027ffffff810000001033a2325b0bfbf6dbe10edf44ecfb372ddffffeef96ffadb335deb6656cefdf6efeb54f6e7d4e953e8b3c43003008c0084000000000000
R2[380] <= 640'h1c803ffee0f80009fc0002cfffff800000000001b951a7a2f39cd78a898c64a9f37db9ce6f7ff3ffa7fed8db76d3e147fc71dfcbd1e7776c7093322e8591b80000000000000000000000
R2[381] <= 640'h39fc01cff81c002080002cff7800000100000005a5f602be6e2bc767befeae8a98dfd4ddffffcfee4fbfeccde1440005ba8378173a970f70f978c4de133800000000000000000000000
R2[382] <= 640'he6ff80ffff3f80000002000080000810fec001b7ae9a3eaf039a46f7acc47e6b0efd3bfffffdfe64fe7581e0078008410c0e76bac090b3ec70067ddc00000000000000000000000000
R2[383] <= 640'h307ff9923f9e8400000106c80001118fef1000651981f307d6d528335dc7a38e22ddd0b13fffff7fd7e2b2000800000000f49d19a654709864a89e8000000000000000000000000000
R2[384] <= 640'h1b0fffffc3fff8c3000356d0077ff3c3fd0000567281d7152a1facc9ae93b2b3adad1887dffbfb7fdff6bc00000000000003aefe8e654e4fb9e4f00000000000000000000000000000
R2[385] <= 640'hcf803ffffff9bf03800382443fffffb7c003127c4e82e5e72d1e2dbaed1dff872655a1dbffbff5fb2c3c000000000000000c7c8d43b2fb595a1800000000000000000000000000000
R2[386] <= 640'h20fe007ffffff0fff400007c9fffff9c3009153d4c828c424779e9fbd62a79b142e5ad73ffff6d4e65f0000000000000000f0829b6d02c86027000000000000000000000000000000
R2[387] <= 640'hc7ff0007fffffc7e723f92520ffff0000070dce3a98b0f78e0edcbf74d6bfe7a1647db0fd91e5c719c0000000000000000e0722cce96d3ec98000000000000000000000000000000
R2[388] <= 640'h301fffe10000ff47376394ba0000c0031fb7bffe33ebd837769ab7a45b45ec0a407c1ea24f57863f300000000000000000207a16008a1c1c88000000000000000000000000000000
R2[389] <= 640'h1901fffffff007e0ffff7f2a000000c0e745fde582d4e429f7ffa7e32091b9e771b17ad77fbbbc68000000000000000000a400140008238000000000000000000000000000000000
R2[390] <= 640'h78000000000000ce0007fffff701ffd9f2c070003e0fa4f20bd4064bdf6ab4d763342cc15de9f2286f8eddfbf889f0000000000000000e0481a0801c0002400000000000000000000000000000000
R2[391] <= 640'h6c00000000000023fe0017066bf4067e66bf9001ff09bee804200e42453d1fb9faa928fa8401f87dc5078d7b363c0000000000000000060b61a244400000000000000000000000000000000000000
R2[392] <= 640'h6c000000000000083ff030180007f180ffffe7165e1807e0040000000ec6fa1af67f757f000061f3dad3ffffe00000000000000000000004c00004000803000000000000000000000000000000000
R2[393] <= 640'h3c0000000000000307ffefffff000ffe17ffcfa0f9b83f60000000000017b2e35ed4eff000001ffd35d80000000000000000000000000003c00004000000000000000000000000000000000000000
R2[394] <= 640'hc07ffffffffe001c1f83c4936fd830000000000000001afe0154a8000000000008000000000000000000000000000000c00006780000000000000000000000000000000000000
R2[395] <= 640'h3f0033ff33cff0000ff7ff82e7800000000000c830fd7cb1def7a0000000000000000000000000000000000000000000182006780000000000000000000000000000000000000
R2[396] <= 640'h1ffc000000000fc7003ff8e008303ffffc8000c1ffffc83dc8ce0c000000000000000000000000000000000000000000182476780000000000000000000000000000000000000
R2[397] <= 640'hc3f800000120027fc01f26863e03ffe0fc000c9fffd6005100040000000000004000000000000000000000000000000182476000000000000000000000000000000000000000
R2[398] <= 640'h301f800003ff00073f8067402703830000000fb00097cd0040000000000000000000000000000000000000000000000dc3030000000000000000000000000000000000000000
R2[399] <= 640'h2031cfff0fffe4001f88be43303880060002030005c430040000000000000000000000000000000000000000000100fc0030000000000000000000000000000000000000000
R2[400] <= 640'h1000003300007fe0009ffff00028000600020300c9fbe80000000000000000000000000000000000000000000000002821e0000000000000000000000000000000000000000
R2[401] <= 640'h4c00000000001fff907fffe103800060001f33fe9ffc8020000000000000000000000000000000000000000000000082000000000000000000000000000000000000000000
R2[402] <= 640'h47e0000000000007f920fff003fc0000001f33ffcfcf8020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[403] <= 640'h1079000000ffc00003fffff803018000000d12ffc02e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[404] <= 640'h501ff1cffffffc0000ffffc0001c000000003fce0060000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[405] <= 640'h110000ff8f8ffffff003fff80000000000003f800060000000000000000000000000000000000000000000000000000000003c00000000000000000000000000000000000
R2[406] <= 640'hc0000000000003fff801ff400000000000017000060800000000000000000000000000000000000000000000000000000003f00000000000000000000000000000000000
R2[407] <= 640'h3c000000000000000bc4cfd80000000000000000040800000000000000000000000000000000000000000000000080100003500000000000000000000000000000000000
R2[408] <= 640'hee00000000000000021fffa0000000000003000060000000000000000000000000000000000000000000000000000110002600000000000000000000000000000000000
R2[409] <= 640'h31f00017e3cffc000001fff8000000000300400000000000000000000000000000000000000000000000000000000000003600000000000000000000000000000000000
R2[410] <= 640'h86877c7e1c00ff8e00071c20000000000e0008000000000000000000000000000000000000000000000000000000000002820000000000000000000000000000000000
R2[411] <= 640'h100000106c0ff0f983800000007400000000000000000000000000000000000000000000000000000000000000286c000000000000000000000000000000000
R2[412] <= 640'h800000000000000001fe7fe2400000001b400800000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000
R2[413] <= 640'h600000000000000000023fb0c000000003500900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[414] <= 640'h18f8000007319f00000001c400000000002203c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[415] <= 640'h408edb3ff0103800c3d17f90000000000380040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[416] <= 640'h4000000000000000001c7e4501000000046000000000000000000000000000000000000000000000000000000000000470000000000000000000000000000000000
R2[417] <= 640'h40000000000000000000001ac2000000010400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[418] <= 640'h38000000000000000000000800000000005600f00000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000
R2[419] <= 640'h7e0000001fe01800000066f000000000004a02c00000000000000000000000000000000000000000000006c0000000000000000000000000000000000000000000
R2[420] <= 640'h337ff8c100000000000081040000000000328090000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000
R2[421] <= 640'h9002000000000000000000600000000000a800a000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[422] <= 640'h42000000000000000000002800000000002cc01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[423] <= 640'h8080000000000000000004a000000000003200c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[424] <= 640'h60600000018000000000002800000000000860300000000000000000000000000000000000000000000000200000000000000000000000000000000000000000
R2[425] <= 640'h1cf00000000000000000000100000000000594000000000000000000000000000000000000000000000003700000000000000000000000000000000000000000
R2[426] <= 640'h6b800000000000000000000c0000000000061000000000000000000000000000000000000000000000003f00000000000000000000000000000000000000000
R2[427] <= 640'h300000000000000000000008f078c0000000e000000000000000000000000000000000000000000000003e00000000000004000000000000000000000000000
R2[428] <= 640'h400000000000000000002007ffe0c66e000a000000000000000000000000000000000000000000000000828000000000004000000000000000000000000000
R2[429] <= 640'h1000016000000000000000047fff00fc0000000000000000000000000000000000000000000000000003060000000000000000000000000000000000000000
R2[430] <= 640'h200c01880000000000000000ffffc3f8000000000000000000000000000000000000000000000000007000000000000000000000000000000000000000000
R2[431] <= 640'h1dfe000000000000000000000ff0f818000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[432] <= 640'hc0000000000001000000008df3c3800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[433] <= 640'h300000000000000000000004ff00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000
R2[434] <= 640'hc000000003c0000000001f80000000000000000000000000000000000000000000000000000000000c78000000000000000000000000000000000000000
R2[435] <= 640'h8000ff7cc000000000fe000000000000000008000000000000000000000000000000000200000000030000000000000000000000000000000000000000
R2[436] <= 640'h7d1fe00000000100fc00000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000
R2[437] <= 640'h197e0000000003fe00000000000000000000000000000000800000000000000000000004c0000000000000000000000000000000000000000000000000
R2[438] <= 640'h6000000001eff000000000000000000800000000000000000000000000000000000000380000000000000000000000000000000000000000000000000
R2[439] <= 640'h1000000e7ffc0000000000000000000fdc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[440] <= 640'h4103ff7ee000000000000000000000fc00e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[441] <= 640'h303cff200000000000000000000000787f60000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[442] <= 640'h87f80000000000000000000000000683fc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[443] <= 640'h3fc000000000000000000000000007c7f80000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[444] <= 640'h3e4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R2[445] <= 640'h12000000000000000000000000000000000000000000000000000000a000000000000000000000000000000000
R2[446] <= 640'h2000000000000000000000000000000000
R2[447] <= 640'h1e00f3100000000000000000000000000000000
R2[448] <= 640'h60000000000000000000000000000000000000000000000000001800000000000a0e460c00000000000000000000000000000000
R2[449] <= 640'h200000000000000000000000000000000000000000000000000000c00000000001985f00000000000000000000000000000000000
R2[450] <= 640'h6e0000000000000000000000000000000140000000800000000000300000000210384400000000000000000000000000000000000
R2[451] <= 640'h6e00000000000000000000000000000000600000000000000000001400000000f0080000000000000000000000000000000000000
R2[452] <= 640'h80060000000000000000000000000000000000001c000340000000000000000000000000000000000000000000000000000000000000
R2[453] <= 640'hfc00000000000000000000000000000000000002033000040000000000000000000008000000000000000000000000000000000000000
R2[454] <= 640'h7e800000000000000000000000000000000000006086401810000000001fc7000000000000000000000000000000000000000000000000
R2[455] <= 640'h60c000000000000000000000000000000000000140019c0018e07f3100000c000000000000000000000000000000000000000000000000
R2[456] <= 640'h6e00000000000000000000000000000011803800000023ff00c70d9e7cc7cb0000000000000000000000007c06e00c0000000000000000
R2[457] <= 640'h60000000000000070105e280000ff1c001801e80000678003f72b4e00401e6000000000000006040001fffe000030e0000000000000000
R2[458] <= 640'h91bc8f738781ff180000003800007ffff0000035b8301c280000000000000c42801ffffe00000000000000000000000
R2[459] <= 640'h1000000000000000000000000000000000041880003ff8000000000000000000000000000d800c03a7800000000400000008000f3c7c00f0000000000000000000
R2[460] <= 640'h80000000000000000000000000000000000004400826504fb83080010000400602c6080ffff7c001c000000000000000000
R2[461] <= 640'h8000000000000040000000000000000000000000000000000000000000000000102000f9419e0000320800100044006c7c24007fffe60008000000000300000000
R2[462] <= 640'h8000000000000140000000000000000000000000010000000000000000000019f3203f0c40e4380024948000004481766404000000e600c0000000000100000300
R2[463] <= 640'h12000000001000000400000000001f2f800000000000000001d7fccfe520033c000187f38800440807e6c6c00ffefe00100000000000000000000
R2[464] <= 640'h7200000000000000042001041e080000000000000000000000ffff3dac0008e80001a18138004000062042c00fc000000c0000000000000000000
R2[465] <= 640'h200000000000000000000000000000000000261088000000000000000000000000000bff7ef00000077bff094d61d00e02001e3c6703f80700001e001810000c01c00000
R2[466] <= 640'h10000000000000000300100000000000000000000000000000000000000100800000000000000000000000000000000000000000300da5cddc50c02003f380701ff07cc007c000018000000000000
R2[467] <= 640'h7ff04400100000000000000000000000000000000000000c01780000000000000000000000000000000000000000000123fb000000000000000000000000000000000000000000
R2[468] <= 640'h1fff94ec0fac00000000000000000000000000000000000084018e00000000000000000000000fffffc000000000081c020018200000000000000000000000000000c00000000000
R2[469] <= 640'h10001fff067ecb900000000000000000000000000000000000008400ed00000000000000000000000f0003400000000000e9870dfee400001c000000e00c1f0000001000400000000000
R2[470] <= 640'h3fffe47fcc8000000000000000000000000000000000000080007a20000000000000000000000400000000008000000094b4001bc1000938c700e000780000180400000000000000
R2[471] <= 640'h103ffffffe470000000000000000000000000000000000000000000043fc3000000000000000000000780008000f01c00000002c01880c100013040000080000007c089d0480007d00e00
R2[472] <= 640'h3f00000000ffffffffff6300c00000000000000000000000000000000000000040007fff00000000000000000000073ff9807601460000000007e0010800042062000c5682231980492cc00353e80800
R2[473] <= 640'hfd800000c7ffffff3fffe700e00000000000000000000000000000000000001000003fe00002000000000000000001007d003981e0000000000007016a00001880000000080cc90770717c0363000000
R2[474] <= 640'hef0000cf47fffffeffffe700000000000000000000000000000000000000001000001f7800000000000000000000037fc00e3901e00000000000001e23c0000000000027f10f83fe0800f60010000000
R2[475] <= 640'hffffffffc7ffffffffffe910000000000000000000000000000000000000000000001f400000000000000000000006c0060239600000000000000000602000000001c1e00008080010050e0000000000
R2[476] <= 640'hffffff4fc7fcffffffffe200000000000000000000000000000000000000000020001f9c1c0001f0000000000000078000031fe0000000000000000000000001813800002ee9463c003b810000000000
R2[477] <= 640'h1000007c3ffffffffffc800000000000000000000000000000000000000000040001f80220002080000000000000000000099000000000000000000000000015274f0e5df050c034c03c100b800000c
R2[478] <= 640'h3ffe3fffffffffb800000000000000000000000000000000000000000004000008000000270000000000000000000006000000000000000000000000000805a075ff00e01efc0000000b30a000b
R2[479] <= 640'hf000e17fc1fffffffff0018400000000000000000800000000000000000000002000000000000178000000000000000000000000000000000000000000000000002d3fd888008fc000b0009026c40a00
end
always @(posedge vga_clk) begin
R3[0] <= 640'h10000000000000000030000000000000180000008000000000000000010004c3ffe366ffdffe7fffff78fff7fffffffffffffffffbffffffffe7ff07997f8e033f81fffc7fe3613900000000
R3[1] <= 640'h4006000400000000000000000000000000000000000000607ffff67ffdfefffffff7ffffeffffffffffffffffffffffffffcffffe9fff8f1f7ffffffffff0e08100000000
R3[2] <= 640'h8c00e000e0000001008100000000000000000000001800061fff7fc3ffffe7fffffeffffffffffffffffffffffffffffffff1ffffc7ffe8f7fe7fffffffffcf8c000000000
R3[3] <= 640'h80000000800000000000000000c00060000000000000000000000000000000000801063ffffc99fffffcfffffefffffffffffffffffffffffffffffffffcfffc7edf9f7fe7fffffffffcdc1c00000000
R3[4] <= 640'h8000000000000000018000000000000600000000180000000000000000000000010100e3fffe99ffff7effffffffffffffffffffffffffffffffffffffffffff7e9ff0ffffffffffffffdc3803000000
R3[5] <= 640'h8000001f0c03070000000018c000000000000000000000010300e3ffdebfffffffffffffffffffffffffffffffffffffffffffffffffe77ffff0ffffe7fffffff78c6181000000
R3[6] <= 640'h31078c00070031070100c10000000000000000000089039dffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff33ffffffffffffffffe3d0000000
R3[7] <= 640'h2100c600660079870300e3000080000000010000039c039d3ffffbe7ffffffffffffffff7fffffffffffffffffffffffffffffffff9f3f3fffffffffffffff73fc09000000
R3[8] <= 640'h100000003f9c300cf3c831e600e000000000000000000c00007fffff3ffffffffffffffffff7ffffffffffff7ffffffffffffffffffffff7fffbff3ffff7ffffffeeefc08000000
R3[9] <= 640'h10000002099df03033e071e600e00000000000000010000e0e0ffffffffffffffffffffffffffffbfffffffffffffffffffffffffffffffffffbffffffffffffffffefe80000000
R3[10] <= 640'h183c0003749f3c1f31c33fff600c00000000000000210107f007ffff7fffffffffffffffffffffffbffffffffffffffffffffffffffffffffffffffeffff7fffffffffff80000000
R3[11] <= 640'h183c000f669f7cfff3e17fef6404f000800000000020030fff0ffffffffffffffffffffffffffffcfefffffffffffffffffffffffffffffffffefffffffffffffeffffff80000000
R3[12] <= 640'h187e000f67f97bffcf7ce7e3660cf8000000000000000ffffff0ffffffffffffffffffdffffffef8fefbfffffffffffffffffffffffffffffffeffffffffffffffffffffc0180000
R3[13] <= 640'h99ff000fe7f9f3ffcefce7f3668c7c000000000000081ffef8fffffffffffffffffffffffffffefcbff3ffffffffffffffffffffffffffffffffffffffffffffffffffffdc100000
R3[14] <= 640'h1dfff8183f9fff37ffffeffff66fc3f80000000000001fffff80fffffffffffffffffffffffffffff1ff7fffffffffeffffffffffffffffffffffffffffffffffffffffffbc810000
R3[15] <= 640'h800000000000003dfffc3c0b99f7b1fffffffffe6fe3f80300000200023feff9ffffffffffffffffe7f7ffeff7fc7ff96ffffffffff3fffffffffffffffffffffffffffffffffffffffffff1c818000
R3[16] <= 640'h100008040187b0bffc78ffcffff9ffeffffffffd3ff1e99001800600006380f3efffffffffffffff9ff9fffbffc7e1f1ecffef97f3b7fffffffbfffffffffff7ffffffffffffeffff7effffe3708000
R3[17] <= 640'h1000000800073f1fffe9efffffeffeeffffffff997c7f99000000600004813f7fffffffffffffffffff9ffffffe7e1f3ffffffb7ffb7bfffffffdfffffffffffffffffffffffefffffffffdff0fc000
R3[18] <= 640'h1008773f1fffefefffffefbefffffffffbffef9fb00800020008083ffffffffffffffffffffffdffff9fe00c13f3c9f19fcf973f8ff7ffdfffffffffffffffffffffffffffffffffd7ccec000
R3[19] <= 640'h620080000007733ffffffffffffffbffffffffffffe7fb661800800080001dfffffdffffffffffffffffffffc03e00c0e138df90fffcfbf8fffffffffffffffffffffffffffffffefffffffffecce000
R3[20] <= 640'h66008030011cff7fffffffffffff7fffffffffffffefff663800c10380073ffffffffffffffffffff6ffffffc33f00c00001fe900f9cf1fcffff3fffffffffffffffffffffff7bffffffffffff8ff000
R3[21] <= 640'h4008070801cfff9ff7ffffffffffffffffffffff77fffe63800c1633c17dfffffffffffff7ffffffeffffff67ff00800083fc11071900fcffff7ffffeffffffffffffffffff7fffffffffffff8f3000
R3[22] <= 640'h880020c0c03efff9ff7ffffffffffffffffffffffffeffeee00800623c33fffffffffffffffffffff9ff777f66610000008600010331000099cffefffeffffffffffffffffffffccfffffffffffc1c00
R3[23] <= 640'h98003083e0fffffffff7fffffffe7fffffffffff67fcfbfcc0803c7cc371fdfffffdfeff66efdec799ff6778600000003186000080f18700998f76ff1fffffffffffffffffffdfff7ffeffffff7f1c00
R3[24] <= 640'hc0ccef0c03f8ffffffffffffffffffffeffff7ffffff3fee383cc387ffffffffffffbffefffe33c79c7c8c0000000010000000000990000fe0f3bcfc7fffffffffffffffcff3fe7fff9ffffffffffc0
R3[25] <= 640'hf8c0dce0f83ffffffffffffffffffffffffffffffffffffff800ff3cfffffffffffffbfee7fc7c666dc780380000000000010000009900007c1e998e0f7fffffffffffffffffff7fffffffffffffff80
R3[26] <= 640'hfcc1fcc0fffffeffffffffffffe7fffffffffffffffffff37838ff9ffb7ffffffffffbf861383ce70984010800000000000000000080000000008c1c187dff3fffffffffffffde3fff7ffffffffffe86
R3[27] <= 640'hcf83f8c0fff7ffffffffffff1fc7fffffffffffffffffffbfc38dfcfffffffffffffff003138383c400c008000000000000000000000000000000d0c1801ff7fffffffffffdece7ffffffffffffffcc6
R3[28] <= 640'h871cf3e0fffffffffffffffffc1ffffffffffffffffffffeff0f8fc4fffffffffffffe0030c00018000c0080000000000000000000000000000019c700c3fff3ffffffffffde71ef7ffeffffffffffe0
R3[29] <= 640'hc0f8e7ffffffffffffffffeff01cfffffffffffffffffffeff078fc0fffffffffffffe0030c00081000000000000000000000000000000000000f1c703c3fbf1fffffffffcff73c73ffffffffffffffc
R3[30] <= 640'hfcf0dffffffffffffffffe4d03001fffffffffffffffffffffc7cff3ffffffffffffe60000000081000000080000000000000000000000000000d08401c771c7fffffffffe7f73ff3fdffffffffffffc
R3[31] <= 640'hffe3deffffff7ffffffffe48e101fcffffffffffff7fffff7ef8ff7fffffffffffff4600000000004000008000008000000000000000000000188808009e3187ffffffff3f31073ff79ddfffffffff3c
R3[32] <= 640'hfff9bffffffbdffffe8e242040030223ffffedfefffee7ffff7e7ffffffffffffff180800100000000000000000400608100000000000000810007628000f83ffffffeec96b9fcbff3c7f7fffffffffc
R3[33] <= 640'hfffffffffffffffefec4800000000c04ffffeffefffffffffffffff7fffffffff300800000000000000000000000000601090000000000000000006080810ffcff00ffee9639fc1ffffefffffffffffc
R3[34] <= 640'hfffffffffffffffeffc0800000000c0cffffeffffcffdfffffffcff7fffffffff1800000010000000000400000800000100900000000000000000020008107e08e0fc306923880011c7cffffffffffff
R3[35] <= 640'hfffffffffffffffff3000100000080047ffffcfffcff9ffffffffffffffffff97c8000000007000000000000c0800000006900000000000000000000000800c084ffc106920100018e3f77ffffffffff
R3[36] <= 640'hffffffffffffff7ff3000100000000033fc0fcffe7e7fbfffffffffffffffef03c00000000c000080000800000000080e069000000000000000000000018c0030000006010c100018707ffffffffffff
R3[37] <= 640'hffffffffffffffff710000000000000333c04d3fe7f773fffffffffffffffef80300000081c000880000000000010000634d008000010000000000000000000321e018601043004283c0feffffffffff
R3[38] <= 640'hfffffffffffffff10000010000800000337c4f3fe7e066fffffffffffffffe8c01000000c303028900000304c01e0499674e800000000000000000000000000000ff00200000000003004effefffffff
R3[39] <= 640'hffffffff7ffffe730c0081000000010023fe4d3f38c066cffffffffffffe9f8c000000013f3880d918403084033c84f8604ec000e30000000000000000000000000001000020000001007effcfffffff
R3[40] <= 640'hfffffbfffcffe7ff00036004c060000001000000c00c00fffeffffffffff38e0000001803f67fffec31c0073fffe19ffceff71e03c66e7980000000000006000000000800000000000713c1cfefbffff
R3[41] <= 640'hfffffffffffff39900010600f06060000000000080c0001fcfffffffffff30000000303cff7effff80c3013ffffcbbffcffff1e1c16700180000000000000000000000000000000000301f3effffffff
R3[42] <= 640'hfffffffffffff8010000660078980000000000000101001fcfffffffffef80000000383fe3fffffffee7831ff9fcff7ff3fffff3e0673c008600810000000000000000000000000000008307bf7f7fff
R3[43] <= 640'hffffffffff1f38000000e00307990600000000000003000ffffffffffeff8000000603e3e3fffffffff7878ff0fffffff3ffffff7c67ff008f000800000000000000000000000000000083001f7fffff
R3[44] <= 640'hffffffffff0fc3c000076f031f99d8c000000000000000077ffffffffcff8000006703e3fffffffffffe1ecefbffffffcfffffff7eefff0901001800420000000000000000000000000000000fffffff
R3[45] <= 640'hfffffffffff8c300000fff037cfffe8401000080002000007ffffffffeff800000e73cfe7ffffffffffc1cfefff7ffffffffffffefef7e993100c100400000000000000000000000000000c101ffffff
R3[46] <= 640'hfffffffffcf88000000ef899f8ff7fc60000000000000007f3fffffffff7000006fffefefffffffffffe1cffffffefffffffffffffef18d978ff8100000000000000000000000000000000e021e7ffff
R3[47] <= 640'hfffffffff81e8000031e9f9de37ff3e00020000000000007e3ffffffff070000077fffdfffffffffffff0fffffffeffffffffffffceffff99cff18381000000000000000000000000001000071c3ffff
R3[48] <= 640'hffffffcff4000c00034fffffff7ffffe990800010004000fc0ffffffe77c000103ffffffffe7ffffffe7fbfffcff3efffffffef3cffe79fffff8f8fe0000000100000000000000000100000001feffff
R3[49] <= 640'hffffffcce080040000cfffffffffffff998000100000000f1fff7ffdfff000087fffffffff77fffffff7ffffffffeffeffffffee86e3ffffc33f9be00000000000000000000000000000000001ffffff
R3[50] <= 640'hfffffffc2360010000cffffffffffffffc8001100000001f3fff7fffffc10018f1ffff7fff7fffffffffffffffffffffffffffce8673ffc7ff078300f00000010000000000000000000000030087ffff
R3[51] <= 640'hfffffefc21200080004dffffffffffffff0001000000010ffeffffff7ec0008121fcf7ffff7ffffffffffffffffffe7ffffffffeff3fffe7ffe3d1fff0000000000000000000000000000001000fffff
R3[52] <= 640'hffe7feff61001000017dffffffffffffe730000200000100ffffffff3c000003ffffe7fffe87fffffffffffffffffefcfffffff9ffffffffc3f1f8fff8000001000000000000000000000000003fffff
R3[53] <= 640'hffe7fffff000180c00e9ffffffffffffff3899780000000007ffffe73c1800063fe7fe0ffc8e9f99fffffffffffffffffffffff9fffffffeffffbffefc000000000000000000000000008000003fffff
R3[54] <= 640'hfffffff1e000080800f9fffffeff9f7fffd19940000000000fffff660000000e7f71fc8ffc988199e79ffffffefffffffffffffffffffffffffffffefc0c0000000000000000000000000000033fffff
R3[55] <= 640'hff7efff1ce808081007dfffffefe9f7fffc1ffc6000000001c7fffe700000006fffefcfe0c1880f983993fffffffffffffe7fffefffefffffffffffffe840000000000000000000000000000c30fffff
R3[56] <= 640'hfffc9d7c0300048388ffff7ceefe00cffefff3ee0c040090771ffcfc00000c0effff03180000600621ff7fceffff7fffffffffff7fffffffffffffffff3000000000000000004000000000000c7fffff
R3[57] <= 640'hffffdffcf0000000890fffff7fe78cc7ffffffee06c000013ffffcfc0000000fffe7fc800000400022ffd7c4ffffffffffffffffffffffffffffffffff400000000000000000000000000000007fffff
R3[58] <= 640'hfee7fffef0000000037fffeffee78cf1fffffefe07c000013fffffe00000018ffffffc400000000000c3810087ffffffffffffffffffffffffffffffffc1000000000000000300000000000000ffffff
R3[59] <= 640'hffcf66ff0380000003ffffdfe3ff00717fffffff73040000e3ffffe0000001ffff7f0860000000000003000103ffffffffffffffffffffffffffffffffe1000018000000010000000000000000ffffff
R3[60] <= 640'hff1c66ff03008000037ffffe03ff000f07ffffff793c0000e3fffee0000000ffff7c016000000000000000217ffffffffffffffffffffffffffffffffef8000008008000000000000000000001ffffff
R3[61] <= 640'hff3c7ffff010800003ffffff3de30104effffffff96000007fbf3ee00000017ffff3e04000000200000000607ffffffffffffffffffffffffffffffffe78000000000000000000000000000003ffffff
R3[62] <= 640'hfc38fbeff000000046ffffe3f8c001c0ffbfffffffe000007cff3ee00000077fffe0e00000003200000000003fffffffffffffffffffffffffffffffffff000081013100003800000000000001ffffff
R3[63] <= 640'h7cfeb9ef03000008efffff339d38800006997b7fffef0000f3ff87e0000007fffffc00000103326e000000001f7ff9ffff7f3ffffffffffffeffffff7ff700107f03317e803f04000000000001cfffff
R3[64] <= 640'hfffc83078c00001bffff87237e610140087f1fffff9f80013fffffff80003f7ffbc60000300000f00100000020f1fe7dffff7ffffffffffeffffffffff7ff1c00080260020803000000000008133ffff
R3[65] <= 640'hfffe01038c00001b7ffb3c603c01000000001fffffdf80017bfffff000000ffff8e60000030701030000000021fffeedffffffffffffffffffffffffffff9dc00080e0002000000000000000000f3fff
R3[66] <= 640'hcfff00c000000019fffff84000000000000007effff3800070ffff00000027ff8020000002c1fb0100000000010f7fedfff7ffffffffffffffffffffffff9f06009806007018000000000000008f03ff
R3[67] <= 640'hfff300e000000009ffffc10000000001000027fffff1000271ffff0000083fff0020040000e0ffe00000000003e77fedff0fffffffffffffffffffffffffdf1f00980700000c000000008000000f03ff
R3[68] <= 640'h3ee780e000000001ffff0000000000100000067ffffc000203ffefc0001c3fff00200400030fff7e0000000013efff7dfddfffffffeffffffffffffffffff93fff9ff0e1f80700000000c00000330f7f
R3[69] <= 640'h1ecf80c000009080ffdc3c00000000830000027ffffe000003ffefc0000f7fff00000400020fff7e00000000138fff7dfcfdffffffefffffff7ffffffffff97fff9f99e1fec78000000000000031bf7f
R3[70] <= 640'h8f8e83030000008fffcc1800000000800000017fffee0000001f7600000fffdf0000060090e0fffe00000000008fff7fffc0ffffffeffffff87f3cceffffffffff9f1f70ffff00000000000000339fff
R3[71] <= 640'hc78c03070000018fffccc000008000108000417fffc60000000f7e00000ffee004010f008603ffee80e0010000cfff6fff03c3fffffffff970733cce9fffdfffffdff878ff7e210100000000008e07cf
R3[72] <= 640'h90180760000000f3ff380000000001000001061f73fec000003f9900033fff38030031300f39fffe3f1c00081c7673fe79b1fe7fffe7ffffff8fff011fffffffcfffce03ff9c0c030c0000000083083f
R3[73] <= 640'h999803740000013f78f00100000000000000001f7cfe3c00003f9900003fce0000003b00003bffff800000000367ffffff817fffffffe7df1f3c00017fffffffffffcfb7fffe0000000000000003003f
R3[74] <= 640'hb98637e0000033ff3f0008000000100000400213fff3c380000800000ff800001803880007fffffe1c080008107fff3f7a43ffffb7e000e00d80000ffffffffffffffbffbff3000200000000033033f
R3[75] <= 640'hff1637e000003e77f9c008000000100001c6101cfffc3fc0000c00001ff0000008000c00327ffffffc080000c03ffffe18c3fffff7e3c8000c00000fffffffffffffffffffff000000061000033833f
R3[76] <= 640'h7e7266200001fe7fc180130e000c000801e6102c7ffe7fe0000000001ff000000000c170087fffffff8010000007ffefc083fffdfff38c0000000001ffffffffffffffefffffc00060071000030033f
R3[77] <= 640'h26e6246000001f7fe398083038008000013e40063ffffffc00000000087e000000007f30000fffffffff300080407ffefc103fffcefbc1c0001800000fffffffffffffffffff8c0084007000003800ff
R3[78] <= 640'h60006000001f3fe380007b3c000f00c07f800030fffffc00006000187e00000000dfe0000fe11fffff00008000fffcf0011ffffefb81000000000003ffffffffffffffffff000080001800008e00ff
R3[79] <= 640'h240060000007fff98100ff3c0188830c7f8031e1fffffc00006000017c800000038f8f833fe038ffffc0000c03eef1c0011df9fbf93c000080000000ffffff7fffffffffff31bf03001c00000600ff
R3[80] <= 640'h1000f08000cc7fffc00077f9fc0f8f1c3ff0000021f7fde00000000037e000000107fffe3ffc000fff900000000ff9c20000399f180808000001c00039dfffffffffffefffffc73ff99a000000003ff
R3[81] <= 640'hc0000000000cdfffc7000fffff8f7fffe17f000000bf7ffc0000000003fe000000123ffff3ff8000ffff80000000e7c600000098ce8080000000c080011ffffffffffffffffffefb07990000000003ff
R3[82] <= 640'h80000c3ffee4001fff7fff3f3f3c7f808080fdfffe000000000afc00000092fffefcff00000fff80000010c38000000066ce80c0008000c000002effffffffffcffffffffc83f90000000030ff
R3[83] <= 640'h1800080000c7ffff800ffff7ffefe3f1effc00080fef7ff0000000002f800000092ffe6fcfe00800fff80000000400880000027e10fc00fc000fc000066ffffff7fffc3fffffffefff90000000023bf
R3[84] <= 640'h10cffe700001fffdffcfc7f0ffec000002ff9bc8000000103f8000000b29fe6deff00003fef81000000180000000026713ce01fc000fce00026ffffff7ff8007fffffffff9f0000000003bf
R3[85] <= 640'h10cffffc0001fffffffffffcfff80000006197e8000000003f800000037fffeffff00000fe68000000018000000000031387107c000e7700006fffffff97c017fffffffffbf0000000003bf
R3[86] <= 640'h6dfffec0803fffffffffffffeec0600000017f800000000ffc60000136ffffffff030001fec000000000000400000003017103d001ef3f000087c039f0000137fffffffff900000000103f
R3[87] <= 640'h8000000669ffff0098ffff63fff37fffffc0708100011e800000003ffc300003367ffffffe070007fe6080000000012c8000008e017183c083ff31000000c018030021033ffffffff800000000383e
R3[88] <= 640'h21004000417fefff00c6ff630fffc7ffffff99e160000067c00000009ff83880009bffffefff00c006ff991883000084e7000000643ff1cffc413cffe1801830030c00010007fffffff720000000703f
R3[89] <= 640'h7ffff0004fffffe7fffffffff7ff600000002fc00000009ff03e80cfbbffffffff000018ff03000080001ffe0000000000f001fc009efff0801820c00400000063ffffffff00000000003f
R3[90] <= 640'hc7ffff00067feffc067ffffffcfff7f2000000ef800000effe0f40001fbfffffffe010c1c7f60c3fee0187ffe00000000000001ff00defff8800000000000000000f8fffffe04010000041f
R3[91] <= 640'hf7ffff800f3fe000367ffffffcffffff000000ffc0001ffffe0f4003efffffffffe010c0f7fe0e77ff9387fff10000000000001ff407fffffc00000000000000000f09ffffc8c000000061f
R3[92] <= 640'hcf7ffef801fbfe000167fffffffffefff8088007ff0000ffff007f393effff0ffffe008c07f367ff3ffff7ff3ff0000000030001f3003f1effe0000000000000000081b9ffff8cc00000061e
R3[93] <= 640'h4dfffff803fefc000080fffffcfeffff80000003ff8000ffff007f3f80fffffffffe0080049b67ff7fffffff8ef000000003040171007f983ff0000001000000000003b8ffff88c00000061e
R3[94] <= 640'h79ffffe003bffc000090fffff9007fff90000003ffc000fffdc1fd7fe7fffffffffe0000803ff9ffffffffff87e0000000010c047100ff080ff000003100000000000067fffc98800000003e
R3[95] <= 640'h40010000613fffe003ffc0008098ffff91017e7ff9800080ffe81cfffd80157ffffc7fffbeff0010003fbbffffffffe31fc000c018008e847800bf0c07f000800301180000000047ffffb9000000019e
R3[96] <= 640'h1b000001d7ffe700fff8000000cffc038c11fffffcc8027ffff0fffff00fffffff3cff9ffff6000cdffbffefff3e0008ff80000383308817b00fe420fe600000001010084005803f6fffc8000001807
R3[97] <= 640'h97fdfe01fff0030e0009e00000008feffcc8002fffffcfffc00ffff8f70873fffff601e093ffffffc7100008ff8000000711e997b80ffe09fe400800000000001000002eeffff8000000900
R3[98] <= 640'h4677fcfc01fff0078fc000000008000787ffc0103fffffefffc80ffff9f00031fffff013c0001ffc7fc2000000ff000000870fc1cffc0fff8effc00900000010021000000ffffffd800000338
R3[99] <= 640'h6e7ffcfc03fff007ffe0000000301003b7ffc0003ffffffffce00ffff1c0001dfffff002000036ffc6600000003f000013ff1f83cffc1fff8e7fc80011800018003800000fffffbd800008110
R3[100] <= 640'h667fff7007efe00fffc20000003100003ffff0001ffffffff8400effe980000ffffff000780016ff02700000000f800203fc3fe7fff997ff966fe6107f80063808e8000009fffffc080000001
R3[101] <= 640'h63fffc00fffe00fffc30003901e00003fffde001ffffffff8003fffcc000000fffe00107800065c100013c030378000007c70fe7ff787ef9efff730ff338f3fcde8300009ffffec180000403
R3[102] <= 640'h10000001fbffc000fffe03fffe60003e1ff000008ffdec00c7ffffff8007fefc8000002fffc00040000060810003ff8002fe000003ff0f67fff007fc8ffff37fff3ffffffec280009dfffeccc0000600
R3[103] <= 640'h80000019ffdf0000effe03ff7fe0001e8f3c00001cfdce01837fffff003feffe180000663fc00000000060000003ff8010ff0000e7fce077fff107fc811fdffffffffffffffc800099fffff8c0000000
R3[104] <= 640'h1e7ffff80007ff603fffffe019ecfd8001000fffc03003fffff003ffffc40000e1f4920000000000000803ffe1900ff00003fcef27fff80078101fffffbffffbffbffc000821cffff80f000000f
R3[105] <= 640'hfffff80077ff607fffff0101e4fff3e0000fffe30003ffffc0067ff4800000007e9000000100c0000b8ffff99e01f80007ffef23fbfc00398000ffffffc7ffffff8e000000effffc1f000000f
R3[106] <= 640'h3808cfffffc0066f700fff7fe0003f4fffff00017fffe0001ffffe90077fc80400000f6800000030480080b8ffffff631fc000f738f2ffbe3c01f80c007f9e8c1ffffff818000087ffffcf10000031
R3[107] <= 640'h10dffffff4006cfb907ff77f080334fffffe003ffffe0000fffff9007ffcc00000107090000013001ec00927fffff771fc000e37137fefe3e83e00cc0331e000fffff7f00000087fffff800000031
R3[108] <= 640'h1033fffff057fcf9a07ff67fc00ffcfbbfff90087fffc0007fee09007de4800008007000000c0300fff009f3f9ffffe1fe00023e3178ffe3fc3e01801013000009f7ffe0010611e7ffff000000031
R3[109] <= 640'h817fffff017fefba8fff87ff1cdece13ffff001c7ffe8403f07c101fce6c0000c00000000000113fee0fbec3dfffff0fe0003fc3b29ff7f181e01080012000001f39fe1800613e7ffff800000030
R3[110] <= 640'h801cc1ff7fff8076fff697ff9fff1ffece23ff7f8108e7fccc01783f321f8ecc000001000200000001fcfce7bffffffffbe7fcc07bdeb2fcf77181e01000000000007ff97f380060dfffffff80000000
R3[111] <= 640'he0c68fdfc7ffa07ffff603ff9fffc33fd266fc7e8103c0fefe013c81361fc7c0000e2100b02000030beefcc19767ee777bf7fec3f1be833fff37c3e0000100080100fff9f8003974cfefffffc0000000
R3[112] <= 640'he3087799fff81ffe7fc873fe77f9bf2e026099b0602019f9d033198001fdf7c000671808c100c0037ef37c0cffbbfffcfc3de390cc423ff7ecfe0c00a010000800033fe3007f0e3f3cfffff08000003
R3[113] <= 640'h807ffffefbff03fff7fc87ffff7f9dfb60000001e6c0811ffc012098003fff608003f081fe810002f5bfffffdffff60fff83fff800cf60f7fffec3d1004000000000ffe4000fffdf3edfffff30800003
R3[114] <= 640'hf8cffcefbff03bffbff07f7fc7ebcff00000001ffc1803ffc187830303fe7400603fefbfff80c033cbffefffffb824dff07fff8001f0ef7ff7fc380004000000000cfc0013fff9ebefffecef0800001
R3[115] <= 640'h1cfe3fceffff0ffdf9ff07f3f8fffbbec00412c0fced00ffe0181026803ffec00f3fffffffec0f03bdbffffffffb006fcf07ffff830f0f37ffffc3800300000000001ec081ffffffcfffeee0f0000000
R3[116] <= 640'hf0fffff08fff9ffffbf807bff8cffffe80663ffc6f3f01ff60000006841ffc4900fbff7ff3e7cf00ff7fffe3fffe026f8fc3ffff0000e137ffffc3f40000016000003f80d9fffefff7fffef8ff00000c
R3[117] <= 640'hc3ffff700eff9ffffffc01bfff7fffff7866bfb80c1f01fe00000006840f3c0b0e99ff3ff367fefc3f37fff1fffc006f0bc0ffff003821b7fffff3e00001006001007f81dffffffb7fffffffff000004
R3[118] <= 640'h6ffff000eff1fffffff01bfff7ffffff83f13180cbf00fe000000030007fc020f89fefff107ffff1c0377ff9ff80c7c7e80ff1fc17b1bf6fffff3e60000180000003e87fffffffffffffffffc000000
R3[119] <= 640'h78fffc0086ff07ffffe1c1ff21f3ff7ff13f00790def00f6000080213007e0021e9f8eff8003fffffc027ffb9f718cbf4600001f803b98b7fff2f13ffc12010000007f0e5fffffffcfffffeff8400021
R3[120] <= 640'hfffffe20827fbffffffc809fc1f00ef1f81936181fff80fb00000000001fc7039f7fbeff81c077fffe80cf7163980039e642227fc83080bffffee0f83fcfc6380001390ffff9ffffffffffffff800300
R3[121] <= 640'hf6fffe00007f266dffe303bff8f0c2fff808f9c727ffc018000000000007e007bf23be3fc0807fffe0009fe1618080396e4208ffc81080bffffe70000bffefe00001f81ffffbffffffffffffff800000
R3[122] <= 640'hf3fffc02007b03cff3f301bffce10361f8016c7f57ff83fe800000000003e0073ff7be7ff8003fffc0181ff06080003c0e0148ffec00003ffffe38000183fff0003ff81fffff7fffffffffffff040000
R3[123] <= 640'h7fffe006807f07cff3ff003fe73f0000f0016f760300077f00010d0000037087ffff3fffe0000e7e80003ff04080c03c0e0d023fbc000133ffffe0000001fff8c17ff87ffff6feffffffffffff000000
R3[124] <= 640'heefc03068007007fcffe003fe63f800f1070bffe94c31ec000010800001f70ffffff3ff80000006600003ff00000003c06e8003f9f400001dfffc0000000fffe00ffe0fefb66ffffffffffffff300004
R3[125] <= 640'hfef838060007817fceff0837fe1c8000f8103031a0037fc0c0608000001bf03fffffcdb8000021c000183f000000813fc04c003817e000019f6f180083801f3fffffe0fff746efffffffffffff700000
R3[126] <= 640'h7ff0700c0000c3effff71836fa1e8300f8010980ff007fc0804018000011f807fec7cc11111ce106000c1f000000011fe00f400083e000339f7e003edfc0001fffff017f779fffffffffffffff700000
R3[127] <= 640'hf1000388d00003cffffb0006f9f9f8fe7c808970dfc383fc00040c00be01ec06fefeec16b11cc00680801c300000381ff0fc6000caefc033dffec37fffd1001fffff0967679fffffffdfffffff8e4001
R3[128] <= 640'h1866019cb00186ffffcec024388016919c430efc0ff981390000018038e7c04979e3c1073fff80618183000100009cf9b8c00027707165118367fbffff9d10037fd09b790efffffffc7effffffe00000
R3[129] <= 640'he100001f120125fffef0180000003641380e0fff007c8647040009004167c00df9f048839fff8020007f1860c0008fc1f100037ff87f6601937e1fffffdd010131c0039d07bfffffff7effffffc00000
R3[130] <= 640'h603fb00025fbfcf098800e0071e0000e01ff807e8607e80079200167d00fffe07c83cfff800000301801c8002f81790003fffc3bfc00123efff7ffdd01603000e3b803effffcfffffffffff00000
R3[131] <= 640'h77f08016fbffc00180060073ec84c600a781ff803ff88069601c6fc07fff00e903cfff800c00303907c0003e00fcc0037fffdbfcc01004fffbffdd904030007ff8f3ffeff8ffc3fffffff00080
R3[132] <= 640'h1000067be8006fc81800180000017bffcf6200061e0007f0f004fc03fffc073e00000e3ffffc01c002001ce48007e00f8e0fe3fffc0e2e60002237fc7ddd94000073fdff8ffe6fffe91fffffefc0000
R3[133] <= 640'h71c0001e3a0087fc0080000004018ffff97e7001e1e0c1ff3318efe6effbc0f3000083c033ffc11f0000018e4481c4007378fc3f7fc1003f8802213ec7008f4000073fff38ffffe77f39defffefc0000
R3[134] <= 640'h7f6003bcfa0087fe00000c000101effff97f79017d80fb1ef0b9fffefffb01b8300003001fffc11fe700810fed9b8000737be0d97f70601bc800600c04008f640064fffc9fff3bc00f301efffffc0000
R3[135] <= 640'h837fc0ffff609ff600008e0000007541f97c01007c430039f9b97ffeffff03383f0016000effc11fffe0df3fef038208f8e200c0f87ff7017c800c060800df76017ffffefffef910c3633bfffffc0000
R3[136] <= 640'h8787c1cfffc13f70100001000000f8000c7381013800011ffcffea37ff9c47e03e60010007c9813ffbf09d9fe7e68000f17e00f0e638bfe61e84240000003fc098917fffff9efe81390c3f7dfffe0000
R3[137] <= 640'hbefff1f33f7837f0800000000000f84080e0180179380003ffffee9fff987ff0306000010761893ff9ff0dbfffff000ef9180004f0001fbe1f8c000000013f039d1fe7ffff723c10180cf8fdfffe0000
R3[138] <= 640'h1effdff21ff97f58800300090666fee000001081f1b483427fff020ff890bdf8000000c3826308ffffff49bffffe000ffc18000cf000239f1cff9e7000007f1ffff9fffffff30000000100c9ffff8000
R3[139] <= 640'h9ffefebe3ff9ff988000000026ffbee700000001e13d9c6873ff011878001efc0201037fc06000fffffce93ffffc001f78f8000cf80024f81c3ffff000c0ff3ef6e3ffffff3b000000010349ffff8000
R3[140] <= 640'h97ffffb007397f184000800366fffe6608800041003fbc7d01ff113878040ef800001f7fc00101fffbffe93fffff00fefcfc0038c8000ef8800ffffc0003fffcf6c7f3fffffe000000000359ffff0000
R3[141] <= 640'hb7ff7b80033f7cc3c000003366fffff01c3000690087ffffc1ff01d1638017e00000feffc0096fdffb7fe13efff8c6feff7c0071c6000dc8003fefde0002fffcff3f5fffffc7000020000059bfff0000
R3[142] <= 640'hb77f668001fffce6c600001cfffffff01f3d804dc007ffbfe070608c03016fe00006feffc4827fdfffffed3f6ff8efffff7c003bc400980000fffffe0040c3ff3b7cfffffe870000000000499fff8000
R3[143] <= 640'h8275e61000fe7eeeee603004fffffffcc0f8008cfc079fff80f8601c3c0047e00006cefec4264bdfbfffbf3f67bf06d3fef0000f600062040d1f7ffc000783cfb967efff7ef00000000000019fffc000
R3[144] <= 640'h10ef6c0017e673e7ed840008ffffffe000011e799013efe807fe88c38813b0008016efcee03f886c6bfdffc1fff817f0e10c71bc000c0036167ff08800019039fff71ff9db0c3000001191c3cffe304
R3[145] <= 640'hfffdc016e677ff7f902001fffff7fe0000164819b36fc00ffc9c0e3003bc000030fffee9f80900ffffffdf1f9c0ffe77e4d1ec8068103767fff008000f831dfffe3ff9b8103006ec018008f7b7800
R3[146] <= 640'h7effc81fe1fdffffd07003fffff7ff800000c001f1379837f498043801bf000078bffffff80020e811fffc3fbffffe3ff1f7efc3f03fffefffffe00000930ffff77ffc38120017ff07c00077f7800
R3[147] <= 640'h2201ffff99f21bfffffd0c10037e8fe3ff00000820415370817f400100c813f00002d97fffbb80420080067d07ff7ff83ff9f6f8fc7981fffefefffc8000032079ff7ffef70070017fff76003fffe1e0
R3[148] <= 640'hefffdff381f1fbffcef8003802e1fc000180000353fc00ffe83000c013f80200fefffffb800000000008e6fff91f1ff937f9fe3fc0ff7ffefff8ec00000071fffffffe00008fffff7e800ffeffe0
R3[149] <= 640'hc5ffffffe03f139bf9effe0000031fc004080000213fc007f49f001c217180100fefeffff088c3e01000064f7790e8f49e201ff82c07f733cffe0fe80000079ffe3fffe4000dffffffe80c3fffee0
R3[150] <= 640'h26803fffff1c07f131bfbfffe0000001ff10cc04500037cc837fe8c103e43301410cfeffffff8c003ffb6000037370008045e0209fc100ffe31cffe7fec680007fffe7fff60003ffffffffc0033ffe40
R3[151] <= 640'h2e8429ffff866018e3bffffff00000831c71cc7c800035c0007fe80018e112ff4c08667effffd807fff9e00001706100186420609dff30f1e798dfe77fcf0000ffff3effe784e3feffff67e09c9ffe00
R3[152] <= 640'h3c6603f9ffcc980000fffffff800100e0fede17f0103cf30003fb93806c086fe81836ffd7f7ffc007fff7c6610701800e03380301f3ecc3ee067ffcffeffc00103e31ffff000ff99c78f3f80009ffffc
R3[153] <= 640'hff640339ffccb8000003fffffc800000077fe11f013effe0001f993843f803b9c038fffdf9fffe007ffff7001800000000b7000ec01f6ffff077ffffffff80003f613ffff000ff98ff9f0ff8002ffffc
R3[154] <= 640'hdf448019ffc07e000003bf3ffc009000077f39ffc03f77c0709ff93c63fe4b10ff7bbffefcfff7007fffffc0000001000096018c910427ff3ffffffffffe840018013fff10008ffeffbf8fd80033ffff
R3[155] <= 640'h1f88c0018340664000031ffff901f30007ef1dfdc4fd3c0978defd0c73cf64007fffbffeff79b9807f7f7f800121e0000002008c191803ff07fffefffffe008000313fffc4001feefffb9af80023ff7f
R3[156] <= 640'h1cd88080000066020000fdffffc0f3c00fefff7fffcc1c0079fe388f7fcf67400f7fbfbfff6df880736ffc00cffff8002003800e1a8c01ffffffff7fffff30c00001f8f3c4001ffefff39ffe000fffff
R3[157] <= 640'h1fdf3800000066028000fff6ffc0f3c00f7fffffbfc8078033ff3c8ff7fe7d7e01e3fe9f7eedf88003fdf9017fff9e000001000e80c000fffff01fffffff71800101feffc0001ffe7ff31fe6000fffff
R3[158] <= 640'hfffffc8101000783fe801ffeff81f2e0077ffff03fc10780637ffffeff7fff7f6601bac77efff88007ffd8017f8f8fc000006000c00381fffff01ffffffff9000001ffff00000fff3ff31fe60003ffff
R3[159] <= 640'hbfb0f43900000f8bfe0001e77ee1f6e000afffe03be90018e17efffeffe7ff7fe0009046ce8140800f4fdc49dc878c78000dc60f6179837fff76007f7fffff0000031ffc3000e7db7ffb07fe0001ffff
R3[160] <= 640'h1ef8c77680801983fe00007bef70df7836ffff67feffb188c7e8d9fbf867f3fbd9c00103f8c0e1039f3e7207080006fe780f8001533fc1f3df800000181fff9c008119c60081fff3fffebfff001bfeff
R3[161] <= 640'hc7f84ce2c3001183ff400f7dff98df78027fffffffff0008004f1fff996ffeffc9c00000ff03e0f09f8f70060200063f3906000040fcc0fffc0000000001ff980000911c00007fffffe4bffff011ffff
R3[162] <= 640'hc7f86c8293000083ff4000fcffb8f3f8027fff7f7ffef028006d7fffc16dfeffcbce0100030080f0fecffc0fc000037f7f0400068c3e41fff80320680000ffc10000811c0001fffffff69ffe0001ffff
R3[163] <= 640'hffbf7cb039800001ff00008099f0f3f893fffffffffe7f2007e87fffc0e1ffffffff00000000017fffeffe8fe90003fbf380c046810f017ef18fe0fcc400ffef800000c00001ff7ffeff8ffe0000ffff
R3[164] <= 640'h7e8ffdb071800000ff40038019b3fff893ffffffffff07a206492fff00e1feeffffe0080008003fb67fffe83ff7003ef66c0006601c0087fe70fe36cce00ffffc00000c30000ffffffff9f9fe000ffff
R3[165] <= 640'hf7c1fd90e39900003fe400000fbefef9107effc77fff028000417ff3041ddffffffc8380068003ff677ffe09fffc030fdfe01866808000831c03ff6f06007ffe8000c71000bfffffffd93fff0000ffff
R3[166] <= 640'he7fbdd92df9980223ffe0400677ffff9007cfe872ffc60880040fff7063dc7ff7fffc3000e00007ffbfbfff8923fffffff600070e680b0011003ffefe70003fff1000000003fffffffd97f7f0f00ffff
R3[167] <= 640'h77fffd1e1cd08003fffc8000667fbdf902e3fc040f3c248800819fe6e0c933ff7ffff820004207fffb79ffe11a33ff7f7f2403391ece3e80000fffbbf7f003bff8000100017ffffffff9e2ff8001ffff
R3[168] <= 640'hbeffffc1c7667003ffe2800003ffffffc10183040080000c0001ffe748c007fffe77c18330401bfebfffff7f0100327fee00467bfff37fe0003365fff7801cf3ff0e000007ffffffefefffe3c003fffc
R3[169] <= 640'h93ffffc6dffe1c0c9ffe0000f0fffffec00080810000c00c00003ffecf807cffff3c489070851ffefffffffe601810414c000cffffffffff803bf77ff6c00cf3fff800000fffffffefffffff0803ffff
R3[170] <= 640'he7ffffce7ff8cedefffe900010dfefffc10100000030004c0006fffecf800efffb7ec89800681ffffffffffefc7800184c0018fefeffe0ffff3f7f7fbee001fffff0068effffffffeffffffe0801ffff
R3[171] <= 640'h774fffee7ff9deffffffc00001c7efffc60000000010014c0007f3e7edf807fefcf7811f00689cbffcfffefffe1f6d80000039fe0ee70003fffffefffff0011ffff307cfffffffffeffffffcc000ffff
R3[172] <= 640'h5e4fff63fffffffffeffc3400007ffffd02480000000007c2003ffe7fdf8dfffcee28118910d1fbfeffffeffff8f7fe1900033fd03ee0000ffff7ffbfff1000ffff30f7fffffffffeffffff8c000fffc
R3[173] <= 640'hf2fff363ffffff7fffdffc000007fffff8c680000f00017c20037f3c78c01fffdf3c02011e0707bffffffffffecfffffba0067f103e80000bfffdff17ff300007fffffffffffffffcdfffff33001ffff
R3[174] <= 640'hb3fdf720fffffefffffffe000007fbfffc63800019800968300fff7e79c0dffffc3e02c74744c6fffdfffdfffcffbef7fa0067f9000080003fff3ffffffb00003fffffffffffffff4dffffff30017fff
R3[175] <= 640'h9f79ff3c7fffffffefffffe1000771ff90a0081cf0809841fc0effff7fc69ffcf0025000934c06f77ffffdfe3c3dbe7f7e0066f8000080001dc77ffffffb00003fffff9bffffffff49cffefc03307fff
R3[176] <= 640'hfd7be7773efffffffffbff9880030ffff902080cc000001db80ffffe3f7d3fe4600400004d7cdfff7ffefffc98c3ff3fff7007f10881000387fffefedf7ff8003edeb946fffffff030effff4810407f9
R3[177] <= 640'hbf79fc7667fff9fbffffff980001063ff80080071f300609f807fffefb690fe4400200404dff9ffffffffffe9873ffffff6063f00800003fff7fff8fdf7ff800273f00007fffffe0004dff7e0806c7ff
R3[178] <= 640'h3f7838e6e3ffffffffcee7fc000000fffc0081113cf002c1c007fffff14186e0000000000fffffffe7ff7ffe801ffffffc0063f80800003fffffff87ffffff18033100003fffffc3806fff7e0000ffff
R3[179] <= 640'hb88000c622ffdfffffceffe7000000ffff013980fcf700e1c01ffffff340cf70000000181f7fffffeffffffe0007ffffff0063ffcc0003ffffffffe0ffffff18000000001f7fff80000dfffe80007fb6
R3[180] <= 640'hd180008f20f3fc9ffff33f7f0400000eff0039f08fff103e803ffff8ffccf370000100091ffffffffffffffc06e1fffffb00039fcc0007ffffdffff07ffffef000000044067fff000000fffec0073ff7
R3[181] <= 640'h8380388fe3f3ff8ffff3fdfff800000eff0003b91bfe80390003ffffffcc7171000000006dfffffffffffffc1c18bffef000019fbce30f7ffecffff3fffffce00001f166007fff300008ff6eb80383ff
R3[182] <= 640'hd9000019e3fffffffef3f9fff0810007fe83033c3ffe80488003ff9fff4800000020018049ffffffffff3fff8007bffe2000001fbdf6cffffee7ff7bfffffcff0effffff001bfec0006d78069000c3f8
R3[183] <= 640'hf838033938fff97ffecc9fffe7c00007fc801ff07fbf8101c090fdfffe610000a00004010ff8feffffffffff80e1bfc700600c0e9f7efffef9713973ffffee7e7effff1f301bfe800000780081083eff
R3[184] <= 640'he601008446ffffff7eb2f9ffff820003ff1807716ffff003780177f99f843080108000300dce7ffffffd768c80009f980098070fffffff66ffcf7f677effe37fffff989fc418fef80001008400209bff
R3[185] <= 640'h1c00fffefffeb21fffffd00303b60002f07f7fffc008017fffb90000030100000083fffffffffd674c80000fc0001801ce3ffffce0800077e7ffffc0ffffff0003fc00ffa0001800000022bfff
R3[186] <= 640'h100000c00fffffffe96fffffffc0713ff0002f0fefeff800c00feff300000010130004003fffffffffdc70181101180013f008e3ffffc80000423e7ffff80fff3008080e6001f800000000000273fff
R3[187] <= 640'h100008100fffffffe96ff7fffe6c011ff060233fe00ffc00004fee6000000000020016000f9ffffffffd8010100390101ff0007bfff1018000c017eff3f03ffe10002803fc00fc00000000000073fff
R3[188] <= 640'h1ffffffe97ffffffe6c0016c060013fa03fff8404c1fee00c4000300010344803ffdffff6d1c018000300000ff780007ffe0180000003efefc077fe10007901cf007f00000180000039fff
R3[189] <= 640'h1ffffffeb3ffffffff9800dcc20003f2c3fff0800f9fec010e0087b00180c6193ff9fff94900008000000000f7fe0003f3e0000000000b7cf80f77f3180318007e07fc00000000000bffff
R3[190] <= 640'he000000021ffc9fceb3fcffffff9800dfe3040772f8fffb900df9f800000038000080fe98fffffff948400000000001007ffe0003f000000000008166300fffff7c3000037f07fc80000000021bffff
R3[191] <= 640'he10080006703bf9f4ef33f9f7ffa9100193c4c6420193ef19108db310c18983b010c0f39c83feffff1401a0000000080013ffec10000038080000018c7000fffff7c000023ff86fec0810000003fffff
R3[192] <= 640'hf00606001f03c64c6dfe9fff7cffc08c0effe13e00032eff7c193ff80f310008f803e7fff08ff77ff8c8002008020080be7fe68000600000861800000c00037fffff9000013f8ff781003000000ee7f9
R3[193] <= 640'hf07e87001f8006cfe7ce9ffcffffc48c0e3ffffe001c0fffe67fe70008000000100307cff80077fffe0800000000000023ff7f98080180000001300000000037fffe000063ff00ff19000100001efff9
R3[194] <= 640'hb237c7ffffc00241e7effb3fdfff87180cbdfffc001cc67fe7ffe7000000040011001be77c017f7fe602708c10080003e7ce1ffc0e0b71000000180000000007ffff9001e7fe03ff3c000000001ffff9
R3[195] <= 640'hb023e7fffff8000007ffff1f3fffe00089f9fffc001ecfffffe6fe3010000000310b19fffc806ffde603f888be4c0033ffc01ffc07dd3180000001000000008633ffb207fffe077ff000c00000c7fff9
R3[196] <= 640'ha0fffffffff800081ffffefee7fff00009fc3e9e00871efffffffe800000000001033bffff004dc6603efe8fbffc003ff3c08ffe00dd870040308300000000060ffff28fffee01dfc32000000307fff9
R3[197] <= 640'hb2dffffffff180020ffffecfff7ff3c0033c3cc100c73bffffffef880000000000033fffff199cc6213ffffffffe803ffcc001ff00cdce980021000e0400000686ffffffffe403fffe200000033ffff9
R3[198] <= 640'hf7bf9ff803ff88be60ffffdf7e7ff3c0032000c000c7f9ffffffff000000000000097fffff9d8c0402bd7ffffdbf807f7c80007fc067fffc0000000c00000006003fffffff6007fffe60c080003ffffc
R3[199] <= 640'hfdfe1ffc03f38f9f70fff7fefe7ef0fca2e00000013f8fffff7ffe90110101000019ffffffdcb02066ff0cc761bf81ffe2000067c07c3ffe00040c1c0380000021cf7fffff60019f4fe200000023fefc
R3[200] <= 640'hfc3d01e0003ff7eff0cffefff99ffbc01dfe81800063ffffbebeffe0011300000001ffffff5f70010ffc0000801fe3fc30008019e01f9f7f103166890000200000ffffff8f8041fff360e2000407fffe
R3[201] <= 640'hf8000060003fffeff81f3ffff9191f808f000100000fffffbf9fffd88100000000e3ffffffffe001bff800000017f7f800006000f8199fff303f06888000000000233f60c000497fff606400000efff7
R3[202] <= 640'hc03a3c00000e7f00fc1cffff380007008fc00000809edfffff97ff9c8886000003eff7ffffff270fffc03c080003fff0000378013c001e7fc0fb60408000000000077c000000090ffff06600016efff3
R3[203] <= 640'h73fe0020004100fe8cf0ff006087001fe0000000feff7ffb92fffe00000000037ffffffff9be0fff817efe8001ffc0000fffe81f803666c4f0e46400000000003ff800000349ffff81c3c001fefffe
R3[204] <= 640'he7fc00700040003fc607f3000080001fc08000c03ffffffab2dfff00100000033ffffff8f1fafbf003ffff82007e00001fff8f1fe0020080060f4080000000007b0700e00048ffff99e700c01fffff
R3[205] <= 640'hfffdf2708002787f660fc000000000cfc38080807fffffff369fff31230000837fe7f1c8007ff90007ffff83c03e00003ffff81ffc004000ccc000000000000030030040034dbfff7cff00c01fff7f
R3[206] <= 640'h3fdfffffff017fc7fc0000011000000e7ef808000ffffc17f36dffff903000003ffe370000026f000bfffffffc00003feffff7807ff400000c0c0000c4000000032f0000307491fff7cfc80601fff77
R3[207] <= 640'h7ffc7fdffff88fee3bc000001be604017fe0810e00df7f387e328ffff800000303fe38700001006403ffcfffffdc8007fffff7ff03ffc48000000000cc60f000003f3ff10000c9fbffe7f9c0e0099fff
R3[208] <= 640'hfff97ff0dfff3ffc3bfc0000390f660efffc786707ffff30cff0813ce01000261fff70204000d8020ff9ff00ffff807fff7e00ffc0ffc04030181607787c0000010373e20004c1c0fefefee93c003cff
R3[209] <= 640'hffffff03ce3ffffe1bfe00003fff7efe3f7f802006ff7ef08f9f987ff6800007ffff9000000084028ff0000080ffc07f0100003fc0fffe60601f90037e383c8170017776000018007ffffffd3d0003ff
R3[210] <= 640'hffffe401001fffff83ff01c17fffffffffff026001ff78000fdfd8fff08800c3ffef88000064bccfce0020000007fcff00000019f831fe38c2f9c003ff7ffcc33398773e00000c007ffffff9680003ff
R3[211] <= 640'hffffe1000008fdff83ffa1e3ffff77ff7eff060089fce000077f7bff800080f9ffc480001067dffffc0400000003fffe00008001fc00ff99c6fffcfffffffffe3f7cf77400000101ffffffd72000003f
R3[212] <= 640'hfffee1030000003f8187ffffffff2480f8ff00000e7dc00300ff7fff00010fbfff800000003ffffffc00000e000010fc083ef8001e811f9fdf3efffc1dc41cfff83fffe2000001007efffffa9100181f
R3[213] <= 640'hfffe7803f800001fc087fffffffc100178ff40009eff000000fefffe00481fffffd80000003fffffc00001280e80010008fffc4007f81f4ffff69ff80000003effffffe7888080000e3f7ff88c000007
R3[214] <= 640'hfff7fc23fe80000ff0007f7fe000000000ffe000fff001fce800ffcc20183fff0f80008c00fbffffc00000e0ffd800001fffffff00fc0efffe6603c000000004ffffffffb9800000007e7ffda6800000
R3[215] <= 640'hfff7cc3fffc3e00478003c18c0010680000f44277ec000bef80018c020093bff838020dc81fb9f7380080e037ffc00019fffffffc01f0008c62001012ee00001077ffffef900208000c3f3ed0e800000
R3[216] <= 640'hfefce03fe7e3ff017c80000061038ff00013c176fe00137fff2100011fe17fff3000067ff0ffef0000031efffffee00ffff3fffff00fc00000001803e0e1ff3019f73ffffcffc8000420243bd31700d0
R3[217] <= 640'hffe7f8ffe33f7f60ffc68000197ffff8800fcf7fcc00bfffff6100011f78ffdf000006fff1fff80000030efffffff03fffe0fffff00dfcc00000d80fffffffc00100fefffffffe80000000c50f160008
R3[218] <= 640'hc1ffc3fee3f83fc00fffc00f7efffff8c007cffd0000fffffffe0011ff7cff8f00062ffffffc380000011fffffffffffffe007ffff017ef3ffffffffffff7ffe000078ffffffff80080000f42c9f84da
R3[219] <= 640'hc07f83fc00e007c003fff8bffffffffcc003ff780007f0f1fffff8bfffffffe0000e7fffffff300000005ffffffffffffff007ffff1007ffffffffffffff3cfe0000043fffffff98003000110a178448
R3[220] <= 640'h603ff000303c0007ffdffffffdfff0003bf480107fc6007ffffffffffffc0031e7fffffff7100001efffffffdfffffffc037ffeb203fffffffffcfbffc01f0000037ffffffff1737000407e17c85c
R3[221] <= 640'h383f7000103cb001ffffffff8c7ff6003fec103ffdc0207ffffffffffff00c3fc7ffffffbe01f00fffffffff9fffffff803fffeb0c13fffffdbf8ff87801ed00001e73fffffe57ff080317557fcf8
R3[222] <= 640'h47eff7000001dffc006ffefff0007fe003b01007ff880403f3fff98eff7c007b3efffffff8e01fffffffffff187ffbfff000ffffb0c00f07ff99707801001ef800006333c3fff57fe6bf5365d1fca2
R3[223] <= 640'h7bf3f000c000ffff0007fe0771713fe000330307f9c0003963fc10047e00013f3e7ffffffc003efffffffffe183f71fef800ff3fb8380000ff980010000083fd8000380018f7b81e6fff2ca3d73978
R3[224] <= 640'h207ff400000c033cffe0008800f861fffc00000ffffc00000000000000060000fff6fffffff0113c7ffffffff0fcdff0c1c000037ffec00000010000000000007f80000400004f7edaedb7b4fdcabff5
R3[225] <= 640'h3ffe000018c0100fff00000000021fffe00007ffffe00000000000000040003fffefffffffc81fcfffffffffa3fff6040000003ffffe00000000000000000003f80000000004f2e1f1fbfaaf44329fe
R3[226] <= 640'hfbfc000003dc0000f0ff0000000000ffff0000ffffe0000000000000000001fffffff3ffff3801fffffffffffd3fc40000000001fffff80000000000000000001fc4000000004a4212ffff661701af7e
R3[227] <= 640'hf9e0000103fe0000001fe0000000007ffe0007feffc03c3c00000000000001ffffffe77cfc1803ffffffffffff5fc000000000018ffffc000000000000008c000ff8c000000001394525deb0b490de1b
R3[228] <= 640'hfdc000030fff0000001ff0800000001ffe001ff0fc003efe00000018700009ffffffff3c800003ffffffffffdfe007200000000087fffc21000000003ab38e0007fce880000011f66c45143621ff433a
R3[229] <= 640'he7c000061fff0002001ffe800000001ffe007fe00000ffffc00c0010f8639fffffff3e0000000dffffffffff87f00f000000000107fffe3133000081fffffffe03ffff80000000f9b41015224db6655f
R3[230] <= 640'hc1c00006ffff800300007f8cc0000007ff81ffc0000fffffffde87e0e3e3fffffeff000000001dffffff7fff07f88400000000011ffffe73fb301fffffffffff80fffff9f8220173e1831014deac06ea
R3[231] <= 640'h106ffffc01e8e001f8fff810007ff8fffc0001fffffffffffffc77efffffeb9800000004dffffff7ff3077cc000000000031fffffffff383fffffffffffe00fffffff6601f3820c08d7e5c96877
R3[232] <= 640'h800101fffffeff9f000fceffe000039fcff880007fffffffffffffffffffffcffc000000000ffffff303ffe6980000000000001ffffffffefc3ffffffffffffc01ffffffcf651c7b39cf79191f2955
R3[233] <= 640'h1e3ffffff1fff0007fffff3800007ffe003c7ffffffffffffffffffffffdffc000000021ffffffc03ffe6800000000000001fffffffffffffffffffff0ffe0003fffffe47c59172bf2547915be9
R3[234] <= 640'h63ffffe30fff0000ffffffefe0017dc003fffeffffffffffffffffe7fffefe000000039ffffefc07fffe810000000000001fffffffffffffffffffff03ff0000c35fffc12a8ce5b12e85b9dbef
R3[235] <= 640'hc0000003ffffe3ffff80001ffffffff0000c8007fffefff3ff7fffffffffc3ff100000000003fffffefe03fffec10000000000001ffffffffffffffe877f3c01f7fe00011fff4a21f3c677762137db2e
R3[236] <= 640'h38000003fffffffffe800007fefffff0801c00fffffcf800033fffc0ffff03ff000000000003ffffffff013fe1c18000000000000ffffffffffffffec31f0403c7fc0000071d555a9b0062c48679dafd
R3[237] <= 640'h380400f07efffffcf8800006fcfffff880080efffffff800001ce0003fff0000000000000803ffffffff011fc1c9c000000000001fffffffffffffffe063000003ff0000009b457cb14ba30a1f01857b
R3[238] <= 640'h380c00003ffffff0f8000006981ffffcc0000ffffffffe00000000000fe10000000000000003ffffffffe3ff99f9e000000000011fffffffffffffcf7c00000401fff3000002a94f55f80008a64136ab
R3[239] <= 640'hfc0800001ffffffff00000000707dfff60200fdffff7ff00000000003fe000000000003c0101ff7f7f7effff98f8e000000080001fffffffffffffc77e00000200ffff180012f982f4b3ee296db13cf5
R3[240] <= 640'hc3380000803fffc01c6000000c03ffff8c310ffffffff000000000007f00000000000082603cffffffff703e7dff7c00000000010ffffffffffffffeff000003e51ffea82a1985cd23b25c31a931367d
R3[241] <= 640'h1f000000c0000c1000000000000fff7fe731fffffe1e000000000027f0000000000008f607ffffffffe316173fffc0000000000dffffffffffffffdf0000003241fff2fbaab3686ca9b92d3e40a8c9a
R3[242] <= 640'h80000800000000000000503ffffffffffc04000000000803c0000800000838f62fffffffffe7fe3d3fffe000000000017fffffffffffff9e0000000064dbcaffb9aa084f2e7d2d2b5efa416
R3[243] <= 640'hc0000180000000000000001ffffffffffc06000000000f8003e71fc0002c7df7ffffffffff6ffeff1dfff0000000000e7fffffffffffff9c0000000044cbc3ebd489eced1e082cd188f6258
R3[244] <= 640'h100781c00000000000000003f7ffffc7bc0000000000138007fffffc18fffffffffffffff63ff1ff85ffff00010000087fffffffffffff9e0000000044c27e7ec57e234eccd6763f2e58e94
R3[245] <= 640'h1007c8300010000000000001e73fe8039c000000000013e03ffffffe3cf7ffffffeffffff73fc0efc1ffffc00000000c7ffffe1fffffffec0000000023c2297eecf22a01e741ac14b66be02
R3[246] <= 640'h7fc100010000000000000c010000008000000000007e07ffffffffcf7ffffffffffff863fc0cfc1fffffc00000f183ffffffffff87fc00000000053c385fde8b3c565e2eecfc657e3735
R3[247] <= 640'hc0002003fff80000c00200000000040000000c800000c63800fe0ffffffffee7f7ff6ffffffff877fe80e31fffffc00001ffc3fffffffcff87fc00000001453c244a1cbadf1557b89d034c2cc5f3
R3[248] <= 640'h270008018c3f80000001e03c8000000000000000000fff3f801ff7fffffffffffffffffffffffffdeff0077ffffff8000037ff0ffffffffc0fff8c300000037adf4865fc09dd6b7293f17bd7a5e62
R3[249] <= 640'he0003fc8000001f8ffef00000000000000003fffffc03ffffffffffffffff7fbfffffffffffff007fffffff000000f1f07ffffff0c0fff07e000081344606c39ee47ffe54a88485b2a21b24
R3[250] <= 640'hc00000003fc107fffc00781fffffff00c20000000006bffffffcfffffffffffffffffbd61fffffffffffff8003ffffff00000043f03fffffc03dfff03c000000d69156533fce31cd6c11b14d8f3af69c
R3[251] <= 640'hf00000007febfffffefff81fffffff80c3800000003ffffffffffffeffffffff7ffff3c21fff1fffc77ffe4001ffe3fe000000031f3fffffe01dfdf018000001ad0f7aa65f393828131b90359e45d91d
R3[252] <= 640'hf00000003bfffffffffffeffffffffe1ff00000ef0fffffffffffffc7fffffff40ffecc3bfc003df01033e0000ff807c000000031f3ffffef3fffc000000005d25934064561784b632028493a1704b1f
R3[253] <= 640'h803bffffffffffffffffffffffff00003ff7ffffffffffffcc7ffffffc003c00421000038e01001e0030ffc13000000000073ffc7e3ffff00000000054b5259a085be79daf541c5bb8c3b8fd7d
R3[254] <= 640'h13ffffffffffffffff01ffffc000c3f73ffffffffffff8cfffffffc401c00060000000407800e0010000000000000000201f4dc7fff400000000030f26770a41a54fcdec9af9361a7d36b8a
R3[255] <= 640'h1000000000ffffffffffffffe010ffffc1c0e3ff3ffffffffffff8edffffffdc01c000c0000100c1d0007f80000000000000080000007fc3ffc000000000029f5e859db711f8f66b83f955e1a70b41f
R3[256] <= 640'h8000000000033f7fffffffffff0117fffc000038c3ffffff7fffff86cffffff1c00000000000000000809c0000010080000000c008003bfe3ffc0000000000936b3f4b3914d5b26a602e10b2d207e103
R3[257] <= 640'h7c000000001b133ffffffffffe0103bffe00007fe3fffffffffffe8407ffffe0e00000000000000000003c0000000100000000c000000ffe000000000000006b6a7dcf3d4d03f48106814b7c086651af
R3[258] <= 640'h3c030000001e03e7fffffff9f80002003f0000fffb9ffffffffffcce07ffffe030040000000000000001700000000100c000008000000e0000000000000320cdbc735aae3088be95ba4a58d7e6a57b3d
R3[259] <= 640'h80000060087ffffffff7ff8e00000001ff03efffffffe7ffffffc8407ff01c000000000000000000000e1000000300002000080000006500000000000003077569bee8ab6623991983a947892522283
R3[260] <= 640'he07087fffff03f01c0fc00c00003f3fffffffffc3fffffff001fff470080010000000000000000000000003820030060000000055000000000000000443f587f26070027e4938ee1b15ab2cf06
R3[261] <= 640'hc00c7fc0c03fff03e0000fc00c00000fffffffffffc1f3fffff003fff1d0080000000000000000000100002007ff303007880000000000400000000000025cbdfd70ccb1e95e6cbb0a42aeb568942
R3[262] <= 640'he001ffe08013fff1e00001c00000000fffffffdfffc3f3fffff0070ff640080000000000000000000c3000a0fffffff83fff80000000008000000000001df9c3e8e81efc42e9b123ff52ef17c6f1c
R3[263] <= 640'he000007effc00103fff700001c00000001e7fffffc7fe03e87ffff80181701c0000000000000000000007000183ffffffffffffe3f800000000000000000c2bd954bd70f99d84fd6acbb272b99458a31
R3[264] <= 640'hfffffc00003ff0000000020000007ffffffefffc7dfffffe101f031f0000008000000000000000c000000fffffffffffffffe00000010000000000a6b01d28a81dc5f21871764fd01f7dffa97d
R3[265] <= 640'h60ffffffc000ffe0000100000000003ffffffffffdff7ffffe103f8140000000000000000000000040000007fffffeffffffffff000000000300000077a31efbc3913f2fbac6d270ec61f273414c
R3[266] <= 640'hc0ffffff03fc3ffff00ff5800040000007fffffefffffe7fffff787f80000000000000000000003fe0000000001fffffffffffffff800140fac7e0800100c7cbd2f37763946d312c8f41861308df49
R3[267] <= 640'h3fffffffc17ffffffffff9000000000005ffffffff3fce3ffffff0ffc1c000000000000000000fffff0000003f3ffe8fffffffffff000068ff03a000015e42f9c6a9fc6efa2f7dedec933ee294ae69
R3[268] <= 640'hc01fffff000ffffffffffe700000000000013cffffff3fc41fffffffffe1c000000000000000003fffffc0e0037ffffc8fffffffffff00000af80000080149a56c564417523a4a58daafbc5585076086
R3[269] <= 640'hc00fffff001ffffffffff0000000000000000000ffff01801fffffffffc00000000000000000003fbffdfffff73ffffc3fffffffffff000003301c00c1000d6bd9eea3496f5b62e0d5796167cc19780a
R3[270] <= 640'hffffc031fe0ffffc0000000000000000000007fff20001ffffff7e3000000000000000000003f07ffffffff3ffffe3fffffffffffffe800200000c008dbb797e279de0bc7fb730e218e6f2deb46f2
R3[271] <= 640'h3ff87fffc0ffffc0000000008000000000007ffff0003ffffff7c1000000000000000000033f00e1fffffe1fffffffffffffffffffe800fa003c0c00984e857cfd06be1f5744791eebdb78e89291
R3[272] <= 640'h7ffcffffec7fffff80000c000000000000004fffff0000ffffff800007c00000000000000001f00ffffbfff1fedfffffffffffffffa000000000000c0ff6da59890967c21f91d1daa7a937be75b3e
R3[273] <= 640'h3ffffff3900fffff0fc000000000000000000fffff8060ffffff800001800000000000000003e00ffff1ffffff9fffffffffffffff800000000000200bf371e2fdf63b7bfe6f92392659f07aba50b
R3[274] <= 640'hfffffe0108ff7c00600000000000000000001ffffc071ffffff800000000000000000000007e00fffffffffcfffffffffffffffff80000000001f070dd77e83151fb2bfc6a15b2ec396c0041bf4e
R3[275] <= 640'h1fffff8387ec11c00000000000000000000000fff7fcfff7ffffc0000000000000000000003ff00fffffffffffffffffffffffffffcf000000000ff630d7b77a2b3b2c7ff439653590eb9450dc9f8
R3[276] <= 640'h1007fffffffc7e8003000000000000000000000003ff3ffffffffffc0000080000000000000007ff3fffffffffffffffffffffffffffffff80000000ff63f7f96bdb7c3998e37f2e2adf8fb0cabed7f7
R3[277] <= 640'h3cfffffffff8000003100000000000000000000001fb3fffffffffff00003c000000000000000fffffffffffffffffffffffffffffffffffe00000000f07393ddcf5c569f25bb2c222d9eac7ed8abf0f
R3[278] <= 640'hfffffffffff0000001000000000000000000000000711fffffffffff18003c000000000000001fffffffffffffffffffffffffffffffffffe0000007401ffae076f62ba7fde1f1eeab569bc5e7de2b6c
R3[279] <= 640'hffffffff0000810000000000000000000000000000200efbffffffff180078000000000000001ffffffffffffffffffffffffffffffffffff0000007003f98de2da2dae15d3cdd1ad3cb329b95708b64
R3[280] <= 640'hffffffff8000000000000000000000000000000001c0077ffffffffef80000800000000000001fff1ffffffffffffffffffffffffffffffffe00ff07ccd55e98226db2fce7d72eb7f718b347afbd7326
R3[281] <= 640'hffffffff800000000000000000000000000000000100017ffffffffcf8c000000000000000001fff3ffffffffffffffffffffffffffffffffe00ff0fcc5df2d323904aef972a5ce9506b8dd1a1fc0e11
R3[282] <= 640'hffffffff800000000000000000000000000000000000007ffffffffcf0e000000000000000001fff7fffffffffffffffffffffffffffffffff00ff1ff04cf6fb57e2ca8f5bdcf17b795fd567fca2ce43
R3[283] <= 640'hffffffff800000000000000000000000000000000000007ffffffffce0f800000000000000001ffffffffffffffffffcfffffffffffffffffff0ff7f70effbeddf0c92c9fde6bbf2a9be6a90dceafd28
R3[284] <= 640'hfff77fffc08000080000000000000000000000000000007ffffffff8c0ff00000000000000001ffffffffffffffffffefffffffffffffffffffcfffff07dd80f3a698f01e1bbf0b2f1cef5be5b81da66
R3[285] <= 640'hfff33fffc00000080000000000000000000000000000007ffffffff800ff00000000000000001ffffffffffffff7fffffffffffffffffffffffefffff04ca3a69363f6bc1b74ff0eaee73ef5b623d1ee
R3[286] <= 640'hff000fffc00000080000000000000000000000000000007ffffffffc000700000000000000001ffffffffffffff7fffffffffffffffffffffffeffffe87ddfcd3789be4ea531fbf4c340faa8131aff30
R3[287] <= 640'h10000f7fc00000000000000000000000000000080000007fff7ffffc0000e0c00000000000001fffffffffffffffffffffffffffffffffffffffffffcc374fa79f674efaae399fc937edba8bbd07d2a9
R3[288] <= 640'h77fe00000000000000000000000000000000000003ffffefff8f80000000000000000181ffffffdffffffffffffffffffffffffffffffffffff8c6e77dd8f9bd7edfedeb727426bf73f1a0d20ab
R3[289] <= 640'h7ffc00000000000000000000000000000000000003fff1fffffe000000000000000003c7ffffff1ffffffffffffffffffffffffffffffffffff837772febe4f6752dff3dfbedbd39d4f3b345106
R3[290] <= 640'h800000000000000000000000000000000000003ffff0ff3e000000000000000000ffffffffffffffffffffffffffffffffffffffffffffff23bf3cdf4ff68eb57b1131dce1ae5a4e25bdea59
R3[291] <= 640'h1000003ffff00f3c0000000000000007ffffffffffffffffffffffffffffffffffffffffffffffff23fd9c7adca07c1e077fdea56a513fd72b1cb775
R3[292] <= 640'h1800003f7f310030000000000001000fffc3fffffffffffffffeffffffffffffffffffe3fffffffe396eed82ef8178915efec96194b1f14f4ea59226
R3[293] <= 640'h3003f3ff000000000000000000007ffc3fffffffffffffffffffffffffffffffff8a0ffffffc0ccf26c5cf1479efa7e8b1f8def63497d7f6357d1
R3[294] <= 640'hf003f1ff080000000000000000000ff817ffffffffffffffbfffffffffffffffff8001ffff800c07ebe3794d866f9fdeeecfa92f60fae0b86638f
R3[295] <= 640'h33e003f038ee0000000000000380000ff001ffffffffffffff3fffffffffffffffffb080fffea00c1adb1697254e308cdc77fbd99068fdff0e39890
R3[296] <= 640'h17e00000f8ce00000000100800cf800e001ffffffffffffffffffffffffffffffff87831ebea080707ddde1b0841aff33f3eee7dafea9cffa77b5df
R3[297] <= 640'h3e0000078cc00000000c0000c7f000f80fffffffffffffffffffffffffffffffffc73eb2b2c08000fdc2b1d9a7836c53cf7bedc8df5d07bb5d6fc6
R3[298] <= 640'h1e00000100000000000c000c00f01fffffff3fffffffffffffffffffffffffffff8070e2328000806e79fe16048e05a1d65eeed2ef9ebdd4e4fd1e
R3[299] <= 640'h6000000000000000051001c3fff3ffffffffffffffefefffffffffffffffffff080e922120000c35faa61feb5a74d7b7bfa63d6e1af57af325dc8
R3[300] <= 640'h300002000000000000000000008033ffffffffffffffffbef8ffffffffffffffffffe000f93782000001afdd83f6073542de57bbf622cf6e18ea7ec55b
R3[301] <= 640'h38000000000000000000000be043e0ffffffffffffffe1ffe3ffffffffffffffffff80003f1282000000d2699eb24770cbc92f43d133a4f97b3954dc4b
R3[302] <= 640'h380000000000000000000007c06e9ffffffffffffffff3ffffffffffffffffffffff0000b750800000003ff99e15b2ea9b7a393e4922469b13f4f9ff26
R3[303] <= 640'h18000000000000000000003f487f561ffffffffffffff07ebfffffffffffffff01ff000179612d00c0001bd45e48fed1e8c4f7ed820026cb569fd1f6bf
R3[304] <= 640'h7ffc0000000000000000006c2c1c9791efdffffcffffff803fbfffffefffffffd869df881320e957dc025febb9df84de3a369feffcec3d7a2daaff2212d
R3[305] <= 640'h1ffe00000000000000001875dc625ca073efffffffffffc3c01ffffff9fffffffbe8fe700d2994bfffde43f2a23ad5adf3725cc5a40e123fd1043fe562b
R3[306] <= 640'hffe00000000000000007bd1656dce603fcffffffffffe03afbffffffffffffffbfff43fe9d154d45ffffcc275a341351dd6739deb143bd4c252ffdc8f4
R3[307] <= 640'hf00000000000000066717d90487800f8fffffffffff001ffff3ffffffffffffffffff734eb5d2ff037fdec6cf81fd0e1ae09596b7af7c73467daac75
R3[308] <= 640'h1f03ffff00000000000000587649fe43d1000107fffffffff8ff1fffffff3ffffffff0c0fee690e9717fff77b409ae8a0358253f2a9fcb32f6fb78d5dee9dd
R3[309] <= 640'h1f0fffff0000000000000023c05fc03eec03f102e007fffffffcffffffffe371ff7cc00800ffb8bf7ef9ffc7ff9692db363fbd5be5a4be3149735d69fd4fbd
R3[310] <= 640'h1800001f7fffff00000000000000410ee19b3ff4038802ff1ffffffffffc0000df20fff8feffffffff7eeff37fff87925f57fca85ef6c9fe595c311ddfc0bfef3eab
R3[311] <= 640'h1800001ffffffc0000000000000083bebe6487fc888c07ffffffe0ff031ffc01807ffffffffebfffff14c657ffffe7e224d8f97d779e8661be1992cc722758b8c3cc
R3[312] <= 640'hf000e31f00001ffcfff8e0000000000007c10797fc83ffaa73efc1021801363fffffffffffff11d97fffff758f70efffbba7e3b21fe6d499c4ac9bca807ca7325ff74fc3
R3[313] <= 640'h400000000000f80f00000000f0e0ffffff00ff0f010000000000213ff3ee031d29cb81768f77ffff8afffffffffffffa7b55fffffd87edfb7fffdaeb946df6bffdd60f1ae156a128dfbc85b96694
R3[314] <= 640'hf0701ff070000ffe7ffffffff00c03f008e47b000007c258e8ffffffffff9ffff75ffffffe5479afffdfd6ae523efffceddd837f595dac62f3fd9d8e3efc7d6673df7d3
R3[315] <= 640'h8000000000400000000000000001ffffffffffffff00fc007fffc007ff09c0a163e31fe848b5fe7f64c7febfffffffffffe0337ffffeff73fbbdbffffee9fd336bb099d3d23f9a49507f62cef3bc2b4e
R3[316] <= 640'h3e7ffffffffffffffef8007eff0c001c00fe00fffff000000038581e1cfcd32c017ffbe3fffe0ffff5fffffff3fffffffffec7bf5d3ffffbb8fb4830cd7f2cec1e1aea488ef78f7fddfe2f
R3[317] <= 640'hfffffff08003ffffffffffffffe0000000007f0001ffffffff000081fcce00ffffeefff9cc2c4ee579feeee7fffbffffffffffcfffffdfd9b6f7ffffb87be369f336a6a3af315ddbab7851f7b2d4dd75
R3[318] <= 640'hff7fff030fc100000ffffffffff0001ffffffffffffeffffe00007071fc4f00730ff188d4c3fb63f8eec947fffffffffff9ff00ffff6da83b35e61ff3e2857ceaacb5546616e69dc025f187935c8f48e
R3[319] <= 640'hc8183ff000073fffffffffffaaabff00e00080f0f0000301f00000001f408000e007e1003cfb71773881e6fffffffffffc9ffc7ffff6ecdcbcd22bffb7353f6f5ba39ce71b17fbdb89e5086fbad05e1d
R3[320] <= 640'hffffc0000000000000000000000000000001603f800000000000003e3cf00001c0003c003c0e800f301fff949ff3fffffffffff70ffe7faaf57ac7d7dc2b3b95ad5dd279a6907a66d15febc57fd81a45
R3[321] <= 640'h700000000000000003fff1f01fc003f1fff808005ffcffff0effe87ffffffffe57ff66a3235e257d79b541ad57411b2e98969b9c66b9a5f95eff9b832
R3[322] <= 640'hfffc7801cc073fe6f800007ff00ff01c05effffffffffe7e7d9393a3df79bcfbe46d6f3cdbed483aa32747b0e7bf754edb570dd
R3[323] <= 640'h107ffc3101ec0433fffdc0000e480008006effffeffffffb3f5fbdd3a5e73a5b6cfb4efb4db30ad80b64baf7a26653dc79795d888
R3[324] <= 640'he000000000000000000000000000000000000000000300000000000001fc80103e000010cffe80fc02000008003dffffffffff97e7e79f2de37fcbaf9835f1bfcd3ddfe1cee30ba50ba28938a6efbfb1
R3[325] <= 640'hf00000000000000000000000000000000000000000030080000000800007000030000003ff3e83f80018070cfeb87fffffffff9aecf399ea36621e7f90b1dbefe6d708c679ff82da5f79efcb3cd615fe
R3[326] <= 640'h80000000000000000000000000000000000000000000ffe8000000c000000000010000071c07fefc039fcff0d37b3f2283ff6ff6d5029bdaed6a1427ffa1e79e2fcde926de7b7fe1a4fdd8e3f50f99bb
R3[327] <= 640'hffffff80000000000000000000000000000000001880fff87c0000047800000001000000002171c1e78078b3f0477f7fffc00615b58e8fffbeff69d79eff6faffd5d6b37d5a7d5ee975a6cf37b7c1714
R3[328] <= 640'h1dffffffffffc0f8023ffeffffffffffffffffffffffffffffffffffffe1000000ffffffefffc00000088400f403183f300007a3f7991d330db27183bf29111fb9d07294967ac05f40bbd0d107fbec4b
R3[329] <= 640'h31fffffffffc0000070f000700000000ffffffffffffff3fff0f00000000061c001ffc0100000007f81fff8021ffffcbfffffeafececfbc9eeaab1dbfd77136f939998cd5abede79cbc7e9a0dddbc583
R3[330] <= 640'h3ffffffffffffffffc00fff8000000ff003c80000000ffffffff00000038000600030007ffffffe7f8fff70100047f833ffffec391cd71b6d7eb79645d7fbdddd6e226ff5a631bea6f1902e96ff9728d
R3[331] <= 640'h4c7c3000008000ffffff0000007fffffffffffffffffffe00000ff7f73fffc07ff3fffff03ff003ffffffffff03ff803c7fffe05065ba9f64d25f9f1d7b97ed65a4005658f06e7a4bbb2c3a90ce19957
R3[332] <= 640'hc51f3fffff00e00000800000001f0000003ecc000000ffc0000fffffe3c001fc000f0ffffffffffffffffffffcffffff0ffffe6ba72b0a57188f9ef1fea9cec1bdd9070d353af4b42bcc176b8aebe7b9
R3[333] <= 640'h590087ffffffffffffffffffc7ffff00fffeffffffffffffffffffffffffffff3fc7f1f8fffffffffffffffffffffffffffe32531f0b730f0755795a377ef9e6f58d18919dbd3e2e5dbff3dafda4db
R3[334] <= 640'hcce1c000000000000000008000830000ffffff000000ff3f1cf0ffcf78fff0fffffffcf8fffff81bc0fffffffffffffffffff5e3edcbcf3d76e675f27ebf51565c24f3d53bed4d7db0d3ef3afea5b7fb
R3[335] <= 640'h30fa0c000000000000000000181c0000000030f81fc02fffff8f0f3ffffeffffffffffffffff7ffdc3fffffffffefffffffff8d7eca245562cf4ded17fe837758f4b729f94dee8e19a909f79ef76c276
R3[336] <= 640'hf83062100000038000000000000000000000000a07000affffeffc3fffffffffffffffffffff7fffff9ff86fffffffffffff99237de5c4bfbf2c505dace8f8ee5bf5fbefdf2cd49dde453cbbfd154e4c
R3[337] <= 640'hef00f09000000000000000000000000000000000070003fffffffeffffffffffffffffffffffffffffffffeffffffffffffff904aa81bd49c957e63e2a28cdaed525f12eba5c449a69854ee3f167fd5f
R3[338] <= 640'h7f1f006f80c10800000000000000000007ffffffffffffffffffffffffffffffffffffffffffffff3ffdfffffffffffffffe6b21e382e1e1976ffc83ba23ece7e497be57b0db91099da123eedbd98dbd
R3[339] <= 640'hcfdc00f38000000000000000000000000fffffffffffffffffffffffffffffffffffffffffffffff9ffffffbfeffffffffff4ec1f61fe7a6d47adcce9539bb5c28adf49d577896768925227fcdd48f6d
R3[340] <= 640'ha27fc20780000000000000000000000007ffffffffffffffffffffffffffffffffffffffffffffffffffff99cfff7ffffff9ee185bbdeb69683bbfedee077a55c2ff5b208072d9affbb7a67de5bdf2bd
R3[341] <= 640'h4cfcc1e00018000000000000000000000000001fffffffffffffffffffffffffffffffffffffdfffffffffff53ff7ffe7ffdbf58c4be5cd188f7ab4b34ec5d5a69d83db0ad14aff28297ad4369ac3d94
R3[342] <= 640'hc9fc02700000000000000000000000000000000fffffffffffffffffffffffffffffffffffff1fffffffffffdbfffffff0fffffe34f439b9ce679dcf5355d40658dd41c37e176ec86838abdfcfe2ad6e
R3[343] <= 640'h2bff4fe80c000018000000000000000000000003ffffffffffffffffffffffffffffffffffffffffffffffe3ffffeefffa4d618d33a7d7d3dde4ec97ddf8857137b083d1ce8bfe39578abf9f9a315ea1
R3[344] <= 640'h23f8e07f0006603000000000000000000000703ffffffffffffffffffffffff6ffffdfffd7fafefdefbf8807fe9e0787f665421f3cb36cd4f0f875d9a9cc7b6789eee8cabafd3c4d84f707524345c84
R3[345] <= 640'h200f870fc701600000000000000000008000070ffffffffffffffffffffffeffff37fbffefd93dfffeff7fc0016cf081b291aeb2f3da73eddc59fbd69a7d7cde77a6eac7aee6b8b637b6f81e308765fc
R3[346] <= 640'h851f8e0ff3f880000000000000000000ff0fffffffffffffffffffffffffffffbf6bffffffbd7ffbdffb7ecffc230800fc3acbb9bc9d478fccff374dea9d22fa476f6ce790ede98f23cc0c65f7885ba3
R3[347] <= 640'h323f0c0007fc99c00000000000000000ff0ffffffffffffffffffffffffffffff343fff5fffdbfb9cc76fcb0000f3e0008076ef7ee64ebd3e7297f75f71933a1bae976db98d3c865eee56fd6f17ce285
R3[348] <= 640'h486707ff3e037fe000000000000000000003ffffffffffffffffffffffa7d1fffdcb99eefffdb581712803ffc007db3e40079b2de73ef25e29f96522b5f947e3275eb6806775c6094009c7b6d2703fc1
R3[349] <= 640'h4efe18007fff0fc00000000000000000000007fffffffffffffffffb01606107fbebe1861778073cc876fc8f0001fe20477c13b1f52edfeecfbb957fe1ef3a5ab65ed04859aa28f61d4fba061d15772f
R3[350] <= 640'h4fffffe3fff0fc07c00000000000000000003ffffffff3ffffffff886f260f247ddadae6800300fc370e43f0200ffffffff73f6d51257b3473fb4efaba132a9ea3f1e43ce024dce9cde387d8e5bde6e
R3[351] <= 640'h1c7fffff00781fe060000000000000000000000b1fffff1ffffffcf9f8e01800bd382d78b85dafe0f73401ce000023ffffbccf8553a8a3aeb9dcfbf1fa27d6025e448b57ef9b15d7fff4bbb29345fa0f
R3[352] <= 640'h53ffffff07c9ec01880000000010002010000201f7ffffffffcfefc01ffffd90bfa6e560c210337f8ffadc00164e3fbfdf6beaae46c8bad42b7b37ffd39eceb7b7d1df2666b6671b506e1d4b3b51f04
R3[353] <= 640'h83ffffffc3ff0708000000000000003190007fff87ffffffd3fe07801ff0e7f06c40eee31f483befa0f9d03ff8e03fffffba4a9d63ecf38d80bd7edfcb962ffcbcb553bd43f8af183424145a7a27edf
R3[354] <= 640'h8e78ffffe03cf813e8f0000040c1fffef1ffcff007ffeffffffc00000ffe0ec40f95acefdea4ffff72fffffffdf83ff7ffbfcb75669d6b38d8ff9d978d9eefe709dc9f2dbdf5b7ab2bd70bd5f80687e
R3[355] <= 640'h88783feffc003fffd9406f90007e7fc3cc7ffff010bf4c1cfffc0000083e275ffbcced57c9c4bdfa579fffffffcffff7fffdcada5f1cd4b9adb6c2b9d59ea4ad7bc873313e5d8b939f62ebb56642d42
R3[356] <= 640'h400007ffffc81fc7e19303800984800a7fffffff801c08377180100700181306387679c799a736bd6e96ffe0f4dfffffef48c7ee3f37cd0c745f8e7d9a75367f75a34b6ab49fea926825acecad8e415
R3[357] <= 640'h1e00000ffff8c40e0039f1c1f0210300447f273bfc07e04c528841e0380000f3c988e3bdfd37c72bc92fddff07c9fffffefce7e7edfbff2bb8b6f88fe42ae1247b5be7f49e446d442100f956e8c36bc3
R3[358] <= 640'h10000003ffffffccf07e0260031d0001f93fbffce60fe07feff041e0008139bba4e8e75eb2dafa4dab95e9dffffdfffffe99de2c450cb165e7dfd55fad397cd8ab2912bd4fcddaa263b2fcbfce1f98d8
R3[359] <= 640'h8a000030fffffffeb19819e5632000061f87f1c7e01ffc06001e01c00186c1ffbfd303cefddeb627cdd8991fffff3ffffd9ff6dfecf4edf6f4dbd6f6f110d97f22bf6995854f364098b55c76e7b2fe3c
R3[360] <= 640'h4400c872ff9cc3ffffc10000c000431ea0001ff87ffff9800008811308007e6fa3550fae8a6afe75fff979ffffe72ffffcdd794aebf860a9f7b7756b97ff8e35706f1a9440657cc1ebe3dddf1eb7b1fd
R3[361] <= 640'h49df1a990ce00000fffff800000f13eff60300fbff3fcafe206701030ff867fbca7c1de8c891fe7a6cf279ffffeffffffefff0eb6cb9ff2f49f037916ae57b1674a750b1a177f0b3bdbddd082e8e3528
R3[362] <= 640'h8a981e10b12000000001fff3ffff07f0aefff0f9c078923b808f30e401fc03e7ddaaab1de4fcfeb75f3bfdfffca6ffffff5ff728fdd9e8f2e99fbe5fec6de3ee905c23e0100584ca89c199cbc8be1d37
R3[363] <= 640'he4aa0c8c8100000000033fffffff1f48a87ff83fdfebf103000f78ed66468feb83a07f58dc3498ff992fcffffc977f7fffd79af38f7275b2f8ff642f84ffda81eb0a6e25210ff74db9cb581abddaef96
R3[364] <= 640'hdf0423dc8080000000030ffcffffff6e717ffc08fe1fddc08101fe6478660fdb2cc5bdb97f01ed3e853f53fffc965e7fff79cb6e351db5df7dca6478f930c48e34c1d271c456fef428d40a64458d0f47
R3[365] <= 640'h2013802d003000000003a0ffffffffd024ffff007e03e1610c0084519cbfa2f9f675f369ecb5bb7ec53e73fffcd6dc6fffedebcef0658fd73bcfb37affdeeea63ea4c269b20621596d9e367ab846865f
R3[366] <= 640'h5012481f05040000000703ff03ffffa05dffff1c03f8961f0f0001a828dc3f739f1f35f67bc2f0a65e30edfffc24f94ffffef3a5c27aff99e0f158fdf9d766cfee57e3a592c85fc96c15239e4bcd13a0
R3[367] <= 640'h8804a1811efe00000707010703fffff0627fffc0107f93807bc38f2a7ef7fff1a6efef8810ddc78cc5256ffffffe3aeefbe4dbaff3e79fb607c7f9e9c8bffe0cc3900751ff2256e2e9220938d8e30550
R3[368] <= 640'h140700bc0024250681000f11603cedffc010bf1ee00edc2e38ebfbfb536de8cfea9454557e750dbfefffda6354bfe5ef45e37cf56fdba7f42def25056be245b64f9d3f962e4e3103997a2e8d93
R3[369] <= 640'hf4004c1c837cc8508fe0307d05afcfff80399fff01fc35fad35c3fffcbecfe017670fa47aaf39cfcffeb64fffff42b57ac24ad907e6af6d9df44f6fa1dff43ac7221fbd50297628394eca3f69
R3[370] <= 640'h1a8004b2ae9b11d00fec63f202e7dfff80c03ffff07ecdde26c8b9dbaa11d8d7d28a3ce1a9f5f7afffcfb3fbf12d7995874714d3b33ee8dea7afee757c1dd86b098373c72857b1f3c36bab382
R3[371] <= 640'h780001c473906667feff08a7931818ff8103ffff01f7fc6b7cc7f9b6daabec42ac3b2d3467bdfffffdb3deffff732713f65feb3ff3efd6fc7bfd06c9e9cd1f6d30bc1860d1d94a762527a087
R3[372] <= 640'hb80001ffcca3dffffff9b722fe1ccdce7070ff00008fc9eaff5fe31525febefdea79c473317d6ffff3fe77df5f9615bb74dbdcd9cf0bd5e1fde3feba2a169d19a8603e98ed9116657c70886
R3[373] <= 640'h7e8028060ea1c1dfffffec00a8e00e30004ffff3f31fa5b23f7d4f786b6d5aacd63a43a3d1da4fffebf7f32ddff7b567b0bf157d62124c37f7d7cce7b527b2974070e555b36a44209de85d5
R3[374] <= 640'h4dd809400e3199fffff000405fff4dc738ff0c4c01a95cbefea338056927e57d13957fb453dfffcffc6dfddff2b7fe16932d52b917765bb5f1d60587320368c4765dd05edca0007eaa0569
R3[375] <= 640'h2c0e800002e6b93effd4120cffff85c06c307c3feefdedee4c53e39cb46e7dd971a1f6d7de740317eef9ffbbf7be5ebffc207ff9feccb1d1f59903b15a30fc900de3376b9058000ad9013a
R3[376] <= 640'h881d800060c766d5b800058fff3c1fe53faef8014bccb61e2be91e122cbdaef1d33cf066e47fffff9bbadf53b0cf153df9efdfebff3f7f87a8173414bb48440be6af17e59d000640023c
R3[377] <= 640'h1fc321880101faae7ec00000f81c007e2077e1190f351dbce0a6dee96709127598358ff767df3d7f77be3f762eb6ae29a3dce44addcd63385e497c39b9a4934054eb71c6a0c00063f0392
R3[378] <= 640'he3c0e0b80003863f74001241001ffe18fcff00966a1cea4a38fbf54fa5f47a0fef3ff8fea7ffb3fbdffbc1544c99e3fbbafd5adfb53e21628ad5825155ef2c0c43b808d60400000c0057
R3[379] <= 640'h510f03cc34001af8e40003b080c3f8ecf423fef904399d03438f09cabe66eebad24f6ae9e7ffcf79ffdde1a843a46aa670ebb72fcee31177fe9392262ff66c0c8070005b980000000023
R3[380] <= 640'h2c803c0620c600962400000c7fff83f83000039241219cec7cfebe4dff29482fe2f1ab3ece9fe7f5b57edeafe965810ac10d018cc9bb730caa0ff750432e041f0028000f800000000022
R3[381] <= 640'h8590c013419ba022ea00434f7780efe1100000f6c64a58bc8e7ac5351a01e0e58fe9b33ddb7ffebeb4f6f79e316081e284065063f67acb1ee2593e5179d5641c00240006000000000022
R3[382] <= 640'he63e80414f30580400411f8080004810fec003309759a6208b67e6abcadedf50ee77adfeffbfcf2e9df679080c31054032eabe2cbdbe798bbdb8ae344c303001260006020000000008
R3[383] <= 640'h1800107ff99238628f0000418989e001118fef10130696605fce6604683cae5b90dfa9dbc413bffbd33f9f76318b052000862621bdd8d80bd4ec201dbc6882016000110003820000000000
R3[384] <= 640'h2000000000002b0fff7fc3f078bc0001dda9f77ff3c3fd08b9a6c8a8eef7b30f14ef2ddbc14438ff3343ffbb7f6edde1e300000001c00ffc9eab697f8062d8d0686000000000000009800000000000
R3[385] <= 640'h15f803fc07ff9b903441dc52a2fffffb7c0183f61ff2462aea80b1fce558f7f998e6d0c6195ffdc9da21a00000000000013e6a71fd51993c9f97600000000000000009800000000000
R3[386] <= 640'h10000000000060ee007f7003f0fffbd002ecbfffff9c4ffc4fade5c77a5ccec4ba125e08775257af733fffbf4d5564c8000000000000039d1086f3cc3f06646c00000000000000009800000000000
R3[387] <= 640'h18000000000003c7ff0007fffffc7e423c6a920ffff017c0d599e12e6f51ade8dff26747faec3857ccfe6b2020b7795e00000000000001813c2c3341d5e72ae7c40000000000000000000000000000
R3[388] <= 640'h10000000000000501effe10000fb47376316088000c00420b5b69c727b20a8b689f63cff69f9408907bcd54f3b4cbec500000000000003c0e8204b3315ec6475000000000000000000000000000000
R3[389] <= 640'h3c000000000002901ffff7ff06760666300f60e0018c610b2d6fa0a212155a29a4c0934ac5ca9d2e92397fff83f9e8000000000000003e0082e69a045dc4f7c030000000000000000000000000000
R3[390] <= 640'h40000000000004e0007ffff8b21de597bff6fffc1f85f85d44b89b3d3c5f4b2c769a626c8f6238c1ee661cdebf54800180000000000110dae477e61fef4800030000000000000000000000000000
R3[391] <= 640'h1200000000000063fe0017066bf4067e6a477c7e00f589569bda13bdb0c98eaecce596d91bfa33f6b77929c6faa3f421b000000000000846124c9afcaebdb88000000000000000000000000000000
R3[392] <= 640'h920000000000000b3ff030180007f180e01f9729a1743a1f1af0067ff1552aa7156f739ebfc1a21a161bc3f018f81001f000000000001f0b39e6ea7817fce00000000000000200000000000000000
R3[393] <= 640'hc20000000000000707ffefffff080ffe161033350e4c069fffc006000468badd09f6dd6ff00060023ba7c07f800000002000000000000f0439266a780fefe00000000000000380000000000000000
R3[394] <= 640'h3c00000000000001407ffffffffe0f1c1d933c4366380e60018004c8007debcddf7d84f04000080cf523a0380f1f0000000800000000000738267884100307c000000000000380000000000000000
R3[395] <= 640'hd70033ff33cff0380ff7f158a46837fffc903b37cf02836dcd149880000000000003e0000f8f80000008000000000006e416f98430000fc000000000000080000000000000000
R3[396] <= 640'h2ffc0000000c0fc7003e0e7b31484300037fff3e3004344283007220000000000503800001f0f0000008000000000000245b8807f0300fc000000000000000000000000000000
R3[397] <= 640'h70000000000000043f800000127f27fc11c90597f87001f02bef3610029d702f6f9e70000000001a10800000e070000000000000000120a65a887fc1f8006000000000000080000000000000000
R3[398] <= 640'h700000000000010111f800003ff01873f87c47cf1877cff7e08704fff22e683308c800c00000f0380000000000000000000000000003fd22744e30c1f8200000000000000080000000000000000
R3[399] <= 640'h8006e31cfff0fff240d9f88b634c8677f797f85fcbfe228081a028000e00001f03a2000003000000000000000000006f9ca56c6684078000000000000000000000000000000000
R3[400] <= 640'h20e70033000078e00099bc0bf857ff89ff85f9bf36fbe2b61c000000000000000000000000000000000000000007e357521e692960000000000000001180000000000000000
R3[401] <= 640'h1cd7e000000001fff907f0012847fff9fe0601e016ec5eb51000000000000000000000000000000000000000000703771bfe69f820000000000000000000000000000000000
R3[402] <= 640'h7e4c13018000007f920f9e98003ffffc02c0c0030376b58000000000000000000000000000000000000000000603ff33fe69fb00100000000000000000000000000000000
R3[403] <= 640'h3679000000ffc03c03ffff7400fe7ffe80122d00bfd47a78000000000000000000000000000000000000000000303ff33fe69fb20000000000000080000000000000000000
R3[404] <= 640'hc00ee1ff1cffffffc0900fc30a07fe3ffe001d3c031bf878700000000000000000000000000000000000000000003f3fb13fc79fc60000000000000080000000000000000000
R3[405] <= 640'h26c000ff8f8ffffff003f844107ff9e00190407f3e259610000000000000000000000000000000000000000001f1e111bc71c260000000000000080000000000000000000
R3[406] <= 640'h30003f00000000103f97801c7607fff8c0018068f611a53010000000000000000000000000000000000000000001b9ec13bc71ce20000000000000080000000000000000000
R3[407] <= 640'h60015c307f0000301f800b44cfd43bfe80000007ffc49d5300000000000000000000000000000000000000000000819f612fc31cdf0000000000000080000000000000000000
R3[408] <= 640'hc3000000000000001660c07f9000002e8e21effb0866c10000c3cff8cf1e210000000000000000000000000000000000000000000c0fe1aac79f2a0000000000000000000000000000000000
R3[409] <= 640'hc4000000000000000c1f00017e3cffc000fc1fef405e0c0000789bf30600010000000000000000000000000000000000000000000c077919c79d58001c000000000000000000000000000000
R3[410] <= 640'h3c000000000000000136877c7e1c00ff8e00071c31c11800009c1394c4000000000000000000000000000000000000000000000000067819c79dd5c01c000000000000000000000000000000
R3[411] <= 640'h3800000000000000005f78000110010106c0ff0f96c184e0000be0881000000000000000000000000000000000000000000000000007f82fc78d1320c3000000000000000000000000000000
R3[412] <= 640'h1fffff783821fffe8e1fe77c008fe00002f210c000000000000000000000000000000000000000000000000007c00607854c4883000000000000000000000000000000
R3[413] <= 640'h2c37fe70100020fde8023fad0fe6000006600810000000000000000000000000000000000000000000000000640004307400d00000000000000000000000000000000
R3[414] <= 640'h200000000000000000028f8007007319f00000001c60d800000103821e0000000000000000000000000000000000000000000000000660004082b27d00000000000000000000000000000000
R3[415] <= 640'h30000000000000000000f08edb3ff0103800c3d17f980000000021180a00000000000000000000000000000000000000000000000007e000008369fd00000000000000000000000000000000
R3[416] <= 640'h1000000000000002bc00000003800108001c7e65450000000230000800200000000000000000000000000000000000000060006e0000003b9fc00000000000000000000000000000100
R3[417] <= 640'he0000000000000dffffee801ff9fffff0006450100000003b820818200000000000000000000000000000000000000002000700000000ff1e00000000000000000000000000000100
R3[418] <= 640'h200000000000001f1ffffe3c0000007f000009c0000008000c806220000000000000000000000000000000000000000000007c0000000200c00000000000000000000000000000000
R3[419] <= 640'h200000000000000fe00001c1fe01800010066f400000000010e01010000000000000000000000000000000000000000000002a0000000000000000000000000000000000000000000
R3[420] <= 640'h10000000000000000537ff8c1000000300100e108200030380c23cc388000000000000000000000000000000000000000010084c0000000000000000000000000000000000000000000
R3[421] <= 640'h100000000000000001a6020000001f8fffbff770f004070e08016b124000000000000000000000000000000000000001801000000000000000000000000000000000000000000000000
R3[422] <= 640'h2009dfdffffc03fffffc7f990941c070c37087c0090000000000000000000000000000000000000018010c021c800000000000000000000000000000000000000000
R3[423] <= 640'h41bf7ffffff000000000600401e20e3f8c1091822000000000000000000000000000000000000000010c830fe00000000000000000000000000000000000000000
R3[424] <= 640'hac9dc00f818018e73c000058013f3c60010020080000060000000000000000000000000000010044188707d24000000000000000000000000000000000000000
R3[425] <= 640'h64f4003800013f0ffffffff90000e3f0008a821900000600000000000000000000000000000007e13986848f6000000000000000000000000000000000000000
R3[426] <= 640'h4000000000000ab8000fc103ffffe7ffff8f20000077f02122000000000000000000000000000000000000000761390605380000000000006000000000000000000000000000
R3[427] <= 640'hc000000000000460ffeffff9ffe00000e0e370c68b0000205400000000000000000000000000000000000000001939871c90000c00000000a000000000000000000000000000
R3[428] <= 640'h40000000f1000000000000ddfff83fff00007efeffdff81f60b59102820000000000000000000000000000000000000000f811c79f65600c00000000a000000000000000000000000000
R3[429] <= 640'h40000000ff000000000000219e396000001fffffffff0480c01fe30360000000000000000000000000000000000000000ec819c784e1e0c30000c0186000000000000000000000000000
R3[430] <= 640'h70000000ff0000000000000c00c0188007fffffffc00033303f3b0638e000000000000000000000000000000000000000f40080388f649830001f8380000000000000000000000000000
R3[431] <= 640'h7f00000000000003dfe03120fffff8000000000138e8c25c00000000000000000000000000000000000000000060000317b07808000700208000000000000000000000000000
R3[432] <= 640'h300ffc00000000000007819fffffffc0100071fff4a72a440000c000001000000000000200800000000000000000270000380383800000000000000000000000000000000000000
R3[433] <= 640'hffc000000000000057ffffe77e00000037ff00003eff80000c0900031000000000000700000000000000000006e0000183e6f800000000000000000000000000000000000000
R3[434] <= 640'h7fe000000000000014fff000003c010300610104fe0e27014c00001c180000000000070000000000000000000ee0000003395e00000080000000000000000000000000000000
R3[435] <= 640'hf0000000000000030300ff7cc038f00000f180000676c37c000036000000000000000018000000000000000500000000fc1e00000000000000000000000000000100000000
R3[436] <= 640'hf000000000000000bd1fe000000c0100e3e000000676fffc0200030000000000800000180000000000000007c4000030000c00000000000000000000000000000100000000
R3[437] <= 640'h30000f8f0000000000000297e000c800003f9800000000477fffc0000000000000007400000000000000000000000a0000000000000000000000000000000000000000000000000
R3[438] <= 640'hfcf00000000000001a000000001ee0fc00000000003fffec720000000000000fc0000000000000000000000760000000000000000000000000000000000000000000000000
R3[439] <= 640'h7cf000000000008003e00000e7f0380000000000023fffccb4219f000000000400000000000000000000000000000000000000000c00000000000000000000000000000000
R3[440] <= 640'h8000018400000000002000f903ff7d1e000000000000037fe7ec037fc300000000000000000000000000000000000c000000000000000600000000000000000000000400000000
R3[441] <= 640'hc000000000000000163cfcde000000000000000033fffcc7804000000000000000000000000000000000000e0000000000008c110000000000000000000000000000e000
R3[442] <= 640'h7000000000000000007e7e00000000000000000013fffcf540e0000000000000000000000000000000000000000000000000000180000000000000000000000000000000
R3[443] <= 640'h71000000000001000402800000000000000000007ffffcfb8040000000000000000000000000000000000000000000000000000000000000000000000000000000000000
R3[444] <= 640'h71000000000003100000000000000000000000017ffffcffbc8000000000000000000000000000000000000f000000000080c06000000000000000000000000000000000
R3[445] <= 640'hf10000000000003000000000ff000000000000203fff7cac000000000000000000000000000000000000000e000000000000002000000000000000000000000000000000
R3[446] <= 640'hfc0000000000000080800000c08c00000000006001c36e80000000000000000000000000000000000000000000000000000001b0f0000000000000000000000000000000
R3[447] <= 640'h800000ce00000000000080300000100fcc00000000006001c34e0000000000000000000000000000000000000060000000000002dcc4daf0000000000000000000000000000000
R3[448] <= 640'h18000000031fe00fe7900000610687e600000000001800000010000000000000040000201c0000008001f8d40f80000000000000000000000000000000
R3[449] <= 640'h100000000000000000000000c0000001ffe040de5e0000060060776000000000000000000a40000010080000000009201000000002d78600c00000000000000000000000000000000
R3[450] <= 640'h3000000000000000000000000000000fffc800fe110000060001726000000000000000000860000389100000000000c83000c0052870060000000e000000000000000000000000000
R3[451] <= 640'h3fb00800fe91000003000333e0000000000000000004ec000004000000000000260000e000603c3f1400000f800008000000000000000000000
R3[452] <= 640'hf0008076fe9000000200803fec00000000000800000207dea0019800000000000000000006080808c4000000000000000000000000000000000
R3[453] <= 640'hc00fe302fe6000000201903b6800000000000000000005dd20041e0000000000000000000044008018000000000008000010000000000000000
R3[454] <= 640'h20fc00fc016fe000000020000000000000000000000000071c4a6180e80000001860d600020031005c86000000800000c000000080800018000400
R3[455] <= 640'h20020f807f01f3ff80000000000000000000000000078000002bcf292300c1fb8511dfe1d00000000020c0000003000002187fffc00fccce3f8000e00
R3[456] <= 640'h441fc18f091e7f0000000608000000200000000012bc8d400fc600a0080470c566538450002000000180137cfb0ffff82691ff2807efe67b2810000
R3[457] <= 640'h1c79dfe1c1ff0000060600f0201154000110ab01040eec00002590638b2daac0d06ec000300c9040dff9fbfbfe0001feffcf1f07ef767be200000
R3[458] <= 640'h18000000000040019bff703ff000004060716532ea37468f0040000005c0000f8806ffe09d3b7680c080f13fddcf0dff3a579e00001fe7fffff00e3723be701300
R3[459] <= 640'h2800000000ee480081fe003fe000000f780a277e00588708800000000000001c000007e00259fc3da75b09ffd9ca09fffe779ff0c383e30ffff80e370e9e303300
R3[460] <= 640'h7000000000ffccff81f80007c000001538000000000000000000040000100018017ebb611f9efb1393100069fdcac99fd21e7f000083f1e3ffcc0f070f9f801000
R3[461] <= 640'h4000000003ffcfb7fffc801f800000080800000000000041000000000000003fefdefe66026ec0bf96f84128ffaac993825bff800019f9f7ffec03838487880700
R3[462] <= 640'h14000000007ffceb7ffff407fe00000000000000002f0180000000000000000260cdfc3f3615c47c3d94cd0b87fab7a899a7bb7ffff19f93ffffe00838687880460
R3[463] <= 640'h180021000000010000000003ffcedfffff403ef80000a400000000020c340c00000000000000228033a361904e2fff521364497aaf79819212f700101ff8fffffe00003b879803e0
R3[464] <= 640'h2000000000300018049000300e1c0000000001ffc8de7fffc8fff800001211528e5f400100000000000000000030000dd5200045a77fc063ae23fab7cc9dfa52ff03ffff713ff1fff0208ff38c3160
R3[465] <= 640'h30300000000020000001803531e300000000023ffcff0ffffc8fff800000008104809080000000000000000000034f082e76040c889f0e39b9c38f0b5c261c298fc07f8fffce1f1e6e80613fa383100
R3[466] <= 640'h6c0c001008000000fdc063003200000000033ffec00ffffe8fffd000006480449800100000000000000000000000000c0000001e5ff29cac34072b5c2c046f8fe00f833fc83f1fee4000e99c01000
R3[467] <= 640'h79fc0000000001f8014bb000e000000000003ffec01ffffe8fffd80008011004fb000000000000000000000000f30000000000000000b4a1c0a011300007ccf39f803000020004000000000000000
R3[468] <= 640'h3c0000001fff60006252c44a000000000003ffe000ffffe8fffd800000114ecf44040000000000000000000010000060e800000013e1e8d218301300000000000000000001000c07a0039cc40200
R3[469] <= 640'h21f80000002fffe000f42d0aec000000000003ffe000ffffe8fffd80000011c2cd15800000000000000000000010fffca01801c10003e1222201105b2663fcef3f1ff3e0fb7fc7fa0700019c000000
R3[470] <= 640'hffc0000001f0ffc00034240300000000000003ffe800ffffe87ff880000010420d199000cc00000000000000000bffff0000095c0000042c398f261a6736c6287f1fff87ff3feff860000000200400
R3[471] <= 640'hfff8000001af4000000366f4180000000000003fff800ffffe87ff8800000106209c14200000000000000000000087cff000109eb6200001dffe74e9ae71ecca77fff7fff9c19de8938180008481700
R3[472] <= 640'h40dc8000071f3e000000a261000000000000003ffffc00ffffe0fffc8000003022030d8e80008000000000000000084686c189f8b83c00000009e1f808e71b359565f3a87c349660408b48043d541700
R3[473] <= 640'h624b80010ffc0000c0006406400000000000003ffffc00fffff0fffc8000002040004dd0800d80000000000000000e00629f467a1ec0000000003b1e86071c35d6053c02107c9506798808042a690000
R3[474] <= 640'h5081073147f0000100006f1ee0000000000003fffff800fffff07ffc8000002040006d70000e20000000000000000d703f11d6fe18000000000001eea7a7000000001048713903e630003e0309000080
R3[475] <= 640'h400107fdc600000000016d2b00000000000003e7fff800ffffe07ffc0000001060006894000000000000000000004abcf905de9ff000000000000001828380000000c2dff397083f9828ab0000000000
R3[476] <= 640'h407fc0b0020300000380c39a00000000000003f7fffc00ffffe07ffc800000004000280e2e000288000000000000097c6604a81e000000000000000020f600021961c17a2ee900330629506000000800
R3[477] <= 640'h1eff38f8260000000fdfa48300000000000000ffffff00ffffe07ffc80000800500020000c004c800000000000000000000366e00000000000000000000200138048f135bd03a00d4e0c6860c6200002
R3[478] <= 640'h7c33c04e200000000144801000000000000037fffff00ffffe07ffc80001c00900013c606004078000000000000000000009800000000000000000000c20001721a840f1fc408eeb001c1100518061b
R3[479] <= 640'h6fff1e8c408000000028034a000000000000037ff7fc00fffff07ffc80000c0001000000000241d10000000000000000000060000000000000000000000e83800c52df176e064930016c0008418d020c
end
//**************************Main Code************************
always @(posedge vga_clk or posedge sys_rst_n) begin
    if(sys_rst_n)   pixel_data <= 12'd0;
    else begin
        pixel_data <= {R0[pixel_y][pixel_x], R1[pixel_y][pixel_x], R2[pixel_y][pixel_x], R3[pixel_y][pixel_x],
                       G0[pixel_y][pixel_x], G1[pixel_y][pixel_x], G2[pixel_y][pixel_x], G3[pixel_y][pixel_x],
                       B0[pixel_y][pixel_x], B1[pixel_y][pixel_x], B2[pixel_y][pixel_x], B3[pixel_y][pixel_x]};
    end
    
end  
endmodule


// The whole VGA 
module VGA_out(
    input sys_clk,
    input sys_rst_n,
    input [1:0] choise,
    //VGA
    output vga_hs,
    output vga_vs,
    output [11:0] vga_rgb);

//Wire define
wire vga_clk_w;
wire [11:0] pixel_data;
wire [9:0] pixel_x;
wire [9:0] pixel_y;

//****************************Main Code**************************
// 这样的话每个VGA输出都有个时钟分频
//优化的时候可以将时钟分频拿出来
clockDiv clkdiv1(
     .sys_clk(sys_clk),         
     .sys_rst_n(sys_rst_n),
     .clk_25M(vga_clk_w));

vga_driver VGAdriver1(
    .vga_clk(vga_clk_w),   
    .sys_rst_n(sys_rst_n),
  
    .vga_hs(vga_hs),      // 行同步
    .vga_vs(vga_vs),      // 场同步
    .vga_rgb(vga_rgb),      //4+4+4
    
    .pixel_data(pixel_data),    //像素点RGB data
    .pixel_x(pixel_x),       //像素点横坐标
    .pixel_y(pixel_y)        //像素点纵坐标
);
 
vga_display vgadisplay1(
    .vga_clk(vga_clk_w),
    .sys_rst_n(sys_rst_n),
    .pixel_x(pixel_x),
    .pixel_y(pixel_y),
    .choise(choise),
    .pixel_data(pixel_data));

endmodule